magic
tech sky130A
magscale 1 2
timestamp 1713426604
<< metal1 >>
rect 19004 11954 21138 12054
rect 10962 11860 15460 11942
rect 10962 11004 11068 11860
rect 15322 11250 15460 11860
rect 15322 11004 15470 11250
rect 10962 10078 15470 11004
rect 19004 11018 19080 11954
rect 21044 11018 21138 11954
rect 19004 10132 21138 11018
rect 23416 11674 26996 11726
rect 23416 10966 23462 11674
rect 26906 10966 26996 11674
rect 23416 10178 26996 10966
rect 21397 8694 21743 8700
rect 20817 8348 21397 8694
rect 21397 8342 21743 8348
rect 10968 3648 16968 4786
rect 10968 2280 11078 3648
rect 12838 3624 16968 3648
rect 12838 2280 14866 3624
rect 10968 2256 14866 2280
rect 16736 2256 16968 3624
rect 10968 2134 16968 2256
rect 18860 3640 21256 7088
rect 25532 4618 29374 4622
rect 18860 2334 18928 3640
rect 21146 2334 21256 3640
rect 23420 3722 29374 4618
rect 23420 2624 23464 3722
rect 25520 3680 29374 3722
rect 25520 2704 27196 3680
rect 29232 2704 29374 3680
rect 25520 2624 29374 2704
rect 23420 2590 29374 2624
rect 23420 2588 25584 2590
rect 18860 2198 21256 2334
<< via1 >>
rect 11068 11004 15322 11860
rect 19080 11018 21044 11954
rect 23462 10966 26906 11674
rect 21397 8348 21743 8694
rect 11078 2280 12838 3648
rect 14866 2256 16736 3624
rect 18928 2334 21146 3640
rect 23464 2624 25520 3722
rect 27196 2704 29232 3680
<< metal2 >>
rect 19004 11954 21138 12054
rect 10986 11860 15414 11924
rect 10986 11004 11068 11860
rect 15322 11004 15414 11860
rect 10986 10940 15414 11004
rect 19004 11018 19080 11954
rect 21044 11018 21138 11954
rect 19004 10132 21138 11018
rect 23432 11674 26964 11700
rect 23432 10966 23462 11674
rect 26906 10966 26964 11674
rect 23432 10934 26964 10966
rect 21391 8348 21397 8694
rect 21743 8348 21749 8694
rect 16782 6190 18184 6310
rect 10398 5888 11182 6062
rect 10398 4363 10572 5888
rect 18064 4741 18184 6190
rect 21397 5968 21743 8348
rect 29228 6110 30226 6230
rect 21397 5966 22782 5968
rect 21397 5814 23612 5966
rect 21397 5810 22350 5814
rect 21445 5282 21619 5810
rect 21441 5118 21450 5282
rect 21614 5118 21623 5282
rect 21445 5113 21619 5118
rect 10398 4189 12003 4363
rect 12177 4189 12186 4363
rect 11030 3648 12972 3784
rect 11030 2280 11078 3648
rect 12838 2280 12972 3648
rect 11030 2170 12972 2280
rect 13346 1868 13466 4676
rect 13806 4544 14010 4664
rect 18060 4631 18069 4741
rect 18179 4631 18188 4741
rect 18064 4626 18184 4631
rect 12260 1748 13466 1868
rect 11287 1076 11397 1080
rect 12260 1076 12380 1748
rect 13890 1595 14010 4544
rect 14732 3624 16882 3770
rect 14732 2256 14866 3624
rect 16736 2256 16882 3624
rect 18870 3640 21196 3732
rect 18870 2334 18928 3640
rect 21146 2334 21196 3640
rect 23438 3722 25564 3772
rect 23438 2624 23464 3722
rect 25520 2624 25564 3722
rect 23438 2606 25564 2624
rect 18870 2290 21196 2334
rect 14732 2158 16882 2256
rect 13886 1485 13895 1595
rect 14005 1485 14014 1595
rect 13890 1480 14010 1485
rect 25794 1433 25914 4582
rect 26314 4122 26434 4572
rect 30106 4147 30226 6110
rect 26901 4122 27011 4126
rect 26314 4117 27016 4122
rect 26314 4007 26901 4117
rect 27011 4007 27016 4117
rect 30102 4037 30111 4147
rect 30221 4037 30230 4147
rect 30106 4032 30226 4037
rect 26314 4002 27016 4007
rect 26901 3998 27011 4002
rect 27168 3680 29272 3734
rect 27168 2704 27196 3680
rect 29232 2704 29272 3680
rect 27168 2678 29272 2704
rect 25790 1323 25799 1433
rect 25909 1323 25918 1433
rect 25794 1318 25914 1323
rect 11282 1071 12380 1076
rect 11282 961 11287 1071
rect 11397 961 12380 1071
rect 11282 956 12380 961
rect 11287 952 11397 956
<< via2 >>
rect 11068 11004 15322 11860
rect 19080 11018 21044 11954
rect 23462 10966 26906 11674
rect 21450 5118 21614 5282
rect 12003 4189 12177 4363
rect 11078 2280 12838 3648
rect 18069 4631 18179 4741
rect 14866 2256 16736 3624
rect 18928 2334 21146 3640
rect 23464 2624 25520 3722
rect 13895 1485 14005 1595
rect 26901 4007 27011 4117
rect 30111 4037 30221 4147
rect 27196 2704 29232 3680
rect 25799 1323 25909 1433
rect 11287 961 11397 1071
<< metal3 >>
rect 19004 11954 21138 12054
rect 10986 11860 15414 11924
rect 10986 11004 11068 11860
rect 15322 11004 15414 11860
rect 10986 10940 15414 11004
rect 19004 11018 19080 11954
rect 21044 11018 21138 11954
rect 19004 10132 21138 11018
rect 23432 11674 26964 11700
rect 23432 10966 23462 11674
rect 26906 10966 26964 11674
rect 23432 10934 26964 10966
rect 17449 5282 21619 5287
rect 17449 5118 21450 5282
rect 21614 5118 21619 5282
rect 17449 5113 21619 5118
rect 11998 4363 12182 4368
rect 17449 4363 17623 5113
rect 11998 4189 12003 4363
rect 12177 4189 17623 4363
rect 18064 4741 18184 4746
rect 18064 4631 18069 4741
rect 18179 4631 18184 4741
rect 11998 4184 12182 4189
rect 11030 3648 12972 3784
rect 11030 2280 11078 3648
rect 12838 2280 12972 3648
rect 11030 2170 12972 2280
rect 14732 3624 16882 3770
rect 14732 2256 14866 3624
rect 16736 2256 16882 3624
rect 14732 2158 16882 2256
rect 13648 1595 14010 1600
rect 13648 1485 13895 1595
rect 14005 1485 14010 1595
rect 13648 1480 14010 1485
rect 9233 1076 9351 1081
rect 9232 1075 11402 1076
rect 9232 957 9233 1075
rect 9351 1071 11402 1075
rect 9351 961 11287 1071
rect 11397 961 11402 1071
rect 9351 957 11402 961
rect 9232 956 11402 957
rect 9233 951 9351 956
rect 13648 567 13768 1480
rect 18064 585 18184 4631
rect 30106 4147 30226 4152
rect 26896 4117 27016 4122
rect 26896 4007 26901 4117
rect 27011 4007 27016 4117
rect 18870 3640 21196 3732
rect 18870 2334 18928 3640
rect 21146 2334 21196 3640
rect 23438 3722 25564 3772
rect 23438 2624 23464 3722
rect 25520 2624 25564 3722
rect 23438 2606 25564 2624
rect 18870 2290 21196 2334
rect 22480 1433 25914 1438
rect 22480 1323 25799 1433
rect 25909 1323 25914 1433
rect 22480 1318 25914 1323
rect 22480 627 22600 1318
rect 26896 673 27016 4007
rect 30106 4037 30111 4147
rect 30221 4037 30226 4147
rect 27168 3680 29272 3734
rect 27168 2704 27196 3680
rect 29232 2704 29272 3680
rect 27168 2678 29272 2704
rect 30106 941 30226 4037
rect 30101 823 30107 941
rect 30225 823 30231 941
rect 30106 822 30226 823
rect 13643 449 13649 567
rect 13767 449 13773 567
rect 18059 467 18065 585
rect 18183 467 18189 585
rect 22475 509 22481 627
rect 22599 509 22605 627
rect 26891 555 26897 673
rect 27015 555 27021 673
rect 30106 614 30226 620
rect 26896 554 27016 555
rect 22480 508 22600 509
rect 30101 495 30106 613
rect 30226 495 30231 613
rect 30106 488 30226 494
rect 18064 466 18184 467
rect 13648 448 13768 449
<< via3 >>
rect 11068 11004 15322 11860
rect 19080 11018 21044 11954
rect 23462 10966 26906 11674
rect 11078 2280 12838 3648
rect 14866 2256 16736 3624
rect 9233 957 9351 1075
rect 18928 2334 21146 3640
rect 23464 2624 25520 3722
rect 27196 2704 29232 3680
rect 30107 823 30225 941
rect 13649 449 13767 567
rect 18065 467 18183 585
rect 22481 509 22599 627
rect 26897 555 27015 673
rect 30106 494 30226 614
<< metal4 >>
rect 798 44634 858 45152
rect 1534 44634 1594 45152
rect 2270 44634 2330 45152
rect 3006 44634 3066 45152
rect 3742 44634 3802 45152
rect 4478 44634 4538 45152
rect 5214 44634 5274 45152
rect 5950 44634 6010 45152
rect 6686 44634 6746 45152
rect 7422 44634 7482 45152
rect 8158 44634 8218 45152
rect 8894 44634 8954 45152
rect 9630 44634 9690 45152
rect 10366 44634 10426 45152
rect 11102 44634 11162 45152
rect 11838 44634 11898 45152
rect 12574 44634 12634 45152
rect 13310 44634 13370 45152
rect 14046 44634 14106 45152
rect 14782 44634 14842 45152
rect 15518 44634 15578 45152
rect 16254 44634 16314 45152
rect 16990 44634 17050 45152
rect 17726 44634 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 798 44574 31358 44634
rect 3742 44572 3802 44574
rect 200 12624 500 44152
rect 31298 44136 31358 44574
rect 200 11954 30536 12624
rect 200 11860 19080 11954
rect 200 11004 11068 11860
rect 15322 11018 19080 11860
rect 21044 11674 30536 11954
rect 21044 11018 23462 11674
rect 15322 11004 23462 11018
rect 200 10966 23462 11004
rect 26906 10966 30536 11674
rect 200 10942 30536 10966
rect 200 10918 18764 10942
rect 21574 10918 30536 10942
rect 200 1000 500 10918
rect 19922 3800 20160 3808
rect 31172 3800 31472 44136
rect 10264 3722 31472 3800
rect 10264 3648 23464 3722
rect 10264 2280 11078 3648
rect 12838 3640 23464 3648
rect 12838 3624 18928 3640
rect 12838 2280 14866 3624
rect 10264 2256 14866 2280
rect 16736 2334 18928 3624
rect 21146 2624 23464 3640
rect 25520 3680 31472 3722
rect 25520 2704 27196 3680
rect 29232 2704 31472 3680
rect 25520 2624 31472 2704
rect 21146 2334 31472 2624
rect 16736 2256 31472 2334
rect 10264 2094 31472 2256
rect 9232 1075 9352 1076
rect 9232 957 9233 1075
rect 9351 957 9352 1075
rect 31172 984 31472 2094
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 957
rect 30106 941 30226 942
rect 30106 823 30107 941
rect 30225 823 30226 941
rect 26896 673 27016 674
rect 22480 627 22600 628
rect 18064 585 18184 586
rect 13648 567 13768 568
rect 13648 449 13649 567
rect 13767 449 13768 567
rect 13648 0 13768 449
rect 18064 467 18065 585
rect 18183 467 18184 585
rect 18064 0 18184 467
rect 22480 509 22481 627
rect 22599 509 22600 627
rect 22480 0 22600 509
rect 26896 555 26897 673
rect 27015 555 27016 673
rect 30106 615 30226 823
rect 26896 0 27016 555
rect 30105 614 30227 615
rect 30105 494 30106 614
rect 30226 494 31432 614
rect 30105 493 30227 494
rect 31312 0 31432 494
use opamp  opamp_0
timestamp 1713422843
transform 1 0 21426 0 1 7506
box 1988 -3100 7988 2900
use opamp  opamp_1
timestamp 1713422843
transform 1 0 8980 0 1 7586
box 1988 -3100 7988 2900
use vbias_resistor  vbias_resistor_0
timestamp 1713420874
transform 1 0 17820 0 1 7778
box 1048 -958 3482 2578
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 31172 984 31472 44136 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>

* NGSPICE file created from p3_opamp_parax.ext - technology: sky130A

.subckt p3_opamp_parax VDD MINUS PLUS VOUT VSS
X0 VDD.t63 a_6022_n861.t13 a_9426_n851.t2 VDD.t62 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X1 VOUT.t19 a_9426_n851.t7 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 VOUT.t18 a_9426_n851.t8 VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 VOUT.t17 a_9426_n851.t9 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 VOUT.t16 a_9426_n851.t10 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X5 VDD.t61 a_6022_n861.t14 a_9426_n851.t5 VDD.t60 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X6 a_6022_n861.t3 a_6022_n861.t2 VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X7 a_9426_n851.t1 a_6022_n861.t15 VDD.t57 VDD.t56 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X8 VOUT.t15 a_9426_n851.t11 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X9 VDD.t35 a_9426_n851.t12 VOUT.t14 VDD.t34 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X10 VDD.t55 a_6022_n861.t4 a_6022_n861.t5 VDD.t54 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X11 VDD.t33 a_9426_n851.t13 VOUT.t13 VDD.t32 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X12 VSS.t32 VBIAS VX.t5 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X13 a_6022_n861.t1 a_6022_n861.t0 VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X14 VDD VBIAS VSS.t2 sky130_fd_pr__res_xhigh_po_0p35 l=2.8
X15 VDD.t31 a_9426_n851.t14 VOUT.t12 VDD.t30 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X16 VBIAS VBIAS VSS.t30 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X17 VOUT.t11 a_9426_n851.t15 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X18 VX.t3 VBIAS VSS.t28 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X19 VDD.t51 a_6022_n861.t16 a_9426_n851.t0 VDD.t50 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X20 a_9426_n851.t3 a_6022_n861.t17 VDD.t49 VDD.t48 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X21 VOUT.t10 a_9426_n851.t16 VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X22 VSS.t26 VBIAS VX.t2 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X23 VOUT.t9 a_9426_n851.t17 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X24 VBIAS VBIAS VSS.t24 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X25 a_9426_n851.t4 a_6022_n861.t18 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X26 VX.t4 VBIAS VSS.t22 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X27 a_6022_n861.t12 MINUS.t0 VX.t0 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.5
X28 a_9426_n851.t6 PLUS.t0 VX.t1 VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.5
X29 VSS.t20 VBIAS VOUT.t26 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X30 VDD.t17 a_9426_n851.t18 VOUT.t8 VDD.t16 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X31 VSS.t18 VBIAS VBIAS VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X32 VDD.t15 a_9426_n851.t19 VOUT.t7 VDD.t14 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X33 VSS.t16 VBIAS VBIAS VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X34 VDD.t13 a_9426_n851.t20 VOUT.t6 VDD.t12 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X35 VOUT.t24 VBIAS VSS.t14 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=2
X36 a_6022_n861.t7 a_6022_n861.t6 VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X37 VDD.t11 a_9426_n851.t21 VOUT.t5 VDD.t10 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X38 VOUT.t21 VBIAS VSS.t12 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X39 VDD.t9 a_9426_n851.t22 VOUT.t4 VDD.t8 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X40 VSS.t10 VBIAS VOUT.t20 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X41 VOUT.t22 VBIAS VSS.t8 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X42 VDD.t7 a_9426_n851.t23 VOUT.t3 VDD.t6 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X43 VSS.t6 VBIAS VOUT.t25 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X44 VDD.t5 a_9426_n851.t24 VOUT.t2 VDD.t4 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X45 VOUT.t1 a_9426_n851.t25 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X46 VDD.t43 a_6022_n861.t8 a_6022_n861.t9 VDD.t42 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
X47 VDD.t41 a_6022_n861.t10 a_6022_n861.t11 VDD.t40 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=2
X48 VOUT.t0 a_9426_n851.t26 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X49 VOUT.t23 VBIAS VSS.t4 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=2
R0 a_6022_n861.n11 a_6022_n861.t1 228.615
R1 a_6022_n861.n7 a_6022_n861.t11 228.284
R2 a_6022_n861.n6 a_6022_n861.n14 200.05
R3 a_6022_n861.n6 a_6022_n861.n12 200.05
R4 a_6022_n861.n4 a_6022_n861.t15 53.2404
R5 a_6022_n861.n8 a_6022_n861.t15 53.0562
R6 a_6022_n861.t16 a_6022_n861.n4 52.0225
R7 a_6022_n861.n8 a_6022_n861.t16 52.0225
R8 a_6022_n861.t18 a_6022_n861.n4 52.0225
R9 a_6022_n861.n8 a_6022_n861.t18 52.0225
R10 a_6022_n861.n5 a_6022_n861.t14 52.0225
R11 a_6022_n861.t14 a_6022_n861.n9 52.0225
R12 a_6022_n861.n5 a_6022_n861.t17 52.0225
R13 a_6022_n861.t17 a_6022_n861.n9 52.0225
R14 a_6022_n861.t13 a_6022_n861.n13 52.0225
R15 a_6022_n861.n10 a_6022_n861.t13 52.0225
R16 a_6022_n861.n2 a_6022_n861.n11 0.72045
R17 a_6022_n861.n2 a_6022_n861.t0 25.6523
R18 a_6022_n861.t4 a_6022_n861.n6 52.0225
R19 a_6022_n861.n3 a_6022_n861.t4 52.0225
R20 a_6022_n861.t10 a_6022_n861.n0 25.5988
R21 a_6022_n861.n7 a_6022_n861.n0 0.827361
R22 a_6022_n861.n1 a_6022_n861.t2 52.0225
R23 a_6022_n861.t2 a_6022_n861.n6 52.0225
R24 a_6022_n861.n1 a_6022_n861.t8 52.0225
R25 a_6022_n861.t8 a_6022_n861.n6 52.0225
R26 a_6022_n861.t6 a_6022_n861.n3 52.0225
R27 a_6022_n861.n6 a_6022_n861.t6 52.0225
R28 a_6022_n861.t12 a_6022_n861.n6 38.0282
R29 a_6022_n861.n14 a_6022_n861.t9 28.5655
R30 a_6022_n861.n14 a_6022_n861.t3 28.5655
R31 a_6022_n861.n12 a_6022_n861.t5 28.5655
R32 a_6022_n861.n12 a_6022_n861.t7 28.5655
R33 a_6022_n861.n1 a_6022_n861.n0 3.41613
R34 a_6022_n861.n3 a_6022_n861.n1 2.58927
R35 a_6022_n861.n5 a_6022_n861.n4 2.43874
R36 a_6022_n861.n13 a_6022_n861.n5 2.36344
R37 a_6022_n861.n11 a_6022_n861.n6 2.22134
R38 a_6022_n861.n6 a_6022_n861.n7 2.20242
R39 a_6022_n861.n11 a_6022_n861.n10 1.70389
R40 a_6022_n861.n3 a_6022_n861.n2 2.01483
R41 a_6022_n861.n13 a_6022_n861.n11 1.34609
R42 a_6022_n861.n9 a_6022_n861.n8 2.06781
R43 a_6022_n861.n10 a_6022_n861.n9 2.06781
R44 a_9426_n851.n4 a_9426_n851.t10 240.778
R45 a_9426_n851.t10 a_9426_n851.n3 240.778
R46 a_9426_n851.n1 a_9426_n851.t9 119.816
R47 a_9426_n851.t18 a_9426_n851.n0 119.504
R48 a_9426_n851.n1 a_9426_n851.t25 119.677
R49 a_9426_n851.t14 a_9426_n851.n1 119.501
R50 a_9426_n851.n0 a_9426_n851.t17 240.349
R51 a_9426_n851.t17 a_9426_n851.n2 240.349
R52 a_9426_n851.t21 a_9426_n851.n0 240.349
R53 a_9426_n851.n2 a_9426_n851.t21 240.349
R54 a_9426_n851.t7 a_9426_n851.n0 240.349
R55 a_9426_n851.n2 a_9426_n851.t7 240.349
R56 a_9426_n851.n0 a_9426_n851.t22 240.349
R57 a_9426_n851.t22 a_9426_n851.n2 240.349
R58 a_9426_n851.n0 a_9426_n851.t8 240.349
R59 a_9426_n851.t8 a_9426_n851.n2 240.349
R60 a_9426_n851.t13 a_9426_n851.n0 240.349
R61 a_9426_n851.n2 a_9426_n851.t13 240.349
R62 a_9426_n851.t16 a_9426_n851.n0 240.349
R63 a_9426_n851.n2 a_9426_n851.t16 240.349
R64 a_9426_n851.n3 a_9426_n851.t19 240.349
R65 a_9426_n851.t19 a_9426_n851.n2 240.349
R66 a_9426_n851.n3 a_9426_n851.t11 240.349
R67 a_9426_n851.t11 a_9426_n851.n4 240.349
R68 a_9426_n851.t20 a_9426_n851.n3 240.349
R69 a_9426_n851.n4 a_9426_n851.t20 240.349
R70 a_9426_n851.t26 a_9426_n851.n3 240.349
R71 a_9426_n851.n4 a_9426_n851.t26 240.349
R72 a_9426_n851.n3 a_9426_n851.t12 240.349
R73 a_9426_n851.t12 a_9426_n851.n4 240.349
R74 a_9426_n851.n3 a_9426_n851.t15 240.349
R75 a_9426_n851.t15 a_9426_n851.n4 240.349
R76 a_9426_n851.t23 a_9426_n851.n3 240.349
R77 a_9426_n851.n4 a_9426_n851.t23 240.349
R78 a_9426_n851.n1 a_9426_n851.t24 119.882
R79 a_9426_n851.n5 a_9426_n851.t2 229.762
R80 a_9426_n851.n1 a_9426_n851.t1 228.216
R81 a_9426_n851.n5 a_9426_n851.n7 200.619
R82 a_9426_n851.n5 a_9426_n851.n6 200.614
R83 a_9426_n851.t6 a_9426_n851.n5 36.3657
R84 a_9426_n851.n6 a_9426_n851.t0 28.5655
R85 a_9426_n851.n6 a_9426_n851.t4 28.5655
R86 a_9426_n851.n7 a_9426_n851.t5 28.5655
R87 a_9426_n851.n7 a_9426_n851.t3 28.5655
R88 a_9426_n851.n0 a_9426_n851.n3 5.15267
R89 a_9426_n851.n4 a_9426_n851.n2 4.72333
R90 a_9426_n851.n5 a_9426_n851.n1 3.16959
R91 a_9426_n851.n2 a_9426_n851.n1 3.15795
R92 a_9426_n851.n1 a_9426_n851.n0 2.68725
R93 VDD.n13 VDD.n12 6857.65
R94 VDD.n15 VDD.n12 6857.65
R95 VDD.n15 VDD.n10 6857.65
R96 VDD.n13 VDD.n10 6857.65
R97 VDD.n44 VDD.n41 6130.59
R98 VDD.n46 VDD.n41 6130.59
R99 VDD.n44 VDD.n43 6130.59
R100 VDD.n46 VDD.n43 6130.59
R101 VDD.n4 VDD.n1 6130.59
R102 VDD.n6 VDD.n1 6130.59
R103 VDD.n4 VDD.n3 6130.59
R104 VDD.n6 VDD.n3 6130.59
R105 VDD.n17 VDD.n9 731.482
R106 VDD.n11 VDD.n9 731.482
R107 VDD.n16 VDD.n11 731.482
R108 VDD.n17 VDD.n16 731.482
R109 VDD.t50 VDD.t56 681.976
R110 VDD.t46 VDD.t50 681.976
R111 VDD.t48 VDD.t60 681.976
R112 VDD.t62 VDD.t48 681.976
R113 VDD.t54 VDD.t52 681.976
R114 VDD.t44 VDD.t54 681.976
R115 VDD.t58 VDD.t42 681.976
R116 VDD.t40 VDD.t58 681.976
R117 VDD.n48 VDD.n47 653.929
R118 VDD.n47 VDD.n42 653.929
R119 VDD.n42 VDD.n40 653.929
R120 VDD.n48 VDD.n40 653.929
R121 VDD.n8 VDD.n7 653.929
R122 VDD.n7 VDD.n2 653.929
R123 VDD.n2 VDD.n0 653.929
R124 VDD.n8 VDD.n0 653.929
R125 VDD.t56 VDD.n44 541.571
R126 VDD.n46 VDD.t62 541.571
R127 VDD.t52 VDD.n4 541.571
R128 VDD.n6 VDD.t40 541.571
R129 VDD.n45 VDD.t46 340.988
R130 VDD.t60 VDD.n45 340.988
R131 VDD.n5 VDD.t44 340.988
R132 VDD.t42 VDD.n5 340.988
R133 VDD.t36 VDD.n10 318.216
R134 VDD.t4 VDD.n12 318.216
R135 VDD.t6 VDD.t36 235.267
R136 VDD.t22 VDD.t6 235.267
R137 VDD.t34 VDD.t22 235.267
R138 VDD.t0 VDD.t34 235.267
R139 VDD.t12 VDD.t0 235.267
R140 VDD.t28 VDD.t12 235.267
R141 VDD.t14 VDD.t28 235.267
R142 VDD.t20 VDD.t14 235.267
R143 VDD.t32 VDD.t20 235.267
R144 VDD.t38 VDD.t8 235.267
R145 VDD.t8 VDD.t24 235.267
R146 VDD.t24 VDD.t10 235.267
R147 VDD.t10 VDD.t18 235.267
R148 VDD.t18 VDD.t30 235.267
R149 VDD.t30 VDD.t2 235.267
R150 VDD.t2 VDD.t16 235.267
R151 VDD.t16 VDD.t26 235.267
R152 VDD.t26 VDD.t4 235.267
R153 VDD.n55 VDD.n54 204.227
R154 VDD.n60 VDD.n59 204.191
R155 VDD.n58 VDD.n57 204.185
R156 VDD.n32 VDD.n31 201.939
R157 VDD.n23 VDD.n22 201.929
R158 VDD.n53 VDD.n52 201.869
R159 VDD.n39 VDD.n38 201.867
R160 VDD.n34 VDD.n28 201.861
R161 VDD.n26 VDD.n18 201.861
R162 VDD.n25 VDD.n19 201.861
R163 VDD.n51 VDD.n50 201.859
R164 VDD.n33 VDD.n29 201.858
R165 VDD.n24 VDD.n20 201.858
R166 VDD.n32 VDD.n30 201.855
R167 VDD.n35 VDD.n27 201.853
R168 VDD.n23 VDD.n21 201.852
R169 VDD.n14 VDD.t32 117.633
R170 VDD.n14 VDD.t38 117.633
R171 VDD.n47 VDD.n46 30.8338
R172 VDD.n44 VDD.n40 30.8338
R173 VDD.n12 VDD.n11 30.8338
R174 VDD.n17 VDD.n10 30.8338
R175 VDD.n7 VDD.n6 30.8338
R176 VDD.n4 VDD.n0 30.8338
R177 VDD.n59 VDD.t59 28.5655
R178 VDD.n59 VDD.t41 28.5655
R179 VDD.n57 VDD.t45 28.5655
R180 VDD.n57 VDD.t43 28.5655
R181 VDD.n54 VDD.t53 28.5655
R182 VDD.n54 VDD.t55 28.5655
R183 VDD.n50 VDD.t47 28.5655
R184 VDD.n50 VDD.t61 28.5655
R185 VDD.n38 VDD.t57 28.5655
R186 VDD.n38 VDD.t51 28.5655
R187 VDD.n52 VDD.t49 28.5655
R188 VDD.n52 VDD.t63 28.5655
R189 VDD.n31 VDD.t27 28.5655
R190 VDD.n31 VDD.t5 28.5655
R191 VDD.n30 VDD.t3 28.5655
R192 VDD.n30 VDD.t17 28.5655
R193 VDD.n29 VDD.t19 28.5655
R194 VDD.n29 VDD.t31 28.5655
R195 VDD.n28 VDD.t25 28.5655
R196 VDD.n28 VDD.t11 28.5655
R197 VDD.n27 VDD.t39 28.5655
R198 VDD.n27 VDD.t9 28.5655
R199 VDD.n18 VDD.t21 28.5655
R200 VDD.n18 VDD.t33 28.5655
R201 VDD.n19 VDD.t29 28.5655
R202 VDD.n19 VDD.t15 28.5655
R203 VDD.n20 VDD.t1 28.5655
R204 VDD.n20 VDD.t13 28.5655
R205 VDD.n21 VDD.t23 28.5655
R206 VDD.n21 VDD.t35 28.5655
R207 VDD.n22 VDD.t37 28.5655
R208 VDD.n22 VDD.t7 28.5655
R209 VDD.n43 VDD.n42 4.5127
R210 VDD.n45 VDD.n43 4.5127
R211 VDD.n48 VDD.n41 4.5127
R212 VDD.n45 VDD.n41 4.5127
R213 VDD.n3 VDD.n2 4.5127
R214 VDD.n5 VDD.n3 4.5127
R215 VDD.n8 VDD.n1 4.5127
R216 VDD.n5 VDD.n1 4.5127
R217 VDD.n13 VDD.n9 3.85467
R218 VDD.n14 VDD.n13 3.85467
R219 VDD.n16 VDD.n15 3.85467
R220 VDD.n15 VDD.n14 3.85467
R221 VDD.n37 VDD.n17 2.37291
R222 VDD VDD.n60 0.810764
R223 VDD.n39 VDD.n37 0.39218
R224 VDD.n49 VDD.n48 0.238962
R225 VDD.n56 VDD.n8 0.238962
R226 VDD.n55 VDD.n53 0.217543
R227 VDD.n56 VDD.n55 0.106715
R228 VDD.n60 VDD.n58 0.106599
R229 VDD.n53 VDD.n51 0.102732
R230 VDD.n49 VDD.n39 0.101393
R231 VDD.n35 VDD.n34 0.0727022
R232 VDD.n24 VDD.n23 0.0722509
R233 VDD.n26 VDD.n25 0.0722509
R234 VDD.n34 VDD.n33 0.0722509
R235 VDD.n25 VDD.n24 0.0713484
R236 VDD.n33 VDD.n32 0.0713484
R237 VDD.n36 VDD.n26 0.0492365
R238 VDD.n37 VDD.n36 0.0353837
R239 VDD.n36 VDD.n35 0.0221607
R240 VDD.n58 VDD.n56 0.000963822
R241 VDD.n51 VDD.n49 0.000723214
R242 VOUT.n4 VOUT.t16 230.594
R243 VOUT.n13 VOUT.t2 230.565
R244 VOUT.n4 VOUT.n3 201.864
R245 VOUT.n7 VOUT.n0 201.857
R246 VOUT.n16 VOUT.n9 201.857
R247 VOUT.n15 VOUT.n10 201.857
R248 VOUT.n17 VOUT.n8 201.857
R249 VOUT.n13 VOUT.n12 201.857
R250 VOUT.n5 VOUT.n2 201.855
R251 VOUT.n6 VOUT.n1 201.855
R252 VOUT.n14 VOUT.n11 201.855
R253 VOUT.n21 VOUT.t24 86.4014
R254 VOUT.n24 VOUT.n23 68.9752
R255 VOUT.n24 VOUT.n22 68.355
R256 VOUT.n21 VOUT.n20 68.3524
R257 VOUT.n3 VOUT.t3 28.5655
R258 VOUT.n3 VOUT.t11 28.5655
R259 VOUT.n2 VOUT.t14 28.5655
R260 VOUT.n2 VOUT.t0 28.5655
R261 VOUT.n1 VOUT.t6 28.5655
R262 VOUT.n1 VOUT.t15 28.5655
R263 VOUT.n0 VOUT.t7 28.5655
R264 VOUT.n0 VOUT.t10 28.5655
R265 VOUT.n8 VOUT.t13 28.5655
R266 VOUT.n8 VOUT.t18 28.5655
R267 VOUT.n9 VOUT.t4 28.5655
R268 VOUT.n9 VOUT.t19 28.5655
R269 VOUT.n10 VOUT.t5 28.5655
R270 VOUT.n10 VOUT.t9 28.5655
R271 VOUT.n11 VOUT.t12 28.5655
R272 VOUT.n11 VOUT.t1 28.5655
R273 VOUT.n12 VOUT.t8 28.5655
R274 VOUT.n12 VOUT.t17 28.5655
R275 VOUT.n23 VOUT.t20 17.4005
R276 VOUT.n23 VOUT.t21 17.4005
R277 VOUT.n22 VOUT.t25 17.4005
R278 VOUT.n22 VOUT.t22 17.4005
R279 VOUT.n20 VOUT.t26 17.4005
R280 VOUT.n20 VOUT.t23 17.4005
R281 VOUT.n26 VOUT.n25 0.798123
R282 VOUT.n19 VOUT.n18 0.546565
R283 VOUT.n25 VOUT.n21 0.298332
R284 VOUT.n25 VOUT.n24 0.283026
R285 VOUT.n6 VOUT.n5 0.129532
R286 VOUT.n15 VOUT.n14 0.129532
R287 VOUT.n7 VOUT.n6 0.127919
R288 VOUT.n5 VOUT.n4 0.127113
R289 VOUT.n17 VOUT.n16 0.127113
R290 VOUT.n16 VOUT.n15 0.127113
R291 VOUT.n14 VOUT.n13 0.127113
R292 VOUT VOUT.n19 0.124047
R293 VOUT VOUT.n19 0.115989
R294 VOUT.n19 VOUT 0.108552
R295 VOUT.n18 VOUT.n7 0.0855806
R296 VOUT.n26 VOUT 0.0767338
R297 VOUT VOUT.n26 0.0746279
R298 VOUT.n18 VOUT.n17 0.0420323
R299 VX.n0 VX.t2 84.9941
R300 VX.n0 VX.t3 83.7178
R301 VX.n0 VX.n1 66.9929
R302 VX VX.t1 37.4299
R303 VX.n0 VX.t0 34.9733
R304 VX.n1 VX.t5 17.4005
R305 VX.n1 VX.t4 17.4005
R306 VX VX.n0 3.89792
R307 VSS.n33 VSS.n32 365574
R308 VSS.n33 VSS.n16 14086.5
R309 VSS.n62 VSS.n16 13436.2
R310 VSS.n49 VSS.n30 11339.1
R311 VSS.n50 VSS.n30 11339.1
R312 VSS.n49 VSS.n31 11339.1
R313 VSS.n50 VSS.n31 11339.1
R314 VSS.n46 VSS.n33 9866.67
R315 VSS.n38 VSS.n16 8581.37
R316 VSS.n64 VSS.n4 7358.53
R317 VSS.n78 VSS.n4 7358.53
R318 VSS.n64 VSS.n5 7358.53
R319 VSS.n78 VSS.n5 7358.53
R320 VSS.n59 VSS.n15 7358.53
R321 VSS.n59 VSS.n13 7358.53
R322 VSS.n67 VSS.n15 7358.53
R323 VSS.n67 VSS.n13 7358.53
R324 VSS.n81 VSS.n3 5446.47
R325 VSS.n86 VSS.n3 5446.47
R326 VSS.n84 VSS.n81 5446.47
R327 VSS.n36 VSS.n17 3377.97
R328 VSS.n57 VSS.n17 3377.97
R329 VSS.n36 VSS.n18 3377.97
R330 VSS.n57 VSS.n18 3377.97
R331 VSS.n44 VSS.n34 3377.97
R332 VSS.n40 VSS.n34 3377.97
R333 VSS.n44 VSS.n35 3377.97
R334 VSS.n40 VSS.n35 3377.97
R335 VSS.n39 VSS.n38 2986.36
R336 VSS.n46 VSS.n45 2416.93
R337 VSS.n38 VSS.n37 2260.52
R338 VSS.t13 VSS.t19 843.886
R339 VSS.t19 VSS.t3 843.886
R340 VSS.t5 VSS.t3 843.886
R341 VSS.t5 VSS.t7 843.886
R342 VSS.t7 VSS.t9 843.886
R343 VSS.t9 VSS.t11 843.886
R344 VSS.t31 VSS.t27 831.354
R345 VSS.n60 VSS.n58 784.159
R346 VSS.n48 VSS.n28 736.754
R347 VSS.n51 VSS.n28 736.754
R348 VSS.n48 VSS.n29 736.754
R349 VSS.n51 VSS.n29 736.754
R350 VSS.n32 VSS.t13 631.994
R351 VSS.t11 VSS.n47 631.819
R352 VSS.t27 VSS.n60 622.607
R353 VSS.t25 VSS.t21 488.652
R354 VSS.t29 VSS.t15 488.652
R355 VSS.t23 VSS.t17 488.652
R356 VSS.n14 VSS.n12 478.118
R357 VSS.n69 VSS.n12 478.118
R358 VSS.n68 VSS.n14 478.118
R359 VSS.n69 VSS.n68 478.118
R360 VSS.n7 VSS.n6 478.118
R361 VSS.n76 VSS.n7 478.118
R362 VSS.n77 VSS.n6 478.118
R363 VSS.n77 VSS.n76 478.118
R364 VSS.n80 VSS.n79 452.377
R365 VSS.n61 VSS.t31 415.678
R366 VSS.n66 VSS.n65 390.495
R367 VSS.n66 VSS.t25 365.955
R368 VSS.n65 VSS.t29 365.955
R369 VSS.n79 VSS.t17 365.955
R370 VSS.n37 VSS.t0 350.33
R371 VSS.n58 VSS.t0 350.33
R372 VSS.n45 VSS.t1 348.892
R373 VSS.n39 VSS.t1 348.892
R374 VSS.n82 VSS.n1 342.51
R375 VSS.n88 VSS.n87 341.447
R376 VSS.n83 VSS.n82 333.476
R377 VSS.n87 VSS.n2 329.12
R378 VSS.n84 VSS.n83 292.5
R379 VSS.n3 VSS.n1 292.5
R380 VSS.t2 VSS.n3 292.5
R381 VSS.n62 VSS.n61 270.462
R382 VSS.n85 VSS.n84 268.889
R383 VSS.t15 VSS.n63 244.327
R384 VSS.n63 VSS.t23 244.327
R385 VSS.n47 VSS.n46 229.582
R386 VSS.n42 VSS.n41 219.482
R387 VSS.n43 VSS.n42 219.482
R388 VSS.n20 VSS.n19 219.482
R389 VSS.n55 VSS.n20 219.482
R390 VSS.n56 VSS.n19 219.482
R391 VSS.n56 VSS.n55 219.482
R392 VSS.n41 VSS.n21 197.23
R393 VSS.n43 VSS.n21 197.23
R394 VSS.n35 VSS.n21 195
R395 VSS.n35 VSS.t1 195
R396 VSS.n42 VSS.n34 195
R397 VSS.n34 VSS.t1 195
R398 VSS.n55 VSS.n18 195
R399 VSS.n18 VSS.t0 195
R400 VSS.n19 VSS.n17 195
R401 VSS.n17 VSS.t0 195
R402 VSS.n86 VSS.n85 170.768
R403 VSS.n80 VSS.t2 157.905
R404 VSS.n30 VSS.n28 117.001
R405 VSS.n32 VSS.n30 117.001
R406 VSS.n31 VSS.n29 117.001
R407 VSS.n47 VSS.n31 117.001
R408 VSS.n59 VSS.n12 117.001
R409 VSS.n60 VSS.n59 117.001
R410 VSS.n78 VSS.n77 117.001
R411 VSS.n79 VSS.n78 117.001
R412 VSS.n64 VSS.n7 117.001
R413 VSS.n65 VSS.n64 117.001
R414 VSS.n68 VSS.n67 117.001
R415 VSS.n67 VSS.n66 117.001
R416 VSS.n26 VSS.t12 86.7617
R417 VSS.n24 VSS.n23 69.3536
R418 VSS.n24 VSS.n22 68.8088
R419 VSS.n26 VSS.n25 68.8088
R420 VSS.n72 VSS.n71 68.5048
R421 VSS.n74 VSS.n73 68.5002
R422 VSS.n10 VSS.n9 67.0731
R423 VSS.n10 VSS.n8 67.0703
R424 VSS.n41 VSS.n40 58.5005
R425 VSS.n40 VSS.n39 58.5005
R426 VSS.n44 VSS.n43 58.5005
R427 VSS.n45 VSS.n44 58.5005
R428 VSS.n57 VSS.n56 58.5005
R429 VSS.n58 VSS.n57 58.5005
R430 VSS.n36 VSS.n20 58.5005
R431 VSS.n37 VSS.n36 58.5005
R432 VSS.t21 VSS.n62 53.7574
R433 VSS.n87 VSS.n86 27.8576
R434 VSS.n82 VSS.n81 27.8576
R435 VSS.n81 VSS.n80 27.8576
R436 VSS.n69 VSS.n13 20.8934
R437 VSS.n61 VSS.n13 20.8934
R438 VSS.n15 VSS.n14 20.8934
R439 VSS.n61 VSS.n15 20.8934
R440 VSS.n76 VSS.n5 20.8934
R441 VSS.n63 VSS.n5 20.8934
R442 VSS.n6 VSS.n4 20.8934
R443 VSS.n63 VSS.n4 20.8934
R444 VSS.n23 VSS.t14 17.4005
R445 VSS.n23 VSS.t20 17.4005
R446 VSS.n22 VSS.t4 17.4005
R447 VSS.n22 VSS.t6 17.4005
R448 VSS.n25 VSS.t8 17.4005
R449 VSS.n25 VSS.t10 17.4005
R450 VSS.n9 VSS.t22 17.4005
R451 VSS.n9 VSS.t26 17.4005
R452 VSS.n8 VSS.t28 17.4005
R453 VSS.n8 VSS.t32 17.4005
R454 VSS.n73 VSS.t24 17.4005
R455 VSS.n73 VSS.t18 17.4005
R456 VSS.n71 VSS.t30 17.4005
R457 VSS.n71 VSS.t16 17.4005
R458 VSS.n51 VSS.n50 12.188
R459 VSS.n50 VSS.t5 12.188
R460 VSS.n49 VSS.n48 12.188
R461 VSS.t5 VSS.n49 12.188
R462 VSS.n85 VSS.t2 9.17195
R463 VSS VSS.n88 6.41514
R464 VSS.n54 VSS.n11 3.71217
R465 VSS.n2 VSS.n0 3.32603
R466 VSS.n53 VSS.n21 3.14022
R467 VSS.n55 VSS.n54 3.13594
R468 VSS.n72 VSS.n70 2.61112
R469 VSS.n83 VSS.n2 0.914786
R470 VSS.n54 VSS.n53 0.586639
R471 VSS.n53 VSS.n52 0.510493
R472 VSS.n88 VSS.n1 0.441879
R473 VSS.n27 VSS.n26 0.415163
R474 VSS.n76 VSS.n75 0.358192
R475 VSS.n70 VSS.n69 0.358192
R476 VSS.n52 VSS.n51 0.202674
R477 VSS.n74 VSS.n0 0.186816
R478 VSS.n27 VSS.n24 0.137519
R479 VSS.n11 VSS.n10 0.0838333
R480 VSS.n75 VSS.n72 0.0687353
R481 VSS.n75 VSS.n74 0.0684412
R482 VSS VSS.n0 0.0363166
R483 VSS.n52 VSS.n27 0.0301526
R484 VSS.n70 VSS.n11 0.000862669
R485 MINUS MINUS.t0 155.806
R486 PLUS.n0 PLUS.t0 156.07
R487 PLUS.n0 PLUS 0.231981
R488 PLUS PLUS.n0 0.0861164
C0 VDD VBIAS 0.335706f
C1 PLUS VX 0.554937f
C2 PLUS MINUS 0.006311f
C3 VOUT VBIAS 1.93193f
C4 VX VBIAS 2.94391f
C5 VBIAS MINUS 0.002585f
C6 VOUT VDD 4.97876f
C7 VDD VX 0.025529f
C8 VDD MINUS 4.98e-19
C9 PLUS VBIAS 0.188144f
C10 PLUS VDD 2.92e-19
C11 VX MINUS 0.396729f
.ends


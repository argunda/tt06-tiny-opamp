VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_argunda_tiny_opamp
  CLASS BLOCK ;
  FOREIGN tt_um_argunda_tiny_opamp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.350000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.350000 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3417.542725 ;
    ANTENNADIFFAREA 662.595642 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 158.080 5.000 159.580 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 10.930 212.215 150.690 213.820 ;
      LAYER pwell ;
        RECT 11.125 211.015 12.495 211.825 ;
        RECT 12.505 211.015 18.015 211.825 ;
        RECT 18.025 211.015 23.535 211.825 ;
        RECT 24.015 211.100 24.445 211.885 ;
        RECT 24.465 211.015 29.975 211.825 ;
        RECT 29.985 211.015 35.495 211.825 ;
        RECT 35.505 211.015 36.875 211.825 ;
        RECT 36.895 211.100 37.325 211.885 ;
        RECT 37.345 211.015 42.855 211.825 ;
        RECT 42.865 211.015 48.375 211.825 ;
        RECT 48.385 211.015 49.755 211.825 ;
        RECT 49.775 211.100 50.205 211.885 ;
        RECT 50.225 211.015 55.735 211.825 ;
        RECT 55.745 211.015 61.255 211.825 ;
        RECT 61.265 211.015 62.635 211.825 ;
        RECT 62.655 211.100 63.085 211.885 ;
        RECT 64.510 211.695 65.855 211.925 ;
        RECT 64.025 211.015 65.855 211.695 ;
        RECT 65.865 211.015 71.375 211.825 ;
        RECT 71.385 211.015 75.055 211.825 ;
        RECT 75.535 211.100 75.965 211.885 ;
        RECT 75.985 211.015 81.495 211.825 ;
        RECT 81.505 211.015 85.175 211.825 ;
        RECT 85.185 211.015 86.555 211.825 ;
        RECT 86.565 211.015 87.935 211.795 ;
        RECT 88.415 211.100 88.845 211.885 ;
        RECT 88.865 211.015 94.375 211.825 ;
        RECT 94.385 211.015 96.215 211.825 ;
        RECT 96.225 211.015 97.595 211.795 ;
        RECT 97.605 211.015 101.275 211.825 ;
        RECT 101.295 211.100 101.725 211.885 ;
        RECT 101.745 211.015 104.495 211.825 ;
        RECT 107.160 211.695 108.080 211.925 ;
        RECT 104.615 211.015 108.080 211.695 ;
        RECT 108.195 211.015 109.545 211.925 ;
        RECT 109.565 211.015 110.935 211.795 ;
        RECT 110.945 211.015 113.695 211.825 ;
        RECT 114.175 211.100 114.605 211.885 ;
        RECT 114.625 211.015 116.455 211.825 ;
        RECT 116.465 211.015 117.835 211.795 ;
        RECT 117.845 211.015 123.355 211.825 ;
        RECT 123.365 211.015 127.035 211.825 ;
        RECT 127.055 211.100 127.485 211.885 ;
        RECT 127.505 211.015 128.875 211.795 ;
        RECT 128.885 211.015 134.395 211.825 ;
        RECT 134.405 211.015 136.235 211.825 ;
        RECT 136.705 211.015 139.445 211.695 ;
        RECT 139.935 211.100 140.365 211.885 ;
        RECT 140.385 211.015 145.895 211.825 ;
        RECT 145.905 211.015 148.655 211.825 ;
        RECT 149.125 211.015 150.495 211.825 ;
        RECT 11.265 210.805 11.435 211.015 ;
        RECT 12.645 210.805 12.815 211.015 ;
        RECT 17.705 210.805 17.875 210.995 ;
        RECT 18.165 210.805 18.335 211.015 ;
        RECT 20.005 210.805 20.175 210.995 ;
        RECT 23.680 210.855 23.800 210.965 ;
        RECT 24.605 210.825 24.775 211.015 ;
        RECT 29.665 210.805 29.835 210.995 ;
        RECT 30.125 210.965 30.295 211.015 ;
        RECT 30.120 210.855 30.295 210.965 ;
        RECT 30.125 210.825 30.295 210.855 ;
        RECT 32.425 210.825 32.595 210.995 ;
        RECT 32.425 210.805 32.590 210.825 ;
        RECT 33.810 210.805 33.980 210.995 ;
        RECT 35.645 210.825 35.815 211.015 ;
        RECT 36.565 210.805 36.735 210.995 ;
        RECT 37.485 210.825 37.655 211.015 ;
        RECT 38.405 210.805 38.575 210.995 ;
        RECT 38.860 210.855 38.980 210.965 ;
        RECT 39.325 210.805 39.495 210.995 ;
        RECT 43.005 210.825 43.175 211.015 ;
        RECT 44.845 210.805 45.015 210.995 ;
        RECT 45.305 210.805 45.475 210.995 ;
        RECT 48.525 210.805 48.695 211.015 ;
        RECT 50.365 210.825 50.535 211.015 ;
        RECT 51.740 210.855 51.860 210.965 ;
        RECT 52.205 210.805 52.375 210.995 ;
        RECT 55.425 210.805 55.595 210.995 ;
        RECT 55.885 210.825 56.055 211.015 ;
        RECT 61.405 210.825 61.575 211.015 ;
        RECT 63.255 210.850 63.415 210.970 ;
        RECT 64.165 210.805 64.335 211.015 ;
        RECT 66.005 210.825 66.175 211.015 ;
        RECT 71.525 210.805 71.695 211.015 ;
        RECT 74.285 210.805 74.455 210.995 ;
        RECT 75.200 210.855 75.320 210.965 ;
        RECT 76.125 210.825 76.295 211.015 ;
        RECT 81.645 210.995 81.815 211.015 ;
        RECT 81.645 210.825 81.820 210.995 ;
        RECT 11.125 209.995 12.495 210.805 ;
        RECT 12.505 209.995 15.255 210.805 ;
        RECT 15.275 210.125 18.015 210.805 ;
        RECT 18.025 209.995 19.855 210.805 ;
        RECT 19.865 210.125 27.175 210.805 ;
        RECT 27.235 210.125 29.975 210.805 ;
        RECT 30.755 210.125 32.590 210.805 ;
        RECT 23.380 209.905 24.290 210.125 ;
        RECT 25.825 209.895 27.175 210.125 ;
        RECT 30.755 209.895 31.685 210.125 ;
        RECT 32.745 209.895 34.095 210.805 ;
        RECT 34.135 210.125 36.875 210.805 ;
        RECT 36.895 209.935 37.325 210.720 ;
        RECT 37.345 210.025 38.715 210.805 ;
        RECT 39.285 209.895 42.395 210.805 ;
        RECT 42.415 210.125 45.155 210.805 ;
        RECT 45.265 209.895 48.375 210.805 ;
        RECT 48.425 209.895 51.595 210.805 ;
        RECT 52.165 209.895 55.275 210.805 ;
        RECT 55.285 210.125 62.595 210.805 ;
        RECT 58.800 209.905 59.710 210.125 ;
        RECT 61.245 209.895 62.595 210.125 ;
        RECT 62.655 209.935 63.085 210.720 ;
        RECT 64.025 210.125 71.335 210.805 ;
        RECT 71.385 210.125 74.125 210.805 ;
        RECT 74.145 210.125 81.455 210.805 ;
        RECT 81.650 210.775 81.820 210.825 ;
        RECT 84.865 210.805 85.035 210.995 ;
        RECT 85.325 210.825 85.495 211.015 ;
        RECT 86.705 210.825 86.875 211.015 ;
        RECT 87.635 210.850 87.795 210.960 ;
        RECT 88.080 210.855 88.200 210.965 ;
        RECT 89.005 210.805 89.175 211.015 ;
        RECT 94.525 210.825 94.695 211.015 ;
        RECT 96.365 210.825 96.535 211.015 ;
        RECT 96.825 210.805 96.995 210.995 ;
        RECT 97.745 210.825 97.915 211.015 ;
        RECT 101.885 210.825 102.055 211.015 ;
        RECT 104.185 210.805 104.355 210.995 ;
        RECT 104.645 210.825 104.815 211.015 ;
        RECT 109.245 210.825 109.415 211.015 ;
        RECT 110.625 210.825 110.795 211.015 ;
        RECT 111.085 210.825 111.255 211.015 ;
        RECT 111.545 210.805 111.715 210.995 ;
        RECT 113.845 210.965 114.015 210.995 ;
        RECT 113.840 210.855 114.015 210.965 ;
        RECT 113.845 210.805 114.015 210.855 ;
        RECT 114.765 210.825 114.935 211.015 ;
        RECT 117.525 210.825 117.695 211.015 ;
        RECT 117.985 210.825 118.155 211.015 ;
        RECT 123.045 210.805 123.215 210.995 ;
        RECT 123.505 210.805 123.675 211.015 ;
        RECT 128.565 210.825 128.735 211.015 ;
        RECT 129.025 210.825 129.195 211.015 ;
        RECT 130.865 210.805 131.035 210.995 ;
        RECT 134.545 210.825 134.715 211.015 ;
        RECT 136.385 210.965 136.555 210.995 ;
        RECT 136.380 210.855 136.555 210.965 ;
        RECT 136.385 210.805 136.555 210.855 ;
        RECT 136.845 210.825 137.015 211.015 ;
        RECT 139.600 210.855 139.720 210.965 ;
        RECT 140.525 210.805 140.695 211.015 ;
        RECT 146.045 210.805 146.215 211.015 ;
        RECT 148.800 210.855 148.920 210.965 ;
        RECT 150.185 210.805 150.355 211.015 ;
        RECT 83.780 210.775 84.715 210.805 ;
        RECT 81.650 210.575 84.715 210.775 ;
        RECT 67.540 209.905 68.450 210.125 ;
        RECT 69.985 209.895 71.335 210.125 ;
        RECT 77.660 209.905 78.570 210.125 ;
        RECT 80.105 209.895 81.455 210.125 ;
        RECT 81.505 210.095 84.715 210.575 ;
        RECT 84.725 210.125 87.465 210.805 ;
        RECT 81.505 209.895 82.435 210.095 ;
        RECT 83.765 209.895 84.715 210.095 ;
        RECT 88.415 209.935 88.845 210.720 ;
        RECT 88.865 210.125 96.595 210.805 ;
        RECT 96.685 210.125 103.995 210.805 ;
        RECT 104.045 210.125 111.355 210.805 ;
        RECT 92.380 209.905 93.290 210.125 ;
        RECT 94.825 209.895 96.595 210.125 ;
        RECT 100.200 209.905 101.110 210.125 ;
        RECT 102.645 209.895 103.995 210.125 ;
        RECT 107.560 209.905 108.470 210.125 ;
        RECT 110.005 209.895 111.355 210.125 ;
        RECT 111.415 209.895 112.765 210.805 ;
        RECT 112.795 209.895 114.145 210.805 ;
        RECT 114.175 209.935 114.605 210.720 ;
        RECT 115.625 210.125 123.355 210.805 ;
        RECT 123.365 210.125 130.675 210.805 ;
        RECT 115.625 209.895 117.395 210.125 ;
        RECT 118.930 209.905 119.840 210.125 ;
        RECT 126.880 209.905 127.790 210.125 ;
        RECT 129.325 209.895 130.675 210.125 ;
        RECT 130.725 209.995 136.235 210.805 ;
        RECT 136.245 209.995 139.915 210.805 ;
        RECT 139.935 209.935 140.365 210.720 ;
        RECT 140.385 209.995 145.895 210.805 ;
        RECT 145.905 209.995 148.655 210.805 ;
        RECT 149.125 209.995 150.495 210.805 ;
      LAYER nwell ;
        RECT 10.930 206.775 150.690 209.605 ;
      LAYER pwell ;
        RECT 11.125 205.575 12.495 206.385 ;
        RECT 12.505 205.575 18.015 206.385 ;
        RECT 18.025 205.575 21.695 206.385 ;
        RECT 22.165 205.575 23.535 206.355 ;
        RECT 24.015 205.660 24.445 206.445 ;
        RECT 24.465 206.285 25.415 206.485 ;
        RECT 26.745 206.285 27.675 206.485 ;
        RECT 24.465 205.805 27.675 206.285 ;
        RECT 24.465 205.605 27.530 205.805 ;
        RECT 24.465 205.575 25.400 205.605 ;
        RECT 11.265 205.365 11.435 205.575 ;
        RECT 12.645 205.365 12.815 205.575 ;
        RECT 18.165 205.365 18.335 205.575 ;
        RECT 21.840 205.415 21.960 205.525 ;
        RECT 23.225 205.385 23.395 205.575 ;
        RECT 23.685 205.525 23.855 205.555 ;
        RECT 23.680 205.415 23.855 205.525 ;
        RECT 23.685 205.365 23.855 205.415 ;
        RECT 27.360 205.385 27.530 205.605 ;
        RECT 27.695 205.575 30.425 206.485 ;
        RECT 30.445 205.575 32.275 206.385 ;
        RECT 32.365 206.255 34.135 206.485 ;
        RECT 35.670 206.255 36.580 206.475 ;
        RECT 32.365 205.575 40.095 206.255 ;
        RECT 40.105 205.575 43.775 206.385 ;
        RECT 43.785 205.575 45.155 206.385 ;
        RECT 46.985 206.255 47.915 206.485 ;
        RECT 45.165 205.575 47.915 206.255 ;
        RECT 47.925 205.575 49.755 206.385 ;
        RECT 49.775 205.660 50.205 206.445 ;
        RECT 50.225 205.575 52.055 206.385 ;
        RECT 52.550 206.255 53.895 206.485 ;
        RECT 52.065 205.575 53.895 206.255 ;
        RECT 53.905 205.575 59.415 206.385 ;
        RECT 59.425 205.575 63.095 206.385 ;
        RECT 63.105 205.575 64.475 206.385 ;
        RECT 66.290 206.285 67.235 206.485 ;
        RECT 64.485 205.605 67.235 206.285 ;
        RECT 69.320 206.255 70.455 206.485 ;
        RECT 27.825 205.385 27.995 205.575 ;
        RECT 29.215 205.410 29.375 205.520 ;
        RECT 30.125 205.365 30.295 205.555 ;
        RECT 30.585 205.385 30.755 205.575 ;
        RECT 32.425 205.365 32.595 205.555 ;
        RECT 36.115 205.410 36.275 205.520 ;
        RECT 37.485 205.365 37.655 205.555 ;
        RECT 39.785 205.385 39.955 205.575 ;
        RECT 40.245 205.385 40.415 205.575 ;
        RECT 41.165 205.365 41.335 205.555 ;
        RECT 41.625 205.365 41.795 205.555 ;
        RECT 43.925 205.385 44.095 205.575 ;
        RECT 44.380 205.415 44.500 205.525 ;
        RECT 44.850 205.365 45.020 205.555 ;
        RECT 45.305 205.385 45.475 205.575 ;
        RECT 48.065 205.555 48.235 205.575 ;
        RECT 46.225 205.365 46.395 205.555 ;
        RECT 48.060 205.385 48.235 205.555 ;
        RECT 48.060 205.365 48.230 205.385 ;
        RECT 49.445 205.365 49.615 205.555 ;
        RECT 50.365 205.385 50.535 205.575 ;
        RECT 52.205 205.385 52.375 205.575 ;
        RECT 53.135 205.410 53.295 205.520 ;
        RECT 54.045 205.365 54.215 205.575 ;
        RECT 57.260 205.415 57.380 205.525 ;
        RECT 57.725 205.365 57.895 205.555 ;
        RECT 59.565 205.385 59.735 205.575 ;
        RECT 60.945 205.365 61.115 205.555 ;
        RECT 63.245 205.365 63.415 205.575 ;
        RECT 64.630 205.385 64.800 205.605 ;
        RECT 66.290 205.575 67.235 205.605 ;
        RECT 67.245 205.575 70.455 206.255 ;
        RECT 70.660 205.575 74.135 206.485 ;
        RECT 74.145 205.575 75.515 206.385 ;
        RECT 75.535 205.660 75.965 206.445 ;
        RECT 75.985 205.575 81.495 206.385 ;
        RECT 82.555 206.255 83.485 206.485 ;
        RECT 81.650 205.575 83.485 206.255 ;
        RECT 83.825 205.575 85.175 206.485 ;
        RECT 88.700 206.255 89.610 206.475 ;
        RECT 91.145 206.255 92.915 206.485 ;
        RECT 85.185 205.575 92.915 206.255 ;
        RECT 93.100 206.255 94.020 206.485 ;
        RECT 98.090 206.255 99.435 206.485 ;
        RECT 93.100 205.575 96.565 206.255 ;
        RECT 97.605 205.575 99.435 206.255 ;
        RECT 99.455 205.575 100.805 206.485 ;
        RECT 101.295 205.660 101.725 206.445 ;
        RECT 101.745 205.575 103.575 206.385 ;
        RECT 107.100 206.255 108.010 206.475 ;
        RECT 109.545 206.255 110.895 206.485 ;
        RECT 114.920 206.255 115.830 206.475 ;
        RECT 117.365 206.255 118.715 206.485 ;
        RECT 103.585 205.575 110.895 206.255 ;
        RECT 111.405 205.575 118.715 206.255 ;
        RECT 118.765 205.575 120.135 206.385 ;
        RECT 122.800 206.255 123.720 206.485 ;
        RECT 120.255 205.575 123.720 206.255 ;
        RECT 123.835 205.575 125.185 206.485 ;
        RECT 125.205 205.575 127.035 206.385 ;
        RECT 127.055 205.660 127.485 206.445 ;
        RECT 127.505 205.575 129.335 206.385 ;
        RECT 129.900 206.255 130.820 206.485 ;
        RECT 129.900 205.575 133.365 206.255 ;
        RECT 133.485 205.575 138.995 206.385 ;
        RECT 139.005 205.575 144.515 206.385 ;
        RECT 144.525 205.575 148.195 206.385 ;
        RECT 149.125 205.575 150.495 206.385 ;
        RECT 67.385 205.385 67.555 205.575 ;
        RECT 68.760 205.415 68.880 205.525 ;
        RECT 69.225 205.365 69.395 205.555 ;
        RECT 72.445 205.365 72.615 205.555 ;
        RECT 73.820 205.385 73.990 205.575 ;
        RECT 74.285 205.385 74.455 205.575 ;
        RECT 76.125 205.365 76.295 205.575 ;
        RECT 81.650 205.555 81.815 205.575 ;
        RECT 77.505 205.365 77.675 205.555 ;
        RECT 79.800 205.415 79.920 205.525 ;
        RECT 80.265 205.385 80.435 205.555 ;
        RECT 81.645 205.385 81.815 205.555 ;
        RECT 80.285 205.365 80.435 205.385 ;
        RECT 83.940 205.365 84.110 205.555 ;
        RECT 84.405 205.365 84.575 205.555 ;
        RECT 84.860 205.385 85.030 205.575 ;
        RECT 85.325 205.385 85.495 205.575 ;
        RECT 88.080 205.415 88.200 205.525 ;
        RECT 89.005 205.365 89.175 205.555 ;
        RECT 90.845 205.365 91.015 205.555 ;
        RECT 96.365 205.385 96.535 205.575 ;
        RECT 96.835 205.420 96.995 205.530 ;
        RECT 97.745 205.385 97.915 205.575 ;
        RECT 98.665 205.365 98.835 205.555 ;
        RECT 99.585 205.385 99.755 205.575 ;
        RECT 100.960 205.415 101.080 205.525 ;
        RECT 101.885 205.385 102.055 205.575 ;
        RECT 103.725 205.385 103.895 205.575 ;
        RECT 104.185 205.365 104.355 205.555 ;
        RECT 111.080 205.415 111.200 205.525 ;
        RECT 111.545 205.385 111.715 205.575 ;
        RECT 113.845 205.365 114.015 205.555 ;
        RECT 114.765 205.365 114.935 205.555 ;
        RECT 118.905 205.385 119.075 205.575 ;
        RECT 120.285 205.365 120.455 205.575 ;
        RECT 124.885 205.385 125.055 205.575 ;
        RECT 125.345 205.385 125.515 205.575 ;
        RECT 125.805 205.365 125.975 205.555 ;
        RECT 127.645 205.385 127.815 205.575 ;
        RECT 129.480 205.415 129.600 205.525 ;
        RECT 131.325 205.365 131.495 205.555 ;
        RECT 133.165 205.385 133.335 205.575 ;
        RECT 133.625 205.385 133.795 205.575 ;
        RECT 136.845 205.365 137.015 205.555 ;
        RECT 139.145 205.385 139.315 205.575 ;
        RECT 139.600 205.415 139.720 205.525 ;
        RECT 140.525 205.365 140.695 205.555 ;
        RECT 144.665 205.385 144.835 205.575 ;
        RECT 146.045 205.365 146.215 205.555 ;
        RECT 148.355 205.420 148.515 205.530 ;
        RECT 148.800 205.415 148.920 205.525 ;
        RECT 150.185 205.365 150.355 205.575 ;
        RECT 11.125 204.555 12.495 205.365 ;
        RECT 12.505 204.555 18.015 205.365 ;
        RECT 18.025 204.555 23.535 205.365 ;
        RECT 23.545 204.555 29.055 205.365 ;
        RECT 29.985 204.685 32.275 205.365 ;
        RECT 31.355 204.455 32.275 204.685 ;
        RECT 32.285 204.555 35.955 205.365 ;
        RECT 36.895 204.495 37.325 205.280 ;
        RECT 37.345 204.555 38.715 205.365 ;
        RECT 38.725 204.685 41.475 205.365 ;
        RECT 38.725 204.455 39.655 204.685 ;
        RECT 41.485 204.555 44.235 205.365 ;
        RECT 44.705 204.455 46.055 205.365 ;
        RECT 46.100 204.455 47.915 205.365 ;
        RECT 47.945 204.455 49.295 205.365 ;
        RECT 49.305 204.555 52.975 205.365 ;
        RECT 54.005 204.455 57.115 205.365 ;
        RECT 57.685 204.455 60.795 205.365 ;
        RECT 60.805 204.555 62.635 205.365 ;
        RECT 62.655 204.495 63.085 205.280 ;
        RECT 63.105 204.555 68.615 205.365 ;
        RECT 69.085 204.455 72.295 205.365 ;
        RECT 72.305 204.555 75.975 205.365 ;
        RECT 75.985 204.555 77.355 205.365 ;
        RECT 77.365 204.685 79.655 205.365 ;
        RECT 78.735 204.455 79.655 204.685 ;
        RECT 80.285 204.545 82.215 205.365 ;
        RECT 81.265 204.455 82.215 204.545 ;
        RECT 82.425 204.455 84.255 205.365 ;
        RECT 84.265 204.555 87.935 205.365 ;
        RECT 88.415 204.495 88.845 205.280 ;
        RECT 88.865 204.555 90.695 205.365 ;
        RECT 90.705 204.685 98.435 205.365 ;
        RECT 94.220 204.465 95.130 204.685 ;
        RECT 96.665 204.455 98.435 204.685 ;
        RECT 98.525 204.555 104.035 205.365 ;
        RECT 104.045 204.555 106.795 205.365 ;
        RECT 106.845 204.685 114.155 205.365 ;
        RECT 106.845 204.455 108.195 204.685 ;
        RECT 109.730 204.465 110.640 204.685 ;
        RECT 114.175 204.495 114.605 205.280 ;
        RECT 114.625 204.555 120.135 205.365 ;
        RECT 120.145 204.555 125.655 205.365 ;
        RECT 125.665 204.555 131.175 205.365 ;
        RECT 131.185 204.555 136.695 205.365 ;
        RECT 136.705 204.555 139.455 205.365 ;
        RECT 139.935 204.495 140.365 205.280 ;
        RECT 140.385 204.555 145.895 205.365 ;
        RECT 145.905 204.555 148.655 205.365 ;
        RECT 149.125 204.555 150.495 205.365 ;
      LAYER nwell ;
        RECT 10.930 201.335 150.690 204.165 ;
      LAYER pwell ;
        RECT 11.125 200.135 12.495 200.945 ;
        RECT 12.505 200.135 16.175 200.945 ;
        RECT 20.160 200.815 21.070 201.035 ;
        RECT 22.605 200.815 23.955 201.045 ;
        RECT 16.645 200.135 23.955 200.815 ;
        RECT 24.015 200.220 24.445 201.005 ;
        RECT 24.560 200.815 25.480 201.045 ;
        RECT 32.580 200.815 33.490 201.035 ;
        RECT 35.025 200.815 36.795 201.045 ;
        RECT 39.150 200.845 40.095 201.045 ;
        RECT 24.560 200.135 28.025 200.815 ;
        RECT 29.065 200.135 36.795 200.815 ;
        RECT 37.345 200.165 40.095 200.845 ;
        RECT 11.265 199.925 11.435 200.135 ;
        RECT 12.645 199.925 12.815 200.135 ;
        RECT 16.320 199.975 16.440 200.085 ;
        RECT 16.785 199.945 16.955 200.135 ;
        RECT 18.165 199.925 18.335 200.115 ;
        RECT 21.845 199.925 22.015 200.115 ;
        RECT 23.225 199.925 23.395 200.115 ;
        RECT 25.070 199.925 25.240 200.115 ;
        RECT 27.825 199.945 27.995 200.135 ;
        RECT 28.295 199.980 28.455 200.090 ;
        RECT 28.745 199.925 28.915 200.115 ;
        RECT 29.205 199.925 29.375 200.135 ;
        RECT 37.490 200.115 37.660 200.165 ;
        RECT 39.150 200.135 40.095 200.165 ;
        RECT 40.105 200.815 41.035 201.045 ;
        RECT 40.105 200.135 42.855 200.815 ;
        RECT 42.880 200.135 44.695 201.045 ;
        RECT 44.705 200.135 48.375 200.945 ;
        RECT 48.385 200.135 49.755 200.945 ;
        RECT 49.775 200.220 50.205 201.005 ;
        RECT 50.235 200.135 52.965 201.045 ;
        RECT 52.985 200.135 58.495 200.945 ;
        RECT 58.505 200.135 61.255 200.945 ;
        RECT 63.085 200.815 64.015 201.045 ;
        RECT 61.265 200.135 64.015 200.815 ;
        RECT 64.035 200.135 66.765 201.045 ;
        RECT 66.785 200.845 67.730 201.045 ;
        RECT 66.785 200.165 69.535 200.845 ;
        RECT 66.785 200.135 67.730 200.165 ;
        RECT 32.885 199.925 33.055 200.115 ;
        RECT 33.345 199.925 33.515 200.115 ;
        RECT 37.020 199.975 37.140 200.085 ;
        RECT 37.485 199.945 37.660 200.115 ;
        RECT 42.545 199.945 42.715 200.135 ;
        RECT 37.485 199.925 37.655 199.945 ;
        RECT 43.005 199.925 43.175 200.135 ;
        RECT 44.845 199.945 45.015 200.135 ;
        RECT 46.695 199.970 46.855 200.080 ;
        RECT 47.610 199.925 47.780 200.115 ;
        RECT 48.525 199.945 48.695 200.135 ;
        RECT 48.980 199.925 49.150 200.115 ;
        RECT 50.365 199.945 50.535 200.135 ;
        RECT 51.285 199.925 51.455 200.115 ;
        RECT 53.125 199.945 53.295 200.135 ;
        RECT 54.505 199.925 54.675 200.115 ;
        RECT 58.645 199.945 58.815 200.135 ;
        RECT 60.025 199.925 60.195 200.115 ;
        RECT 61.405 199.945 61.575 200.135 ;
        RECT 63.245 199.925 63.415 200.115 ;
        RECT 64.165 199.945 64.335 200.135 ;
        RECT 68.775 199.970 68.935 200.080 ;
        RECT 69.220 199.945 69.390 200.165 ;
        RECT 69.545 200.135 70.915 200.945 ;
        RECT 71.235 200.815 72.165 201.045 ;
        RECT 71.235 200.135 73.070 200.815 ;
        RECT 73.245 200.135 74.595 201.045 ;
        RECT 75.535 200.220 75.965 201.005 ;
        RECT 75.985 200.135 81.495 200.945 ;
        RECT 81.505 200.135 82.875 200.945 ;
        RECT 82.885 200.845 83.815 201.045 ;
        RECT 85.145 200.845 86.095 201.045 ;
        RECT 82.885 200.365 86.095 200.845 ;
        RECT 83.030 200.165 86.095 200.365 ;
        RECT 69.685 199.945 69.855 200.135 ;
        RECT 72.905 200.115 73.070 200.135 ;
        RECT 11.125 199.115 12.495 199.925 ;
        RECT 12.505 199.115 18.015 199.925 ;
        RECT 18.025 199.115 21.695 199.925 ;
        RECT 21.705 199.115 23.075 199.925 ;
        RECT 23.100 199.015 24.915 199.925 ;
        RECT 24.925 199.015 26.755 199.925 ;
        RECT 26.765 199.245 29.055 199.925 ;
        RECT 26.765 199.015 27.685 199.245 ;
        RECT 29.065 199.115 31.815 199.925 ;
        RECT 31.825 199.145 33.195 199.925 ;
        RECT 33.205 199.115 36.875 199.925 ;
        RECT 36.895 199.055 37.325 199.840 ;
        RECT 37.345 199.115 42.855 199.925 ;
        RECT 42.865 199.115 46.535 199.925 ;
        RECT 47.465 199.015 48.815 199.925 ;
        RECT 48.865 199.015 50.215 199.925 ;
        RECT 51.245 199.015 54.355 199.925 ;
        RECT 54.365 199.115 59.875 199.925 ;
        RECT 59.885 199.115 62.635 199.925 ;
        RECT 62.655 199.055 63.085 199.840 ;
        RECT 63.105 199.115 68.615 199.925 ;
        RECT 69.545 199.895 70.490 199.925 ;
        RECT 71.980 199.895 72.150 200.115 ;
        RECT 72.445 199.925 72.615 200.115 ;
        RECT 72.905 199.945 73.075 200.115 ;
        RECT 73.360 199.945 73.530 200.135 ;
        RECT 74.755 199.980 74.915 200.090 ;
        RECT 76.125 200.085 76.295 200.135 ;
        RECT 76.120 199.975 76.295 200.085 ;
        RECT 76.125 199.945 76.295 199.975 ;
        RECT 76.585 199.925 76.755 200.115 ;
        RECT 78.880 199.975 79.000 200.085 ;
        RECT 79.345 199.925 79.515 200.115 ;
        RECT 81.645 199.925 81.815 200.135 ;
        RECT 83.030 200.115 83.200 200.165 ;
        RECT 85.160 200.135 86.095 200.165 ;
        RECT 86.105 200.135 88.855 200.945 ;
        RECT 88.865 200.135 90.235 200.915 ;
        RECT 90.245 200.135 95.755 200.945 ;
        RECT 95.765 200.135 99.435 200.945 ;
        RECT 99.905 200.135 101.275 200.915 ;
        RECT 101.295 200.220 101.725 201.005 ;
        RECT 101.785 200.815 103.135 201.045 ;
        RECT 104.670 200.815 105.580 201.035 ;
        RECT 112.220 200.815 113.140 201.045 ;
        RECT 101.785 200.135 109.095 200.815 ;
        RECT 109.675 200.135 113.140 200.815 ;
        RECT 113.245 200.135 114.615 200.945 ;
        RECT 118.140 200.815 119.050 201.035 ;
        RECT 120.585 200.815 122.355 201.045 ;
        RECT 114.625 200.135 122.355 200.815 ;
        RECT 122.445 200.135 126.115 200.945 ;
        RECT 127.055 200.220 127.485 201.005 ;
        RECT 127.505 200.135 133.015 200.945 ;
        RECT 133.025 200.135 138.535 200.945 ;
        RECT 138.545 200.135 144.055 200.945 ;
        RECT 144.065 200.135 147.735 200.945 ;
        RECT 147.745 200.135 149.115 200.945 ;
        RECT 149.125 200.135 150.495 200.945 ;
        RECT 83.025 199.945 83.200 200.115 ;
        RECT 83.030 199.925 83.195 199.945 ;
        RECT 85.325 199.925 85.495 200.115 ;
        RECT 86.245 199.945 86.415 200.135 ;
        RECT 88.080 199.975 88.200 200.085 ;
        RECT 89.005 199.925 89.175 200.135 ;
        RECT 90.385 199.945 90.555 200.135 ;
        RECT 90.840 199.975 90.960 200.085 ;
        RECT 91.305 199.925 91.475 200.115 ;
        RECT 94.525 199.925 94.695 200.115 ;
        RECT 95.905 199.945 96.075 200.135 ;
        RECT 98.200 199.975 98.320 200.085 ;
        RECT 98.665 199.925 98.835 200.115 ;
        RECT 99.580 199.975 99.700 200.085 ;
        RECT 100.045 199.945 100.215 200.135 ;
        RECT 104.185 199.925 104.355 200.115 ;
        RECT 104.640 199.975 104.760 200.085 ;
        RECT 105.105 199.925 105.275 200.115 ;
        RECT 108.785 199.945 108.955 200.135 ;
        RECT 109.240 199.975 109.360 200.085 ;
        RECT 109.705 199.945 109.875 200.135 ;
        RECT 112.925 199.925 113.095 200.115 ;
        RECT 113.385 199.945 113.555 200.135 ;
        RECT 114.765 199.945 114.935 200.135 ;
        RECT 114.785 199.925 114.935 199.945 ;
        RECT 117.985 199.925 118.155 200.115 ;
        RECT 118.445 199.925 118.615 200.115 ;
        RECT 122.135 199.970 122.295 200.080 ;
        RECT 122.585 199.945 122.755 200.135 ;
        RECT 126.275 199.980 126.435 200.090 ;
        RECT 127.645 199.945 127.815 200.135 ;
        RECT 129.945 199.925 130.115 200.115 ;
        RECT 130.405 199.925 130.575 200.115 ;
        RECT 133.165 199.945 133.335 200.135 ;
        RECT 135.925 199.925 136.095 200.115 ;
        RECT 138.685 199.945 138.855 200.135 ;
        RECT 139.600 199.975 139.720 200.085 ;
        RECT 140.525 199.925 140.695 200.115 ;
        RECT 144.205 199.945 144.375 200.135 ;
        RECT 146.045 199.925 146.215 200.115 ;
        RECT 147.885 199.945 148.055 200.135 ;
        RECT 148.800 199.975 148.920 200.085 ;
        RECT 150.185 199.925 150.355 200.135 ;
        RECT 69.545 199.215 72.295 199.895 ;
        RECT 69.545 199.015 70.490 199.215 ;
        RECT 72.305 199.115 75.975 199.925 ;
        RECT 76.445 199.245 78.735 199.925 ;
        RECT 79.205 199.245 81.495 199.925 ;
        RECT 77.815 199.015 78.735 199.245 ;
        RECT 80.575 199.015 81.495 199.245 ;
        RECT 81.505 199.115 82.875 199.925 ;
        RECT 83.030 199.245 84.865 199.925 ;
        RECT 83.935 199.015 84.865 199.245 ;
        RECT 85.185 199.115 87.935 199.925 ;
        RECT 88.415 199.055 88.845 199.840 ;
        RECT 88.865 199.115 90.695 199.925 ;
        RECT 91.205 199.015 94.375 199.925 ;
        RECT 94.385 199.115 98.055 199.925 ;
        RECT 98.525 199.245 100.815 199.925 ;
        RECT 99.895 199.015 100.815 199.245 ;
        RECT 100.920 199.245 104.385 199.925 ;
        RECT 104.965 199.245 112.695 199.925 ;
        RECT 100.920 199.015 101.840 199.245 ;
        RECT 108.480 199.025 109.390 199.245 ;
        RECT 110.925 199.015 112.695 199.245 ;
        RECT 112.785 199.115 114.155 199.925 ;
        RECT 114.175 199.055 114.605 199.840 ;
        RECT 114.785 199.105 116.715 199.925 ;
        RECT 116.925 199.145 118.295 199.925 ;
        RECT 118.305 199.115 121.975 199.925 ;
        RECT 122.945 199.245 130.255 199.925 ;
        RECT 115.765 199.015 116.715 199.105 ;
        RECT 122.945 199.015 124.295 199.245 ;
        RECT 125.830 199.025 126.740 199.245 ;
        RECT 130.265 199.115 135.775 199.925 ;
        RECT 135.785 199.115 139.455 199.925 ;
        RECT 139.935 199.055 140.365 199.840 ;
        RECT 140.385 199.115 145.895 199.925 ;
        RECT 145.905 199.115 148.655 199.925 ;
        RECT 149.125 199.115 150.495 199.925 ;
      LAYER nwell ;
        RECT 10.930 195.895 150.690 198.725 ;
      LAYER pwell ;
        RECT 11.125 194.695 12.495 195.505 ;
        RECT 12.505 194.695 18.015 195.505 ;
        RECT 18.025 194.695 23.535 195.505 ;
        RECT 24.015 194.780 24.445 195.565 ;
        RECT 24.465 194.695 29.975 195.505 ;
        RECT 29.985 194.695 35.495 195.505 ;
        RECT 35.505 194.695 38.255 195.505 ;
        RECT 40.085 195.375 41.015 195.605 ;
        RECT 42.830 195.405 43.775 195.605 ;
        RECT 38.265 194.695 41.015 195.375 ;
        RECT 41.025 194.725 43.775 195.405 ;
        RECT 11.265 194.485 11.435 194.695 ;
        RECT 12.645 194.485 12.815 194.695 ;
        RECT 14.945 194.485 15.115 194.675 ;
        RECT 15.400 194.535 15.520 194.645 ;
        RECT 15.865 194.485 16.035 194.675 ;
        RECT 18.165 194.505 18.335 194.695 ;
        RECT 23.225 194.485 23.395 194.675 ;
        RECT 23.680 194.535 23.800 194.645 ;
        RECT 24.605 194.505 24.775 194.695 ;
        RECT 30.125 194.505 30.295 194.695 ;
        RECT 30.590 194.485 30.760 194.675 ;
        RECT 34.265 194.485 34.435 194.675 ;
        RECT 35.645 194.505 35.815 194.695 ;
        RECT 36.115 194.530 36.275 194.640 ;
        RECT 37.490 194.485 37.660 194.675 ;
        RECT 38.405 194.505 38.575 194.695 ;
        RECT 41.170 194.505 41.340 194.725 ;
        RECT 42.830 194.695 43.775 194.725 ;
        RECT 43.785 194.695 45.615 195.605 ;
        RECT 45.625 194.695 49.295 195.505 ;
        RECT 49.775 194.780 50.205 195.565 ;
        RECT 50.225 194.695 55.735 195.505 ;
        RECT 55.745 194.695 57.575 195.505 ;
        RECT 57.585 195.405 58.515 195.605 ;
        RECT 59.845 195.405 60.795 195.605 ;
        RECT 57.585 194.925 60.795 195.405 ;
        RECT 64.320 195.375 65.230 195.595 ;
        RECT 66.765 195.375 68.115 195.605 ;
        RECT 57.730 194.725 60.795 194.925 ;
        RECT 43.005 194.485 43.175 194.675 ;
        RECT 43.460 194.535 43.580 194.645 ;
        RECT 43.925 194.485 44.095 194.675 ;
        RECT 45.300 194.505 45.470 194.695 ;
        RECT 45.765 194.505 45.935 194.695 ;
        RECT 47.145 194.485 47.315 194.675 ;
        RECT 49.440 194.535 49.560 194.645 ;
        RECT 50.365 194.485 50.535 194.695 ;
        RECT 55.885 194.675 56.055 194.695 ;
        RECT 53.120 194.535 53.240 194.645 ;
        RECT 55.880 194.505 56.055 194.675 ;
        RECT 57.730 194.505 57.900 194.725 ;
        RECT 59.860 194.695 60.795 194.725 ;
        RECT 60.805 194.695 68.115 195.375 ;
        RECT 68.165 194.695 69.995 195.505 ;
        RECT 70.005 195.405 70.950 195.605 ;
        RECT 70.005 194.725 72.755 195.405 ;
        RECT 70.005 194.695 70.950 194.725 ;
        RECT 11.125 193.675 12.495 194.485 ;
        RECT 12.505 193.675 13.875 194.485 ;
        RECT 13.885 193.705 15.255 194.485 ;
        RECT 15.725 193.805 23.035 194.485 ;
        RECT 23.085 193.805 30.395 194.485 ;
        RECT 30.445 193.805 34.115 194.485 ;
        RECT 34.125 193.805 35.955 194.485 ;
        RECT 19.240 193.585 20.150 193.805 ;
        RECT 21.685 193.575 23.035 193.805 ;
        RECT 26.600 193.585 27.510 193.805 ;
        RECT 29.045 193.575 30.395 193.805 ;
        RECT 32.525 193.575 34.115 193.805 ;
        RECT 34.610 193.575 35.955 193.805 ;
        RECT 36.895 193.615 37.325 194.400 ;
        RECT 37.345 193.575 40.265 194.485 ;
        RECT 40.565 193.805 43.315 194.485 ;
        RECT 40.565 193.575 41.495 193.805 ;
        RECT 43.825 193.575 46.995 194.485 ;
        RECT 47.105 193.575 50.215 194.485 ;
        RECT 50.225 193.675 52.975 194.485 ;
        RECT 53.445 194.455 54.390 194.485 ;
        RECT 55.880 194.455 56.050 194.505 ;
        RECT 58.185 194.485 58.355 194.675 ;
        RECT 58.645 194.485 58.815 194.675 ;
        RECT 60.480 194.535 60.600 194.645 ;
        RECT 60.945 194.485 61.115 194.695 ;
        RECT 62.320 194.535 62.440 194.645 ;
        RECT 63.250 194.485 63.420 194.675 ;
        RECT 67.380 194.485 67.550 194.675 ;
        RECT 67.845 194.485 68.015 194.675 ;
        RECT 68.305 194.505 68.475 194.695 ;
        RECT 69.680 194.535 69.800 194.645 ;
        RECT 71.065 194.485 71.235 194.675 ;
        RECT 71.525 194.485 71.695 194.675 ;
        RECT 72.440 194.505 72.610 194.725 ;
        RECT 72.765 194.695 75.515 195.505 ;
        RECT 75.535 194.780 75.965 195.565 ;
        RECT 75.985 194.695 77.815 195.505 ;
        RECT 78.875 195.375 79.805 195.605 ;
        RECT 81.175 195.375 82.105 195.605 ;
        RECT 77.970 194.695 79.805 195.375 ;
        RECT 80.270 194.695 82.105 195.375 ;
        RECT 82.425 195.405 83.355 195.605 ;
        RECT 84.685 195.405 85.635 195.605 ;
        RECT 82.425 194.925 85.635 195.405 ;
        RECT 82.570 194.725 85.635 194.925 ;
        RECT 72.905 194.505 73.075 194.695 ;
        RECT 76.125 194.505 76.295 194.695 ;
        RECT 77.970 194.675 78.135 194.695 ;
        RECT 80.270 194.675 80.435 194.695 ;
        RECT 77.045 194.505 77.215 194.675 ;
        RECT 77.965 194.505 78.135 194.675 ;
        RECT 79.340 194.535 79.460 194.645 ;
        RECT 77.065 194.485 77.215 194.505 ;
        RECT 53.445 193.775 56.195 194.455 ;
        RECT 56.205 193.805 58.495 194.485 ;
        RECT 53.445 193.575 54.390 193.775 ;
        RECT 56.205 193.575 57.125 193.805 ;
        RECT 58.505 193.675 60.335 194.485 ;
        RECT 60.805 193.705 62.175 194.485 ;
        RECT 62.655 193.615 63.085 194.400 ;
        RECT 63.105 193.575 66.025 194.485 ;
        RECT 66.345 193.575 67.695 194.485 ;
        RECT 67.705 193.675 69.535 194.485 ;
        RECT 70.015 193.575 71.365 194.485 ;
        RECT 71.385 193.675 76.895 194.485 ;
        RECT 77.065 193.665 78.995 194.485 ;
        RECT 79.810 194.455 79.980 194.675 ;
        RECT 80.265 194.505 80.435 194.675 ;
        RECT 82.570 194.505 82.740 194.725 ;
        RECT 84.700 194.695 85.635 194.725 ;
        RECT 85.645 194.695 87.475 195.505 ;
        RECT 87.945 194.695 89.315 195.475 ;
        RECT 92.840 195.375 93.750 195.595 ;
        RECT 95.285 195.375 97.055 195.605 ;
        RECT 89.325 194.695 97.055 195.375 ;
        RECT 97.145 194.695 100.815 195.505 ;
        RECT 101.295 194.780 101.725 195.565 ;
        RECT 103.115 195.375 104.035 195.605 ;
        RECT 101.745 194.695 104.035 195.375 ;
        RECT 104.355 195.375 105.285 195.605 ;
        RECT 104.355 194.695 106.190 195.375 ;
        RECT 106.345 194.695 107.715 195.475 ;
        RECT 107.725 194.695 111.395 195.505 ;
        RECT 115.525 195.375 116.455 195.605 ;
        RECT 112.555 194.695 116.455 195.375 ;
        RECT 116.465 194.695 120.135 195.505 ;
        RECT 120.145 194.695 121.975 195.605 ;
        RECT 121.985 194.695 125.655 195.505 ;
        RECT 125.665 194.695 127.035 195.505 ;
        RECT 127.055 194.780 127.485 195.565 ;
        RECT 127.505 194.695 133.015 195.505 ;
        RECT 133.025 194.695 138.535 195.505 ;
        RECT 138.545 194.695 144.055 195.505 ;
        RECT 144.065 194.695 147.735 195.505 ;
        RECT 147.745 194.695 149.115 195.505 ;
        RECT 149.125 194.695 150.495 195.505 ;
        RECT 83.025 194.485 83.195 194.675 ;
        RECT 84.405 194.485 84.575 194.675 ;
        RECT 85.785 194.485 85.955 194.695 ;
        RECT 87.620 194.535 87.740 194.645 ;
        RECT 88.085 194.505 88.255 194.695 ;
        RECT 89.005 194.485 89.175 194.675 ;
        RECT 89.465 194.505 89.635 194.695 ;
        RECT 96.825 194.485 96.995 194.675 ;
        RECT 97.285 194.505 97.455 194.695 ;
        RECT 98.205 194.485 98.375 194.675 ;
        RECT 100.960 194.535 101.080 194.645 ;
        RECT 101.435 194.530 101.595 194.640 ;
        RECT 101.885 194.505 102.055 194.695 ;
        RECT 106.025 194.675 106.190 194.695 ;
        RECT 102.350 194.485 102.520 194.675 ;
        RECT 106.025 194.485 106.195 194.675 ;
        RECT 107.405 194.505 107.575 194.695 ;
        RECT 107.865 194.645 108.035 194.695 ;
        RECT 107.860 194.535 108.035 194.645 ;
        RECT 107.865 194.505 108.035 194.535 ;
        RECT 108.600 194.485 108.770 194.675 ;
        RECT 111.555 194.540 111.715 194.650 ;
        RECT 112.465 194.485 112.635 194.675 ;
        RECT 114.765 194.485 114.935 194.675 ;
        RECT 115.870 194.505 116.040 194.695 ;
        RECT 116.605 194.505 116.775 194.695 ;
        RECT 120.290 194.505 120.460 194.695 ;
        RECT 120.745 194.485 120.915 194.675 ;
        RECT 81.940 194.455 82.875 194.485 ;
        RECT 79.810 194.255 82.875 194.455 ;
        RECT 78.045 193.575 78.995 193.665 ;
        RECT 79.665 193.775 82.875 194.255 ;
        RECT 79.665 193.575 80.595 193.775 ;
        RECT 81.925 193.575 82.875 193.775 ;
        RECT 82.885 193.675 84.255 194.485 ;
        RECT 84.265 193.705 85.635 194.485 ;
        RECT 85.645 193.675 88.395 194.485 ;
        RECT 88.415 193.615 88.845 194.400 ;
        RECT 88.865 193.805 96.595 194.485 ;
        RECT 92.380 193.585 93.290 193.805 ;
        RECT 94.825 193.575 96.595 193.805 ;
        RECT 96.685 193.675 98.055 194.485 ;
        RECT 98.065 193.575 101.275 194.485 ;
        RECT 102.205 193.805 105.875 194.485 ;
        RECT 102.205 193.575 103.130 193.805 ;
        RECT 105.885 193.675 107.715 194.485 ;
        RECT 108.185 193.805 112.085 194.485 ;
        RECT 108.185 193.575 109.115 193.805 ;
        RECT 112.325 193.675 114.155 194.485 ;
        RECT 114.175 193.615 114.605 194.400 ;
        RECT 114.625 193.675 118.295 194.485 ;
        RECT 118.315 193.575 121.045 194.485 ;
        RECT 121.205 194.455 121.375 194.675 ;
        RECT 122.125 194.505 122.295 194.695 ;
        RECT 124.890 194.485 125.060 194.675 ;
        RECT 125.345 194.505 125.515 194.675 ;
        RECT 125.805 194.505 125.975 194.695 ;
        RECT 125.365 194.485 125.515 194.505 ;
        RECT 127.645 194.485 127.815 194.695 ;
        RECT 133.165 194.505 133.335 194.695 ;
        RECT 135.465 194.485 135.635 194.675 ;
        RECT 138.685 194.505 138.855 194.695 ;
        RECT 139.155 194.530 139.315 194.640 ;
        RECT 140.525 194.485 140.695 194.675 ;
        RECT 144.205 194.505 144.375 194.695 ;
        RECT 146.045 194.485 146.215 194.675 ;
        RECT 147.885 194.505 148.055 194.695 ;
        RECT 148.800 194.535 148.920 194.645 ;
        RECT 150.185 194.485 150.355 194.695 ;
        RECT 122.405 194.455 123.785 194.485 ;
        RECT 121.080 193.775 123.785 194.455 ;
        RECT 122.405 193.575 123.785 193.775 ;
        RECT 123.825 193.575 125.175 194.485 ;
        RECT 125.365 193.665 127.295 194.485 ;
        RECT 127.505 193.805 135.235 194.485 ;
        RECT 126.345 193.575 127.295 193.665 ;
        RECT 131.020 193.585 131.930 193.805 ;
        RECT 133.465 193.575 135.235 193.805 ;
        RECT 135.325 193.675 138.995 194.485 ;
        RECT 139.935 193.615 140.365 194.400 ;
        RECT 140.385 193.675 145.895 194.485 ;
        RECT 145.905 193.675 148.655 194.485 ;
        RECT 149.125 193.675 150.495 194.485 ;
      LAYER nwell ;
        RECT 10.930 190.455 150.690 193.285 ;
      LAYER pwell ;
        RECT 11.125 189.255 12.495 190.065 ;
        RECT 16.020 189.935 16.930 190.155 ;
        RECT 18.465 189.935 19.815 190.165 ;
        RECT 12.505 189.255 19.815 189.935 ;
        RECT 19.865 189.935 21.210 190.165 ;
        RECT 19.865 189.255 21.695 189.935 ;
        RECT 21.705 189.255 23.075 190.035 ;
        RECT 24.015 189.340 24.445 190.125 ;
        RECT 24.465 189.255 27.215 190.065 ;
        RECT 27.225 189.935 28.570 190.165 ;
        RECT 30.870 189.965 31.815 190.165 ;
        RECT 27.225 189.255 29.055 189.935 ;
        RECT 29.065 189.285 31.815 189.965 ;
        RECT 11.265 189.045 11.435 189.255 ;
        RECT 12.645 189.045 12.815 189.255 ;
        RECT 16.325 189.045 16.495 189.235 ;
        RECT 16.780 189.095 16.900 189.205 ;
        RECT 17.245 189.045 17.415 189.235 ;
        RECT 19.545 189.045 19.715 189.235 ;
        RECT 21.385 189.065 21.555 189.255 ;
        RECT 22.765 189.065 22.935 189.255 ;
        RECT 23.235 189.205 23.395 189.210 ;
        RECT 23.220 189.100 23.395 189.205 ;
        RECT 23.220 189.095 23.340 189.100 ;
        RECT 23.685 189.045 23.855 189.235 ;
        RECT 24.605 189.065 24.775 189.255 ;
        RECT 26.905 189.045 27.075 189.235 ;
        RECT 27.365 189.045 27.535 189.235 ;
        RECT 28.745 189.065 28.915 189.255 ;
        RECT 29.210 189.065 29.380 189.285 ;
        RECT 30.870 189.255 31.815 189.285 ;
        RECT 32.285 189.965 33.235 190.165 ;
        RECT 34.565 189.965 35.495 190.165 ;
        RECT 32.285 189.485 35.495 189.965 ;
        RECT 32.285 189.285 35.350 189.485 ;
        RECT 32.285 189.255 33.220 189.285 ;
        RECT 30.120 189.095 30.240 189.205 ;
        RECT 30.580 189.045 30.750 189.235 ;
        RECT 31.965 189.205 32.135 189.235 ;
        RECT 31.960 189.095 32.135 189.205 ;
        RECT 31.965 189.045 32.135 189.095 ;
        RECT 35.180 189.065 35.350 189.285 ;
        RECT 35.505 189.255 39.175 190.065 ;
        RECT 39.185 189.255 41.000 190.165 ;
        RECT 41.025 189.255 46.535 190.065 ;
        RECT 46.545 189.255 49.295 190.065 ;
        RECT 49.775 189.340 50.205 190.125 ;
        RECT 50.225 189.255 52.975 190.065 ;
        RECT 53.295 189.935 54.225 190.165 ;
        RECT 53.295 189.255 55.130 189.935 ;
        RECT 55.285 189.255 56.655 190.035 ;
        RECT 56.665 189.255 62.175 190.065 ;
        RECT 62.185 189.255 67.695 190.065 ;
        RECT 67.705 189.255 69.535 190.065 ;
        RECT 70.025 189.255 71.375 190.165 ;
        RECT 71.385 189.255 75.055 190.065 ;
        RECT 75.535 189.340 75.965 190.125 ;
        RECT 75.985 189.255 77.815 190.065 ;
        RECT 78.285 189.255 79.655 190.035 ;
        RECT 79.665 189.255 85.175 190.065 ;
        RECT 85.185 189.255 86.555 190.065 ;
        RECT 86.650 189.255 95.755 189.935 ;
        RECT 95.765 189.255 99.420 190.165 ;
        RECT 99.445 189.255 101.275 190.065 ;
        RECT 101.295 189.340 101.725 190.125 ;
        RECT 101.745 189.255 110.850 189.935 ;
        RECT 110.945 189.255 114.115 190.165 ;
        RECT 114.165 189.255 115.995 190.065 ;
        RECT 116.465 189.255 121.055 190.165 ;
        RECT 121.065 189.255 124.275 190.165 ;
        RECT 124.285 189.255 127.035 190.065 ;
        RECT 127.055 189.340 127.485 190.125 ;
        RECT 127.505 189.255 130.715 190.165 ;
        RECT 130.725 189.255 132.095 190.035 ;
        RECT 132.105 189.255 137.615 190.065 ;
        RECT 137.625 189.255 143.135 190.065 ;
        RECT 143.145 189.255 148.655 190.065 ;
        RECT 149.125 189.255 150.495 190.065 ;
        RECT 35.645 189.045 35.815 189.255 ;
        RECT 37.485 189.045 37.655 189.235 ;
        RECT 40.240 189.095 40.360 189.205 ;
        RECT 40.705 189.045 40.875 189.255 ;
        RECT 41.165 189.065 41.335 189.255 ;
        RECT 43.925 189.045 44.095 189.235 ;
        RECT 46.685 189.065 46.855 189.255 ;
        RECT 49.440 189.095 49.560 189.205 ;
        RECT 50.365 189.045 50.535 189.255 ;
        RECT 54.965 189.235 55.130 189.255 ;
        RECT 50.835 189.090 50.995 189.200 ;
        RECT 51.740 189.045 51.910 189.235 ;
        RECT 53.125 189.045 53.295 189.235 ;
        RECT 54.965 189.065 55.135 189.235 ;
        RECT 55.425 189.045 55.595 189.255 ;
        RECT 56.805 189.065 56.975 189.255 ;
        RECT 62.325 189.065 62.495 189.255 ;
        RECT 67.845 189.235 68.015 189.255 ;
        RECT 66.465 189.045 66.635 189.235 ;
        RECT 66.935 189.090 67.095 189.200 ;
        RECT 67.845 189.065 68.020 189.235 ;
        RECT 69.680 189.095 69.800 189.205 ;
        RECT 70.140 189.065 70.310 189.255 ;
        RECT 71.525 189.235 71.695 189.255 ;
        RECT 71.525 189.065 71.700 189.235 ;
        RECT 67.850 189.045 68.020 189.065 ;
        RECT 11.125 188.235 12.495 189.045 ;
        RECT 12.505 188.235 13.875 189.045 ;
        RECT 13.885 188.365 16.635 189.045 ;
        RECT 17.105 188.365 19.395 189.045 ;
        RECT 13.885 188.135 14.815 188.365 ;
        RECT 18.475 188.135 19.395 188.365 ;
        RECT 19.405 188.235 23.075 189.045 ;
        RECT 23.545 188.365 25.835 189.045 ;
        RECT 24.915 188.135 25.835 188.365 ;
        RECT 25.845 188.265 27.215 189.045 ;
        RECT 27.225 188.235 29.975 189.045 ;
        RECT 30.465 188.135 31.815 189.045 ;
        RECT 31.825 188.235 35.495 189.045 ;
        RECT 35.505 188.235 36.875 189.045 ;
        RECT 36.895 188.175 37.325 188.960 ;
        RECT 37.345 188.235 40.095 189.045 ;
        RECT 40.665 188.135 43.775 189.045 ;
        RECT 43.785 188.235 49.295 189.045 ;
        RECT 49.315 188.135 50.665 189.045 ;
        RECT 51.625 188.135 52.975 189.045 ;
        RECT 52.985 188.365 55.275 189.045 ;
        RECT 55.285 188.365 62.595 189.045 ;
        RECT 54.355 188.135 55.275 188.365 ;
        RECT 58.800 188.145 59.710 188.365 ;
        RECT 61.245 188.135 62.595 188.365 ;
        RECT 62.655 188.175 63.085 188.960 ;
        RECT 63.105 188.365 66.775 189.045 ;
        RECT 63.105 188.135 64.035 188.365 ;
        RECT 67.705 188.135 71.360 189.045 ;
        RECT 71.530 189.015 71.700 189.065 ;
        RECT 74.290 189.045 74.460 189.235 ;
        RECT 75.200 189.095 75.320 189.205 ;
        RECT 75.660 189.095 75.780 189.205 ;
        RECT 76.125 189.065 76.295 189.255 ;
        RECT 77.965 189.205 78.135 189.235 ;
        RECT 77.960 189.095 78.135 189.205 ;
        RECT 77.965 189.045 78.135 189.095 ;
        RECT 78.435 189.065 78.605 189.255 ;
        RECT 79.805 189.065 79.975 189.255 ;
        RECT 73.190 189.015 74.135 189.045 ;
        RECT 71.385 188.335 74.135 189.015 ;
        RECT 73.190 188.135 74.135 188.335 ;
        RECT 74.145 188.135 75.495 189.045 ;
        RECT 75.985 188.135 78.275 189.045 ;
        RECT 79.205 189.015 80.155 189.045 ;
        RECT 82.560 189.015 82.730 189.235 ;
        RECT 83.025 189.015 83.195 189.235 ;
        RECT 85.325 189.065 85.495 189.255 ;
        RECT 85.785 189.045 85.955 189.235 ;
        RECT 88.085 189.045 88.255 189.235 ;
        RECT 89.005 189.045 89.175 189.235 ;
        RECT 90.840 189.095 90.960 189.205 ;
        RECT 91.305 189.045 91.475 189.235 ;
        RECT 94.525 189.045 94.695 189.235 ;
        RECT 95.445 189.065 95.615 189.255 ;
        RECT 95.910 189.205 96.080 189.255 ;
        RECT 95.900 189.095 96.080 189.205 ;
        RECT 95.910 189.065 96.080 189.095 ;
        RECT 84.240 189.015 85.635 189.045 ;
        RECT 79.205 188.335 82.875 189.015 ;
        RECT 82.900 188.335 85.635 189.015 ;
        RECT 79.205 188.135 80.155 188.335 ;
        RECT 84.225 188.135 85.635 188.335 ;
        RECT 85.645 188.235 87.015 189.045 ;
        RECT 87.035 188.135 88.385 189.045 ;
        RECT 88.415 188.175 88.845 188.960 ;
        RECT 88.865 188.235 90.695 189.045 ;
        RECT 91.165 188.135 94.375 189.045 ;
        RECT 94.395 188.135 95.745 189.045 ;
        RECT 96.225 189.015 97.170 189.045 ;
        RECT 98.660 189.015 98.830 189.235 ;
        RECT 99.125 189.045 99.295 189.235 ;
        RECT 99.585 189.065 99.755 189.255 ;
        RECT 101.885 189.065 102.055 189.255 ;
        RECT 103.720 189.045 103.890 189.235 ;
        RECT 104.185 189.045 104.355 189.235 ;
        RECT 106.485 189.045 106.655 189.235 ;
        RECT 106.945 189.045 107.115 189.235 ;
        RECT 112.465 189.045 112.635 189.235 ;
        RECT 113.845 189.065 114.015 189.255 ;
        RECT 114.305 189.065 114.475 189.255 ;
        RECT 114.765 189.045 114.935 189.235 ;
        RECT 116.140 189.095 116.260 189.205 ;
        RECT 116.610 189.065 116.780 189.255 ;
        RECT 117.985 189.045 118.155 189.235 ;
        RECT 121.205 189.065 121.375 189.255 ;
        RECT 123.505 189.045 123.675 189.235 ;
        RECT 124.425 189.065 124.595 189.255 ;
        RECT 129.025 189.045 129.195 189.235 ;
        RECT 130.405 189.065 130.575 189.255 ;
        RECT 131.785 189.065 131.955 189.255 ;
        RECT 132.245 189.065 132.415 189.255 ;
        RECT 134.545 189.045 134.715 189.235 ;
        RECT 137.765 189.065 137.935 189.255 ;
        RECT 140.525 189.045 140.695 189.235 ;
        RECT 143.285 189.065 143.455 189.255 ;
        RECT 146.045 189.045 146.215 189.235 ;
        RECT 148.800 189.095 148.920 189.205 ;
        RECT 150.185 189.045 150.355 189.255 ;
        RECT 96.225 188.335 98.975 189.015 ;
        RECT 96.225 188.135 97.170 188.335 ;
        RECT 98.985 188.235 100.355 189.045 ;
        RECT 100.380 188.135 104.035 189.045 ;
        RECT 104.045 188.235 105.415 189.045 ;
        RECT 105.435 188.135 106.785 189.045 ;
        RECT 106.805 188.235 112.315 189.045 ;
        RECT 112.325 188.235 114.155 189.045 ;
        RECT 114.175 188.175 114.605 188.960 ;
        RECT 114.625 188.365 117.835 189.045 ;
        RECT 116.700 188.135 117.835 188.365 ;
        RECT 117.845 188.235 123.355 189.045 ;
        RECT 123.365 188.235 128.875 189.045 ;
        RECT 128.885 188.235 134.395 189.045 ;
        RECT 134.405 188.235 139.915 189.045 ;
        RECT 139.935 188.175 140.365 188.960 ;
        RECT 140.385 188.235 145.895 189.045 ;
        RECT 145.905 188.235 148.655 189.045 ;
        RECT 149.125 188.235 150.495 189.045 ;
      LAYER nwell ;
        RECT 10.930 185.015 150.690 187.845 ;
      LAYER pwell ;
        RECT 11.125 183.815 12.495 184.625 ;
        RECT 12.505 183.815 16.175 184.625 ;
        RECT 18.155 184.495 19.085 184.725 ;
        RECT 17.250 183.815 19.085 184.495 ;
        RECT 19.405 183.815 20.755 184.725 ;
        RECT 20.785 183.815 23.535 184.625 ;
        RECT 24.015 183.900 24.445 184.685 ;
        RECT 24.475 183.815 27.205 184.725 ;
        RECT 27.225 183.815 29.055 184.725 ;
        RECT 31.035 184.495 31.965 184.725 ;
        RECT 30.130 183.815 31.965 184.495 ;
        RECT 32.285 183.815 35.495 184.725 ;
        RECT 35.525 183.815 36.875 184.725 ;
        RECT 37.345 183.815 39.635 184.725 ;
        RECT 41.910 184.525 42.855 184.725 ;
        RECT 40.105 183.845 42.855 184.525 ;
        RECT 11.265 183.605 11.435 183.815 ;
        RECT 12.645 183.605 12.815 183.815 ;
        RECT 17.250 183.795 17.415 183.815 ;
        RECT 15.400 183.655 15.520 183.765 ;
        RECT 16.335 183.660 16.495 183.770 ;
        RECT 17.245 183.605 17.415 183.795 ;
        RECT 17.715 183.650 17.875 183.760 ;
        RECT 20.470 183.625 20.640 183.815 ;
        RECT 20.925 183.625 21.095 183.815 ;
        RECT 21.845 183.605 22.015 183.795 ;
        RECT 22.305 183.605 22.475 183.795 ;
        RECT 23.680 183.655 23.800 183.765 ;
        RECT 24.605 183.625 24.775 183.815 ;
        RECT 27.825 183.605 27.995 183.795 ;
        RECT 28.740 183.625 28.910 183.815 ;
        RECT 30.130 183.795 30.295 183.815 ;
        RECT 29.215 183.660 29.375 183.770 ;
        RECT 30.125 183.625 30.295 183.795 ;
        RECT 30.585 183.625 30.755 183.795 ;
        RECT 32.425 183.625 32.595 183.815 ;
        RECT 30.590 183.605 30.755 183.625 ;
        RECT 32.885 183.605 33.055 183.795 ;
        RECT 35.640 183.625 35.810 183.815 ;
        RECT 37.490 183.795 37.660 183.815 ;
        RECT 36.560 183.655 36.680 183.765 ;
        RECT 37.020 183.655 37.140 183.765 ;
        RECT 37.485 183.625 37.660 183.795 ;
        RECT 39.780 183.655 39.900 183.765 ;
        RECT 40.250 183.625 40.420 183.845 ;
        RECT 41.910 183.815 42.855 183.845 ;
        RECT 42.865 183.815 45.615 184.625 ;
        RECT 46.085 183.815 48.375 184.725 ;
        RECT 48.385 183.815 49.755 184.625 ;
        RECT 49.775 183.900 50.205 184.685 ;
        RECT 50.515 183.815 53.435 184.725 ;
        RECT 53.445 183.815 58.955 184.625 ;
        RECT 58.965 183.815 62.635 184.625 ;
        RECT 63.105 183.815 64.935 184.725 ;
        RECT 64.945 183.815 66.775 184.625 ;
        RECT 68.295 184.495 69.225 184.725 ;
        RECT 67.390 183.815 69.225 184.495 ;
        RECT 69.545 183.815 70.915 184.625 ;
        RECT 70.925 184.525 71.880 184.725 ;
        RECT 70.925 183.845 73.205 184.525 ;
        RECT 70.925 183.815 71.880 183.845 ;
        RECT 37.485 183.605 37.655 183.625 ;
        RECT 41.165 183.605 41.335 183.795 ;
        RECT 43.005 183.625 43.175 183.815 ;
        RECT 43.925 183.605 44.095 183.795 ;
        RECT 44.385 183.605 44.555 183.795 ;
        RECT 45.760 183.655 45.880 183.765 ;
        RECT 48.065 183.625 48.235 183.815 ;
        RECT 48.525 183.625 48.695 183.815 ;
        RECT 11.125 182.795 12.495 183.605 ;
        RECT 12.505 182.795 15.255 183.605 ;
        RECT 15.725 182.695 17.540 183.605 ;
        RECT 18.580 182.925 22.045 183.605 ;
        RECT 18.580 182.695 19.500 182.925 ;
        RECT 22.165 182.795 27.675 183.605 ;
        RECT 27.685 182.795 30.435 183.605 ;
        RECT 30.590 182.925 32.425 183.605 ;
        RECT 31.495 182.695 32.425 182.925 ;
        RECT 32.745 182.795 36.415 183.605 ;
        RECT 36.895 182.735 37.325 183.520 ;
        RECT 37.345 182.795 41.015 183.605 ;
        RECT 41.025 182.795 42.395 183.605 ;
        RECT 42.405 182.925 44.235 183.605 ;
        RECT 42.405 182.695 43.750 182.925 ;
        RECT 44.245 182.795 49.755 183.605 ;
        RECT 49.765 183.575 50.720 183.605 ;
        RECT 51.750 183.575 51.920 183.795 ;
        RECT 52.205 183.605 52.375 183.795 ;
        RECT 53.120 183.625 53.290 183.815 ;
        RECT 53.585 183.625 53.755 183.815 ;
        RECT 56.345 183.605 56.515 183.795 ;
        RECT 56.805 183.605 56.975 183.795 ;
        RECT 59.105 183.625 59.275 183.815 ;
        RECT 60.480 183.655 60.600 183.765 ;
        RECT 62.325 183.605 62.495 183.795 ;
        RECT 62.780 183.655 62.900 183.765 ;
        RECT 63.250 183.625 63.420 183.815 ;
        RECT 65.085 183.625 65.255 183.815 ;
        RECT 67.390 183.795 67.555 183.815 ;
        RECT 66.460 183.605 66.630 183.795 ;
        RECT 66.925 183.765 67.095 183.795 ;
        RECT 66.920 183.655 67.095 183.765 ;
        RECT 66.925 183.605 67.095 183.655 ;
        RECT 67.385 183.625 67.555 183.795 ;
        RECT 69.685 183.625 69.855 183.815 ;
        RECT 72.445 183.605 72.615 183.795 ;
        RECT 72.910 183.625 73.080 183.845 ;
        RECT 73.225 183.815 75.055 184.625 ;
        RECT 75.535 183.900 75.965 184.685 ;
        RECT 76.965 183.815 78.735 184.725 ;
        RECT 79.230 184.495 80.575 184.725 ;
        RECT 78.745 183.815 80.575 184.495 ;
        RECT 80.585 183.815 84.255 184.625 ;
        RECT 84.765 183.815 87.935 184.725 ;
        RECT 87.945 183.815 89.315 184.625 ;
        RECT 89.325 184.495 90.245 184.725 ;
        RECT 89.325 183.815 91.615 184.495 ;
        RECT 91.625 183.815 97.135 184.625 ;
        RECT 97.145 183.815 100.815 184.625 ;
        RECT 101.295 183.900 101.725 184.685 ;
        RECT 101.745 183.815 104.915 184.725 ;
        RECT 104.965 183.815 107.715 184.625 ;
        RECT 107.795 183.815 111.855 184.725 ;
        RECT 111.865 183.815 114.905 184.725 ;
        RECT 115.105 183.815 116.455 184.725 ;
        RECT 116.465 183.815 118.295 184.625 ;
        RECT 118.765 183.815 121.685 184.725 ;
        RECT 125.885 184.635 126.835 184.725 ;
        RECT 121.985 183.815 124.735 184.625 ;
        RECT 124.905 183.815 126.835 184.635 ;
        RECT 127.055 183.900 127.485 184.685 ;
        RECT 131.020 184.495 131.930 184.715 ;
        RECT 133.465 184.495 135.235 184.725 ;
        RECT 127.505 183.815 135.235 184.495 ;
        RECT 135.325 183.815 140.835 184.625 ;
        RECT 140.845 183.815 146.355 184.625 ;
        RECT 146.365 183.815 149.115 184.625 ;
        RECT 149.125 183.815 150.495 184.625 ;
        RECT 73.365 183.625 73.535 183.815 ;
        RECT 75.200 183.655 75.320 183.765 ;
        RECT 76.135 183.660 76.295 183.770 ;
        RECT 77.045 183.625 77.215 183.795 ;
        RECT 77.045 183.605 77.210 183.625 ;
        RECT 77.505 183.605 77.675 183.795 ;
        RECT 78.420 183.625 78.590 183.815 ;
        RECT 78.885 183.625 79.055 183.815 ;
        RECT 80.725 183.625 80.895 183.815 ;
        RECT 83.025 183.605 83.195 183.795 ;
        RECT 84.400 183.655 84.520 183.765 ;
        RECT 84.865 183.625 85.035 183.815 ;
        RECT 88.085 183.625 88.255 183.815 ;
        RECT 89.000 183.655 89.120 183.765 ;
        RECT 89.465 183.605 89.635 183.795 ;
        RECT 91.305 183.625 91.475 183.815 ;
        RECT 91.765 183.625 91.935 183.815 ;
        RECT 92.685 183.605 92.855 183.795 ;
        RECT 97.285 183.625 97.455 183.815 ;
        RECT 98.205 183.605 98.375 183.795 ;
        RECT 100.960 183.655 101.080 183.765 ;
        RECT 101.880 183.655 102.000 183.765 ;
        RECT 102.345 183.605 102.515 183.795 ;
        RECT 104.645 183.625 104.815 183.815 ;
        RECT 105.105 183.625 105.275 183.815 ;
        RECT 111.545 183.605 111.715 183.815 ;
        RECT 114.760 183.795 114.905 183.815 ;
        RECT 112.005 183.605 112.175 183.795 ;
        RECT 113.840 183.655 113.960 183.765 ;
        RECT 114.760 183.625 114.935 183.795 ;
        RECT 116.140 183.625 116.310 183.815 ;
        RECT 116.605 183.625 116.775 183.815 ;
        RECT 118.440 183.655 118.560 183.765 ;
        RECT 118.910 183.625 119.080 183.815 ;
        RECT 114.765 183.605 114.935 183.625 ;
        RECT 119.820 183.605 119.990 183.795 ;
        RECT 120.275 183.605 120.445 183.795 ;
        RECT 122.125 183.625 122.295 183.815 ;
        RECT 124.905 183.795 125.055 183.815 ;
        RECT 123.500 183.655 123.620 183.765 ;
        RECT 123.965 183.605 124.135 183.795 ;
        RECT 124.885 183.625 125.055 183.795 ;
        RECT 127.185 183.605 127.355 183.795 ;
        RECT 127.645 183.625 127.815 183.815 ;
        RECT 130.865 183.605 131.035 183.795 ;
        RECT 131.325 183.605 131.495 183.795 ;
        RECT 135.465 183.625 135.635 183.815 ;
        RECT 136.845 183.605 137.015 183.795 ;
        RECT 139.600 183.655 139.720 183.765 ;
        RECT 140.525 183.605 140.695 183.795 ;
        RECT 140.985 183.625 141.155 183.815 ;
        RECT 146.045 183.605 146.215 183.795 ;
        RECT 146.505 183.625 146.675 183.815 ;
        RECT 148.800 183.655 148.920 183.765 ;
        RECT 150.185 183.605 150.355 183.815 ;
        RECT 49.765 182.895 52.045 183.575 ;
        RECT 49.765 182.695 50.720 182.895 ;
        RECT 52.065 182.795 54.815 183.605 ;
        RECT 54.825 182.695 56.640 183.605 ;
        RECT 56.665 182.795 60.335 183.605 ;
        RECT 60.805 182.695 62.620 183.605 ;
        RECT 62.655 182.735 63.085 183.520 ;
        RECT 63.300 182.695 66.775 183.605 ;
        RECT 66.785 182.795 72.295 183.605 ;
        RECT 72.305 182.795 75.055 183.605 ;
        RECT 75.375 182.925 77.210 183.605 ;
        RECT 75.375 182.695 76.305 182.925 ;
        RECT 77.365 182.795 82.875 183.605 ;
        RECT 82.885 182.795 88.395 183.605 ;
        RECT 88.415 182.735 88.845 183.520 ;
        RECT 89.365 182.695 92.535 183.605 ;
        RECT 92.545 182.795 98.055 183.605 ;
        RECT 98.065 182.795 101.735 183.605 ;
        RECT 102.205 182.925 109.935 183.605 ;
        RECT 105.720 182.705 106.630 182.925 ;
        RECT 108.165 182.695 109.935 182.925 ;
        RECT 110.025 182.695 111.840 183.605 ;
        RECT 111.865 182.795 113.695 183.605 ;
        RECT 114.175 182.735 114.605 183.520 ;
        RECT 114.625 182.795 116.455 183.605 ;
        RECT 116.550 182.925 120.135 183.605 ;
        RECT 119.215 182.695 120.135 182.925 ;
        RECT 120.145 182.695 123.355 183.605 ;
        RECT 123.825 182.695 127.035 183.605 ;
        RECT 127.045 182.795 129.795 183.605 ;
        RECT 129.805 182.825 131.175 183.605 ;
        RECT 131.185 182.795 136.695 183.605 ;
        RECT 136.705 182.795 139.455 183.605 ;
        RECT 139.935 182.735 140.365 183.520 ;
        RECT 140.385 182.795 145.895 183.605 ;
        RECT 145.905 182.795 148.655 183.605 ;
        RECT 149.125 182.795 150.495 183.605 ;
      LAYER nwell ;
        RECT 10.930 179.575 150.690 182.405 ;
      LAYER pwell ;
        RECT 11.125 178.375 12.495 179.185 ;
        RECT 16.940 179.055 17.850 179.275 ;
        RECT 19.385 179.055 21.155 179.285 ;
        RECT 13.425 178.375 21.155 179.055 ;
        RECT 22.165 178.375 23.980 179.285 ;
        RECT 24.015 178.460 24.445 179.245 ;
        RECT 27.980 179.055 28.890 179.275 ;
        RECT 30.425 179.055 31.775 179.285 ;
        RECT 24.465 178.375 31.775 179.055 ;
        RECT 31.825 179.055 33.170 179.285 ;
        RECT 31.825 178.375 33.655 179.055 ;
        RECT 34.605 178.375 35.955 179.285 ;
        RECT 39.480 179.055 40.390 179.275 ;
        RECT 41.925 179.055 43.275 179.285 ;
        RECT 35.965 178.375 43.275 179.055 ;
        RECT 43.325 178.375 47.855 179.285 ;
        RECT 47.925 178.375 49.755 179.185 ;
        RECT 49.775 178.460 50.205 179.245 ;
        RECT 50.225 179.085 51.170 179.285 ;
        RECT 52.505 179.085 53.435 179.285 ;
        RECT 50.225 178.605 53.435 179.085 ;
        RECT 50.225 178.405 53.295 178.605 ;
        RECT 50.225 178.375 51.170 178.405 ;
        RECT 11.265 178.165 11.435 178.375 ;
        RECT 12.645 178.165 12.815 178.355 ;
        RECT 13.565 178.185 13.735 178.375 ;
        RECT 16.335 178.210 16.495 178.320 ;
        RECT 18.620 178.165 18.790 178.355 ;
        RECT 19.085 178.165 19.255 178.355 ;
        RECT 21.395 178.220 21.555 178.330 ;
        RECT 23.685 178.185 23.855 178.375 ;
        RECT 24.605 178.185 24.775 178.375 ;
        RECT 25.980 178.165 26.150 178.355 ;
        RECT 26.445 178.165 26.615 178.355 ;
        RECT 31.960 178.215 32.080 178.325 ;
        RECT 33.345 178.185 33.515 178.375 ;
        RECT 33.815 178.220 33.975 178.330 ;
        RECT 34.265 178.185 34.435 178.355 ;
        RECT 34.265 178.165 34.415 178.185 ;
        RECT 34.730 178.165 34.900 178.355 ;
        RECT 35.640 178.185 35.810 178.375 ;
        RECT 36.105 178.185 36.275 178.375 ;
        RECT 36.560 178.215 36.680 178.325 ;
        RECT 43.470 178.185 43.640 178.375 ;
        RECT 46.225 178.165 46.395 178.355 ;
        RECT 46.695 178.210 46.855 178.320 ;
        RECT 47.605 178.165 47.775 178.355 ;
        RECT 48.065 178.185 48.235 178.375 ;
        RECT 53.125 178.185 53.295 178.405 ;
        RECT 53.445 178.375 55.275 179.185 ;
        RECT 55.300 178.375 58.955 179.285 ;
        RECT 59.905 178.375 61.255 179.285 ;
        RECT 61.265 178.375 64.935 179.185 ;
        RECT 64.945 178.375 66.315 179.185 ;
        RECT 66.425 178.375 68.615 179.285 ;
        RECT 68.625 178.375 74.135 179.185 ;
        RECT 74.145 178.375 75.515 179.185 ;
        RECT 75.535 178.460 75.965 179.245 ;
        RECT 75.985 178.375 77.815 179.185 ;
        RECT 78.305 178.375 79.655 179.285 ;
        RECT 83.640 179.055 84.550 179.275 ;
        RECT 86.085 179.055 87.435 179.285 ;
        RECT 80.125 178.375 87.435 179.055 ;
        RECT 87.485 178.375 91.545 179.285 ;
        RECT 91.720 179.055 92.640 179.285 ;
        RECT 91.720 178.375 95.185 179.055 ;
        RECT 95.305 178.375 98.415 179.285 ;
        RECT 98.525 178.375 99.875 179.285 ;
        RECT 99.905 178.375 101.275 179.185 ;
        RECT 101.295 178.460 101.725 179.245 ;
        RECT 101.745 178.375 103.115 179.185 ;
        RECT 103.125 178.375 104.495 179.155 ;
        RECT 104.505 178.375 110.015 179.185 ;
        RECT 110.025 178.375 111.855 179.185 ;
        RECT 112.325 178.375 115.075 179.285 ;
        RECT 115.085 178.375 117.295 179.285 ;
        RECT 118.505 179.195 119.455 179.285 ;
        RECT 118.505 178.375 120.435 179.195 ;
        RECT 120.605 178.375 123.355 179.185 ;
        RECT 123.365 179.085 124.320 179.285 ;
        RECT 123.365 178.405 125.645 179.085 ;
        RECT 123.365 178.375 124.320 178.405 ;
        RECT 53.585 178.185 53.755 178.375 ;
        RECT 58.640 178.185 58.810 178.375 ;
        RECT 60.940 178.355 61.110 178.375 ;
        RECT 59.115 178.220 59.275 178.330 ;
        RECT 60.940 178.185 61.115 178.355 ;
        RECT 60.945 178.165 61.115 178.185 ;
        RECT 61.405 178.165 61.575 178.375 ;
        RECT 65.085 178.185 65.255 178.375 ;
        RECT 11.125 177.355 12.495 178.165 ;
        RECT 12.505 177.355 16.175 178.165 ;
        RECT 17.105 177.255 18.935 178.165 ;
        RECT 18.945 177.355 24.455 178.165 ;
        RECT 24.465 177.255 26.295 178.165 ;
        RECT 26.305 177.355 31.815 178.165 ;
        RECT 32.485 177.345 34.415 178.165 ;
        RECT 32.485 177.255 33.435 177.345 ;
        RECT 34.585 177.255 36.415 178.165 ;
        RECT 36.895 177.295 37.325 178.080 ;
        RECT 37.430 177.485 46.535 178.165 ;
        RECT 47.465 177.485 56.570 178.165 ;
        RECT 56.675 178.125 57.595 178.165 ;
        RECT 56.665 177.935 57.595 178.125 ;
        RECT 59.685 177.935 61.255 178.165 ;
        RECT 56.665 177.575 61.255 177.935 ;
        RECT 56.675 177.485 61.255 177.575 ;
        RECT 56.675 177.255 59.675 177.485 ;
        RECT 61.265 177.355 62.635 178.165 ;
        RECT 63.105 178.135 64.040 178.165 ;
        RECT 66.000 178.135 66.170 178.355 ;
        RECT 66.465 178.165 66.635 178.355 ;
        RECT 68.300 178.185 68.470 178.375 ;
        RECT 68.765 178.185 68.935 178.375 ;
        RECT 69.225 178.165 69.395 178.355 ;
        RECT 71.065 178.165 71.235 178.355 ;
        RECT 74.285 178.185 74.455 178.375 ;
        RECT 76.125 178.185 76.295 178.375 ;
        RECT 77.960 178.215 78.080 178.325 ;
        RECT 79.340 178.185 79.510 178.375 ;
        RECT 80.265 178.355 80.435 178.375 ;
        RECT 79.800 178.215 79.920 178.325 ;
        RECT 80.265 178.185 80.440 178.355 ;
        RECT 62.655 177.295 63.085 178.080 ;
        RECT 63.105 177.935 66.170 178.135 ;
        RECT 63.105 177.455 66.315 177.935 ;
        RECT 63.105 177.255 64.055 177.455 ;
        RECT 65.385 177.255 66.315 177.455 ;
        RECT 66.335 177.255 69.065 178.165 ;
        RECT 69.085 177.355 70.915 178.165 ;
        RECT 70.925 177.485 78.235 178.165 ;
        RECT 74.440 177.265 75.350 177.485 ;
        RECT 76.885 177.255 78.235 177.485 ;
        RECT 78.285 178.135 79.240 178.165 ;
        RECT 80.270 178.135 80.440 178.185 ;
        RECT 80.725 178.165 80.895 178.355 ;
        RECT 82.565 178.165 82.735 178.355 ;
        RECT 85.325 178.165 85.495 178.355 ;
        RECT 87.625 178.185 87.795 178.375 ;
        RECT 88.080 178.215 88.200 178.325 ;
        RECT 89.005 178.165 89.175 178.355 ;
        RECT 90.840 178.215 90.960 178.325 ;
        RECT 94.525 178.165 94.695 178.355 ;
        RECT 94.985 178.185 95.155 178.375 ;
        RECT 95.900 178.165 96.070 178.355 ;
        RECT 96.365 178.165 96.535 178.355 ;
        RECT 98.205 178.185 98.375 178.375 ;
        RECT 99.590 178.185 99.760 178.375 ;
        RECT 100.045 178.165 100.215 178.375 ;
        RECT 101.885 178.185 102.055 178.375 ;
        RECT 102.810 178.165 102.980 178.355 ;
        RECT 103.265 178.185 103.435 178.375 ;
        RECT 104.645 178.185 104.815 178.375 ;
        RECT 106.490 178.165 106.660 178.355 ;
        RECT 110.165 178.165 110.335 178.375 ;
        RECT 112.000 178.215 112.120 178.325 ;
        RECT 113.840 178.215 113.960 178.325 ;
        RECT 114.765 178.165 114.935 178.375 ;
        RECT 115.230 178.185 115.400 178.375 ;
        RECT 120.285 178.355 120.435 178.375 ;
        RECT 117.530 178.165 117.700 178.355 ;
        RECT 118.905 178.165 119.075 178.355 ;
        RECT 120.285 178.185 120.455 178.355 ;
        RECT 120.745 178.185 120.915 178.375 ;
        RECT 121.660 178.215 121.780 178.325 ;
        RECT 122.125 178.185 122.295 178.355 ;
        RECT 125.350 178.185 125.520 178.405 ;
        RECT 125.665 178.375 127.035 179.185 ;
        RECT 127.055 178.460 127.485 179.245 ;
        RECT 127.505 178.375 129.335 179.285 ;
        RECT 129.345 178.375 134.855 179.185 ;
        RECT 134.865 178.375 140.375 179.185 ;
        RECT 140.385 178.375 145.895 179.185 ;
        RECT 145.905 178.375 148.655 179.185 ;
        RECT 149.125 178.375 150.495 179.185 ;
        RECT 122.125 178.165 122.325 178.185 ;
        RECT 125.805 178.165 125.975 178.375 ;
        RECT 129.020 178.185 129.190 178.375 ;
        RECT 129.485 178.185 129.655 178.375 ;
        RECT 131.325 178.165 131.495 178.355 ;
        RECT 135.005 178.185 135.175 178.375 ;
        RECT 136.845 178.165 137.015 178.355 ;
        RECT 139.600 178.215 139.720 178.325 ;
        RECT 140.525 178.165 140.695 178.375 ;
        RECT 146.045 178.165 146.215 178.375 ;
        RECT 148.800 178.215 148.920 178.325 ;
        RECT 150.185 178.165 150.355 178.375 ;
        RECT 78.285 177.455 80.565 178.135 ;
        RECT 78.285 177.255 79.240 177.455 ;
        RECT 80.585 177.355 82.415 178.165 ;
        RECT 82.425 177.255 85.175 178.165 ;
        RECT 85.185 177.355 87.935 178.165 ;
        RECT 88.415 177.295 88.845 178.080 ;
        RECT 88.865 177.355 90.695 178.165 ;
        RECT 91.165 177.485 94.835 178.165 ;
        RECT 91.165 177.255 92.095 177.485 ;
        RECT 94.865 177.255 96.215 178.165 ;
        RECT 96.225 177.355 99.895 178.165 ;
        RECT 99.905 177.485 102.655 178.165 ;
        RECT 101.725 177.255 102.655 177.485 ;
        RECT 102.665 177.255 106.335 178.165 ;
        RECT 106.345 177.255 110.015 178.165 ;
        RECT 110.025 177.355 113.695 178.165 ;
        RECT 114.175 177.295 114.605 178.080 ;
        RECT 114.625 177.355 117.375 178.165 ;
        RECT 117.385 177.255 118.735 178.165 ;
        RECT 118.765 177.355 121.515 178.165 ;
        RECT 122.125 177.485 125.655 178.165 ;
        RECT 122.830 177.255 125.655 177.485 ;
        RECT 125.665 177.355 131.175 178.165 ;
        RECT 131.185 177.355 136.695 178.165 ;
        RECT 136.705 177.355 139.455 178.165 ;
        RECT 139.935 177.295 140.365 178.080 ;
        RECT 140.385 177.355 145.895 178.165 ;
        RECT 145.905 177.355 148.655 178.165 ;
        RECT 149.125 177.355 150.495 178.165 ;
      LAYER nwell ;
        RECT 10.930 174.135 150.690 176.965 ;
      LAYER pwell ;
        RECT 11.125 172.935 12.495 173.745 ;
        RECT 12.505 172.935 16.175 173.745 ;
        RECT 16.185 172.935 17.555 173.715 ;
        RECT 17.565 172.935 23.075 173.745 ;
        RECT 24.015 173.020 24.445 173.805 ;
        RECT 24.465 172.935 29.975 173.745 ;
        RECT 29.985 172.935 35.495 173.745 ;
        RECT 35.505 172.935 37.335 173.745 ;
        RECT 37.345 172.935 38.695 173.845 ;
        RECT 38.725 172.935 41.475 173.745 ;
        RECT 44.025 173.615 45.615 173.845 ;
        RECT 41.945 172.935 45.615 173.615 ;
        RECT 45.625 172.935 49.295 173.745 ;
        RECT 49.775 173.020 50.205 173.805 ;
        RECT 51.365 173.755 52.315 173.845 ;
        RECT 50.385 172.935 52.315 173.755 ;
        RECT 52.605 172.935 54.815 173.845 ;
        RECT 54.825 172.935 56.655 173.845 ;
        RECT 56.665 172.935 62.175 173.745 ;
        RECT 62.185 172.935 64.015 173.745 ;
        RECT 64.025 172.935 65.395 173.715 ;
        RECT 65.405 172.935 67.235 173.745 ;
        RECT 67.245 172.935 70.455 173.845 ;
        RECT 70.465 172.935 72.295 173.745 ;
        RECT 72.320 172.935 74.135 173.845 ;
        RECT 74.145 172.935 75.515 173.745 ;
        RECT 75.535 173.020 75.965 173.805 ;
        RECT 75.985 172.935 77.815 173.845 ;
        RECT 77.825 172.935 81.495 173.745 ;
        RECT 82.520 173.615 83.440 173.845 ;
        RECT 82.520 172.935 85.985 173.615 ;
        RECT 86.105 172.935 89.775 173.745 ;
        RECT 89.785 173.615 90.715 173.845 ;
        RECT 89.785 172.935 93.685 173.615 ;
        RECT 93.925 172.935 97.595 173.745 ;
        RECT 98.075 172.935 100.815 173.615 ;
        RECT 101.295 173.020 101.725 173.805 ;
        RECT 101.755 172.935 103.105 173.845 ;
        RECT 103.125 172.935 108.635 173.745 ;
        RECT 109.105 172.935 112.025 173.845 ;
        RECT 112.325 172.935 114.155 173.845 ;
        RECT 115.745 173.755 116.695 173.845 ;
        RECT 114.165 172.935 115.535 173.745 ;
        RECT 115.745 172.935 117.675 173.755 ;
        RECT 118.765 172.935 120.595 173.845 ;
        RECT 120.605 172.935 123.815 173.845 ;
        RECT 123.825 172.935 126.575 173.745 ;
        RECT 127.055 173.020 127.485 173.805 ;
        RECT 127.505 172.935 133.015 173.745 ;
        RECT 133.025 172.935 138.535 173.745 ;
        RECT 138.545 172.935 144.055 173.745 ;
        RECT 144.065 172.935 147.735 173.745 ;
        RECT 147.745 172.935 149.115 173.745 ;
        RECT 149.125 172.935 150.495 173.745 ;
        RECT 11.265 172.725 11.435 172.935 ;
        RECT 12.645 172.725 12.815 172.935 ;
        RECT 14.480 172.775 14.600 172.885 ;
        RECT 14.945 172.725 15.115 172.915 ;
        RECT 17.245 172.745 17.415 172.935 ;
        RECT 17.705 172.745 17.875 172.935 ;
        RECT 22.315 172.770 22.475 172.880 ;
        RECT 23.235 172.780 23.395 172.890 ;
        RECT 24.605 172.745 24.775 172.935 ;
        RECT 25.065 172.725 25.235 172.915 ;
        RECT 25.525 172.725 25.695 172.915 ;
        RECT 11.125 171.915 12.495 172.725 ;
        RECT 12.505 171.915 14.335 172.725 ;
        RECT 14.805 172.045 22.115 172.725 ;
        RECT 18.320 171.825 19.230 172.045 ;
        RECT 20.765 171.815 22.115 172.045 ;
        RECT 23.085 172.045 25.375 172.725 ;
        RECT 23.085 171.815 24.005 172.045 ;
        RECT 25.385 171.915 28.135 172.725 ;
        RECT 28.290 172.695 28.460 172.915 ;
        RECT 30.125 172.745 30.295 172.935 ;
        RECT 31.515 172.770 31.675 172.880 ;
        RECT 32.430 172.725 32.600 172.915 ;
        RECT 35.645 172.725 35.815 172.935 ;
        RECT 37.490 172.915 37.660 172.935 ;
        RECT 37.485 172.745 37.660 172.915 ;
        RECT 38.865 172.915 39.035 172.935 ;
        RECT 42.090 172.915 42.260 172.935 ;
        RECT 38.865 172.745 39.040 172.915 ;
        RECT 41.620 172.775 41.740 172.885 ;
        RECT 37.485 172.725 37.655 172.745 ;
        RECT 30.420 172.695 31.355 172.725 ;
        RECT 28.290 172.495 31.355 172.695 ;
        RECT 28.145 172.015 31.355 172.495 ;
        RECT 28.145 171.815 29.075 172.015 ;
        RECT 30.405 171.815 31.355 172.015 ;
        RECT 32.285 171.815 35.205 172.725 ;
        RECT 35.505 171.915 36.875 172.725 ;
        RECT 36.895 171.855 37.325 172.640 ;
        RECT 37.345 171.915 38.715 172.725 ;
        RECT 38.870 172.695 39.040 172.745 ;
        RECT 42.080 172.745 42.260 172.915 ;
        RECT 41.000 172.695 41.935 172.725 ;
        RECT 42.080 172.695 42.250 172.745 ;
        RECT 44.390 172.725 44.560 172.915 ;
        RECT 45.765 172.745 45.935 172.935 ;
        RECT 50.385 172.915 50.535 172.935 ;
        RECT 46.685 172.725 46.855 172.915 ;
        RECT 48.525 172.745 48.695 172.915 ;
        RECT 49.440 172.775 49.560 172.885 ;
        RECT 50.365 172.745 50.535 172.915 ;
        RECT 48.530 172.725 48.695 172.745 ;
        RECT 50.825 172.725 50.995 172.915 ;
        RECT 54.500 172.745 54.670 172.935 ;
        RECT 54.970 172.745 55.140 172.935 ;
        RECT 56.345 172.725 56.515 172.915 ;
        RECT 56.805 172.745 56.975 172.935 ;
        RECT 43.280 172.695 44.235 172.725 ;
        RECT 38.870 172.495 41.935 172.695 ;
        RECT 38.725 172.015 41.935 172.495 ;
        RECT 41.955 172.015 44.235 172.695 ;
        RECT 38.725 171.815 39.655 172.015 ;
        RECT 40.985 171.815 41.935 172.015 ;
        RECT 43.280 171.815 44.235 172.015 ;
        RECT 44.245 171.815 46.535 172.725 ;
        RECT 46.545 171.915 48.375 172.725 ;
        RECT 48.530 172.045 50.365 172.725 ;
        RECT 49.435 171.815 50.365 172.045 ;
        RECT 50.685 171.915 56.195 172.725 ;
        RECT 56.205 171.915 58.035 172.725 ;
        RECT 58.180 172.695 58.350 172.915 ;
        RECT 60.485 172.725 60.655 172.915 ;
        RECT 62.325 172.885 62.495 172.935 ;
        RECT 62.320 172.775 62.495 172.885 ;
        RECT 62.325 172.745 62.495 172.775 ;
        RECT 63.245 172.725 63.415 172.915 ;
        RECT 64.165 172.745 64.335 172.935 ;
        RECT 65.545 172.745 65.715 172.935 ;
        RECT 70.145 172.745 70.315 172.935 ;
        RECT 70.605 172.725 70.775 172.935 ;
        RECT 72.445 172.885 72.615 172.935 ;
        RECT 74.285 172.915 74.455 172.935 ;
        RECT 72.440 172.775 72.615 172.885 ;
        RECT 72.445 172.745 72.615 172.775 ;
        RECT 73.825 172.725 73.995 172.915 ;
        RECT 74.280 172.745 74.455 172.915 ;
        RECT 76.130 172.745 76.300 172.935 ;
        RECT 77.965 172.745 78.135 172.935 ;
        RECT 59.380 172.695 60.335 172.725 ;
        RECT 58.055 172.015 60.335 172.695 ;
        RECT 59.380 171.815 60.335 172.015 ;
        RECT 60.345 171.915 62.175 172.725 ;
        RECT 62.655 171.855 63.085 172.640 ;
        RECT 63.105 172.045 70.415 172.725 ;
        RECT 66.620 171.825 67.530 172.045 ;
        RECT 69.065 171.815 70.415 172.045 ;
        RECT 70.465 171.915 72.295 172.725 ;
        RECT 72.775 171.815 74.125 172.725 ;
        RECT 74.280 172.695 74.450 172.745 ;
        RECT 78.425 172.725 78.595 172.915 ;
        RECT 78.885 172.725 79.055 172.915 ;
        RECT 81.655 172.780 81.815 172.890 ;
        RECT 85.785 172.745 85.955 172.935 ;
        RECT 86.245 172.745 86.415 172.935 ;
        RECT 86.705 172.725 86.875 172.915 ;
        RECT 89.000 172.775 89.120 172.885 ;
        RECT 75.480 172.695 76.435 172.725 ;
        RECT 74.155 172.015 76.435 172.695 ;
        RECT 75.480 171.815 76.435 172.015 ;
        RECT 76.445 172.045 78.735 172.725 ;
        RECT 78.745 172.045 86.475 172.725 ;
        RECT 76.445 171.815 77.365 172.045 ;
        RECT 82.260 171.825 83.170 172.045 ;
        RECT 84.705 171.815 86.475 172.045 ;
        RECT 86.565 171.915 88.395 172.725 ;
        RECT 89.470 172.695 89.640 172.915 ;
        RECT 90.200 172.745 90.370 172.935 ;
        RECT 91.130 172.695 92.075 172.725 ;
        RECT 92.230 172.695 92.400 172.915 ;
        RECT 94.065 172.745 94.235 172.935 ;
        RECT 94.985 172.725 95.155 172.915 ;
        RECT 97.740 172.775 97.860 172.885 ;
        RECT 100.505 172.725 100.675 172.935 ;
        RECT 100.960 172.775 101.080 172.885 ;
        RECT 101.885 172.745 102.055 172.935 ;
        RECT 102.805 172.725 102.975 172.915 ;
        RECT 103.265 172.725 103.435 172.935 ;
        RECT 109.250 172.915 109.420 172.935 ;
        RECT 113.840 172.915 114.010 172.935 ;
        RECT 108.780 172.775 108.900 172.885 ;
        RECT 109.245 172.745 109.420 172.915 ;
        RECT 109.245 172.725 109.415 172.745 ;
        RECT 109.705 172.725 109.875 172.915 ;
        RECT 111.540 172.775 111.660 172.885 ;
        RECT 113.840 172.745 114.015 172.915 ;
        RECT 114.305 172.745 114.475 172.935 ;
        RECT 117.525 172.915 117.675 172.935 ;
        RECT 113.845 172.725 114.010 172.745 ;
        RECT 114.765 172.725 114.935 172.915 ;
        RECT 116.600 172.775 116.720 172.885 ;
        RECT 117.065 172.745 117.235 172.915 ;
        RECT 117.525 172.745 117.695 172.915 ;
        RECT 117.995 172.780 118.155 172.890 ;
        RECT 118.910 172.745 119.080 172.935 ;
        RECT 117.070 172.725 117.235 172.745 ;
        RECT 119.365 172.725 119.535 172.915 ;
        RECT 120.745 172.745 120.915 172.935 ;
        RECT 123.045 172.725 123.215 172.915 ;
        RECT 123.965 172.745 124.135 172.935 ;
        RECT 126.720 172.775 126.840 172.885 ;
        RECT 127.645 172.745 127.815 172.935 ;
        RECT 130.865 172.725 131.035 172.915 ;
        RECT 133.165 172.745 133.335 172.935 ;
        RECT 136.385 172.725 136.555 172.915 ;
        RECT 138.685 172.745 138.855 172.935 ;
        RECT 140.525 172.725 140.695 172.915 ;
        RECT 144.205 172.745 144.375 172.935 ;
        RECT 146.045 172.725 146.215 172.915 ;
        RECT 147.885 172.745 148.055 172.935 ;
        RECT 148.800 172.775 148.920 172.885 ;
        RECT 150.185 172.725 150.355 172.935 ;
        RECT 93.890 172.695 94.835 172.725 ;
        RECT 88.415 171.855 88.845 172.640 ;
        RECT 89.325 172.015 92.075 172.695 ;
        RECT 92.085 172.015 94.835 172.695 ;
        RECT 91.130 171.815 92.075 172.015 ;
        RECT 93.890 171.815 94.835 172.015 ;
        RECT 94.845 171.915 100.355 172.725 ;
        RECT 100.365 171.915 101.735 172.725 ;
        RECT 101.755 171.815 103.105 172.725 ;
        RECT 103.125 171.915 105.875 172.725 ;
        RECT 105.980 172.045 109.445 172.725 ;
        RECT 105.980 171.815 106.900 172.045 ;
        RECT 109.565 171.915 111.395 172.725 ;
        RECT 112.175 172.045 114.010 172.725 ;
        RECT 112.175 171.815 113.105 172.045 ;
        RECT 114.175 171.855 114.605 172.640 ;
        RECT 114.640 171.815 116.455 172.725 ;
        RECT 117.070 172.045 118.905 172.725 ;
        RECT 117.975 171.815 118.905 172.045 ;
        RECT 119.225 171.915 122.895 172.725 ;
        RECT 122.905 172.045 130.635 172.725 ;
        RECT 126.420 171.825 127.330 172.045 ;
        RECT 128.865 171.815 130.635 172.045 ;
        RECT 130.725 171.915 136.235 172.725 ;
        RECT 136.245 171.915 139.915 172.725 ;
        RECT 139.935 171.855 140.365 172.640 ;
        RECT 140.385 171.915 145.895 172.725 ;
        RECT 145.905 171.915 148.655 172.725 ;
        RECT 149.125 171.915 150.495 172.725 ;
      LAYER nwell ;
        RECT 10.930 168.695 150.690 171.525 ;
      LAYER pwell ;
        RECT 11.125 167.495 12.495 168.305 ;
        RECT 12.505 167.495 15.255 168.305 ;
        RECT 15.265 168.205 16.195 168.405 ;
        RECT 17.525 168.205 18.475 168.405 ;
        RECT 15.265 167.725 18.475 168.205 ;
        RECT 15.410 167.525 18.475 167.725 ;
        RECT 11.265 167.285 11.435 167.495 ;
        RECT 12.645 167.285 12.815 167.495 ;
        RECT 15.410 167.305 15.580 167.525 ;
        RECT 17.540 167.495 18.475 167.525 ;
        RECT 18.485 167.495 20.315 168.305 ;
        RECT 20.325 167.495 21.675 168.405 ;
        RECT 22.015 168.175 22.945 168.405 ;
        RECT 22.015 167.495 23.850 168.175 ;
        RECT 24.015 167.580 24.445 168.365 ;
        RECT 24.665 168.315 25.615 168.405 ;
        RECT 24.665 167.495 26.595 168.315 ;
        RECT 26.765 167.495 28.595 168.405 ;
        RECT 32.580 168.175 33.490 168.395 ;
        RECT 35.025 168.175 36.375 168.405 ;
        RECT 29.065 167.495 36.375 168.175 ;
        RECT 36.425 167.495 37.795 168.305 ;
        RECT 37.805 168.175 38.725 168.405 ;
        RECT 37.805 167.495 40.095 168.175 ;
        RECT 40.105 167.495 41.475 168.305 ;
        RECT 41.485 167.495 43.300 168.405 ;
        RECT 43.325 167.495 48.835 168.305 ;
        RECT 49.775 167.580 50.205 168.365 ;
        RECT 50.225 167.495 53.335 168.405 ;
        RECT 53.445 167.495 56.555 168.405 ;
        RECT 56.665 167.495 59.415 168.405 ;
        RECT 59.435 167.495 60.785 168.405 ;
        RECT 60.805 167.495 66.315 168.305 ;
        RECT 70.300 168.175 71.210 168.395 ;
        RECT 72.745 168.175 74.095 168.405 ;
        RECT 66.785 167.495 74.095 168.175 ;
        RECT 74.145 167.495 75.515 168.305 ;
        RECT 75.535 167.580 75.965 168.365 ;
        RECT 76.070 167.495 85.175 168.175 ;
        RECT 85.685 167.495 88.855 168.405 ;
        RECT 88.865 167.495 94.375 168.305 ;
        RECT 94.385 167.495 98.055 168.305 ;
        RECT 98.065 167.495 101.275 168.405 ;
        RECT 101.295 167.580 101.725 168.365 ;
        RECT 105.260 168.175 106.170 168.395 ;
        RECT 107.705 168.175 109.475 168.405 ;
        RECT 101.745 167.495 109.475 168.175 ;
        RECT 109.565 167.495 113.685 168.405 ;
        RECT 113.705 167.495 116.455 168.305 ;
        RECT 116.465 168.175 117.385 168.405 ;
        RECT 116.465 167.495 118.755 168.175 ;
        RECT 118.765 167.495 120.115 168.405 ;
        RECT 122.205 168.315 123.155 168.405 ;
        RECT 121.225 167.495 123.155 168.315 ;
        RECT 124.285 167.495 125.655 168.275 ;
        RECT 125.665 167.495 127.035 168.305 ;
        RECT 127.055 167.580 127.485 168.365 ;
        RECT 127.505 167.495 133.015 168.305 ;
        RECT 133.025 167.495 138.535 168.305 ;
        RECT 138.545 167.495 144.055 168.305 ;
        RECT 144.065 167.495 147.735 168.305 ;
        RECT 147.745 167.495 149.115 168.305 ;
        RECT 149.125 167.495 150.495 168.305 ;
        RECT 18.165 167.285 18.335 167.475 ;
        RECT 18.625 167.305 18.795 167.495 ;
        RECT 20.470 167.305 20.640 167.495 ;
        RECT 23.685 167.475 23.850 167.495 ;
        RECT 26.445 167.475 26.595 167.495 ;
        RECT 23.685 167.285 23.855 167.475 ;
        RECT 25.520 167.335 25.640 167.445 ;
        RECT 25.985 167.285 26.155 167.475 ;
        RECT 26.445 167.305 26.615 167.475 ;
        RECT 28.280 167.305 28.450 167.495 ;
        RECT 28.740 167.335 28.860 167.445 ;
        RECT 29.205 167.305 29.375 167.495 ;
        RECT 29.660 167.335 29.780 167.445 ;
        RECT 30.125 167.285 30.295 167.475 ;
        RECT 33.805 167.285 33.975 167.475 ;
        RECT 34.265 167.285 34.435 167.475 ;
        RECT 36.565 167.305 36.735 167.495 ;
        RECT 37.485 167.285 37.655 167.475 ;
        RECT 39.785 167.305 39.955 167.495 ;
        RECT 40.245 167.305 40.415 167.495 ;
        RECT 41.165 167.285 41.335 167.475 ;
        RECT 43.005 167.305 43.175 167.495 ;
        RECT 43.465 167.305 43.635 167.495 ;
        RECT 44.385 167.285 44.555 167.475 ;
        RECT 48.995 167.340 49.155 167.450 ;
        RECT 49.905 167.285 50.075 167.475 ;
        RECT 51.740 167.335 51.860 167.445 ;
        RECT 53.125 167.305 53.295 167.495 ;
        RECT 53.585 167.285 53.755 167.475 ;
        RECT 54.045 167.285 54.215 167.475 ;
        RECT 56.345 167.305 56.515 167.495 ;
        RECT 56.805 167.305 56.975 167.495 ;
        RECT 59.565 167.285 59.735 167.475 ;
        RECT 60.485 167.305 60.655 167.495 ;
        RECT 60.945 167.305 61.115 167.495 ;
        RECT 66.925 167.475 67.095 167.495 ;
        RECT 62.320 167.335 62.440 167.445 ;
        RECT 63.245 167.285 63.415 167.475 ;
        RECT 66.460 167.335 66.580 167.445 ;
        RECT 66.920 167.305 67.095 167.475 ;
        RECT 66.920 167.285 67.090 167.305 ;
        RECT 69.225 167.285 69.395 167.475 ;
        RECT 69.685 167.285 69.855 167.475 ;
        RECT 73.360 167.335 73.480 167.445 ;
        RECT 73.825 167.285 73.995 167.475 ;
        RECT 74.285 167.305 74.455 167.495 ;
        RECT 79.800 167.285 79.970 167.475 ;
        RECT 80.265 167.285 80.435 167.475 ;
        RECT 84.865 167.305 85.035 167.495 ;
        RECT 85.320 167.335 85.440 167.445 ;
        RECT 85.785 167.285 85.955 167.495 ;
        RECT 89.005 167.285 89.175 167.495 ;
        RECT 91.765 167.285 91.935 167.475 ;
        RECT 94.525 167.305 94.695 167.495 ;
        RECT 94.985 167.285 95.155 167.475 ;
        RECT 96.825 167.285 96.995 167.475 ;
        RECT 100.515 167.330 100.675 167.440 ;
        RECT 100.975 167.305 101.145 167.495 ;
        RECT 101.425 167.285 101.595 167.475 ;
        RECT 101.885 167.305 102.055 167.495 ;
        RECT 103.265 167.285 103.435 167.475 ;
        RECT 106.955 167.330 107.115 167.440 ;
        RECT 108.140 167.285 108.310 167.475 ;
        RECT 109.705 167.305 109.875 167.495 ;
        RECT 111.545 167.305 111.715 167.495 ;
        RECT 113.380 167.285 113.550 167.475 ;
        RECT 113.845 167.445 114.015 167.495 ;
        RECT 113.840 167.335 114.015 167.445 ;
        RECT 113.845 167.305 114.015 167.335 ;
        RECT 114.765 167.285 114.935 167.475 ;
        RECT 118.445 167.285 118.615 167.495 ;
        RECT 119.830 167.305 120.000 167.495 ;
        RECT 121.225 167.475 121.375 167.495 ;
        RECT 120.285 167.285 120.455 167.475 ;
        RECT 121.205 167.305 121.375 167.475 ;
        RECT 123.515 167.340 123.675 167.450 ;
        RECT 123.965 167.285 124.135 167.475 ;
        RECT 125.345 167.305 125.515 167.495 ;
        RECT 125.805 167.305 125.975 167.495 ;
        RECT 127.645 167.475 127.815 167.495 ;
        RECT 127.640 167.305 127.815 167.475 ;
        RECT 127.640 167.285 127.810 167.305 ;
        RECT 128.105 167.285 128.275 167.475 ;
        RECT 133.165 167.305 133.335 167.495 ;
        RECT 133.625 167.285 133.795 167.475 ;
        RECT 138.685 167.305 138.855 167.495 ;
        RECT 139.155 167.330 139.315 167.440 ;
        RECT 140.525 167.285 140.695 167.475 ;
        RECT 144.205 167.305 144.375 167.495 ;
        RECT 146.045 167.285 146.215 167.475 ;
        RECT 147.885 167.305 148.055 167.495 ;
        RECT 148.800 167.335 148.920 167.445 ;
        RECT 150.185 167.285 150.355 167.495 ;
        RECT 11.125 166.475 12.495 167.285 ;
        RECT 12.505 166.475 18.015 167.285 ;
        RECT 18.025 166.475 23.535 167.285 ;
        RECT 23.545 166.475 25.375 167.285 ;
        RECT 25.955 166.605 29.420 167.285 ;
        RECT 29.985 166.605 32.725 167.285 ;
        RECT 28.500 166.375 29.420 166.605 ;
        RECT 32.745 166.505 34.115 167.285 ;
        RECT 34.125 166.475 36.875 167.285 ;
        RECT 36.895 166.415 37.325 167.200 ;
        RECT 37.345 166.475 41.015 167.285 ;
        RECT 41.125 166.375 44.235 167.285 ;
        RECT 44.245 166.475 49.755 167.285 ;
        RECT 49.765 166.475 51.595 167.285 ;
        RECT 52.065 166.375 53.880 167.285 ;
        RECT 53.905 166.475 59.415 167.285 ;
        RECT 59.425 166.475 62.175 167.285 ;
        RECT 62.655 166.415 63.085 167.200 ;
        RECT 63.215 166.605 66.680 167.285 ;
        RECT 65.760 166.375 66.680 166.605 ;
        RECT 66.805 166.375 68.155 167.285 ;
        RECT 68.165 166.505 69.535 167.285 ;
        RECT 69.545 166.475 73.215 167.285 ;
        RECT 73.685 166.605 76.425 167.285 ;
        RECT 76.640 166.375 80.115 167.285 ;
        RECT 80.125 166.475 85.635 167.285 ;
        RECT 85.645 166.475 88.395 167.285 ;
        RECT 88.415 166.415 88.845 167.200 ;
        RECT 88.865 166.475 91.615 167.285 ;
        RECT 91.665 166.375 94.835 167.285 ;
        RECT 94.860 166.375 96.675 167.285 ;
        RECT 96.685 166.475 100.355 167.285 ;
        RECT 101.300 166.375 103.115 167.285 ;
        RECT 103.125 166.475 106.795 167.285 ;
        RECT 107.725 166.605 111.625 167.285 ;
        RECT 107.725 166.375 108.655 166.605 ;
        RECT 111.865 166.375 113.695 167.285 ;
        RECT 114.175 166.415 114.605 167.200 ;
        RECT 114.625 166.475 118.295 167.285 ;
        RECT 118.305 166.605 120.135 167.285 ;
        RECT 118.790 166.375 120.135 166.605 ;
        RECT 120.145 166.475 123.815 167.285 ;
        RECT 123.825 166.475 125.195 167.285 ;
        RECT 125.345 166.375 127.955 167.285 ;
        RECT 127.965 166.475 133.475 167.285 ;
        RECT 133.485 166.475 138.995 167.285 ;
        RECT 139.935 166.415 140.365 167.200 ;
        RECT 140.385 166.475 145.895 167.285 ;
        RECT 145.905 166.475 148.655 167.285 ;
        RECT 149.125 166.475 150.495 167.285 ;
      LAYER nwell ;
        RECT 10.930 163.255 150.690 166.085 ;
      LAYER pwell ;
        RECT 11.125 162.055 12.495 162.865 ;
        RECT 12.505 162.055 16.175 162.865 ;
        RECT 19.700 162.735 20.610 162.955 ;
        RECT 22.145 162.735 23.915 162.965 ;
        RECT 16.185 162.055 23.915 162.735 ;
        RECT 24.015 162.140 24.445 162.925 ;
        RECT 24.465 162.055 28.135 162.865 ;
        RECT 29.165 162.055 32.275 162.965 ;
        RECT 32.385 162.055 35.495 162.965 ;
        RECT 35.505 162.055 37.335 162.865 ;
        RECT 37.805 162.735 38.940 162.965 ;
        RECT 44.225 162.735 45.155 162.965 ;
        RECT 37.805 162.055 41.015 162.735 ;
        RECT 41.485 162.055 45.155 162.735 ;
        RECT 45.165 162.055 46.535 162.865 ;
        RECT 46.645 162.055 49.755 162.965 ;
        RECT 49.775 162.140 50.205 162.925 ;
        RECT 50.225 162.055 51.595 162.865 ;
        RECT 51.895 162.055 54.815 162.965 ;
        RECT 54.825 162.055 58.035 162.965 ;
        RECT 58.045 162.055 63.555 162.865 ;
        RECT 63.565 162.055 66.315 162.865 ;
        RECT 66.785 162.765 67.715 162.965 ;
        RECT 69.045 162.765 69.995 162.965 ;
        RECT 66.785 162.285 69.995 162.765 ;
        RECT 66.930 162.085 69.995 162.285 ;
        RECT 11.265 161.845 11.435 162.055 ;
        RECT 12.645 161.845 12.815 162.055 ;
        RECT 16.325 161.865 16.495 162.055 ;
        RECT 18.165 161.845 18.335 162.035 ;
        RECT 21.845 161.845 22.015 162.035 ;
        RECT 23.225 161.845 23.395 162.035 ;
        RECT 24.605 161.865 24.775 162.055 ;
        RECT 28.295 161.900 28.455 162.010 ;
        RECT 29.205 161.865 29.375 162.055 ;
        RECT 31.045 161.845 31.215 162.035 ;
        RECT 32.425 161.865 32.595 162.055 ;
        RECT 35.645 161.865 35.815 162.055 ;
        RECT 37.485 162.005 37.655 162.035 ;
        RECT 36.560 161.895 36.680 162.005 ;
        RECT 37.480 161.895 37.655 162.005 ;
        RECT 11.125 161.035 12.495 161.845 ;
        RECT 12.505 161.035 18.015 161.845 ;
        RECT 18.025 161.035 21.695 161.845 ;
        RECT 21.705 161.035 23.075 161.845 ;
        RECT 23.085 161.165 30.815 161.845 ;
        RECT 26.600 160.945 27.510 161.165 ;
        RECT 29.045 160.935 30.815 161.165 ;
        RECT 30.905 161.035 36.415 161.845 ;
        RECT 36.895 160.975 37.325 161.760 ;
        RECT 37.485 161.615 37.655 161.895 ;
        RECT 40.705 161.865 40.875 162.055 ;
        RECT 41.160 161.895 41.280 162.005 ;
        RECT 41.625 161.845 41.795 162.055 ;
        RECT 43.460 161.895 43.580 162.005 ;
        RECT 44.845 161.845 45.015 162.035 ;
        RECT 45.305 161.845 45.475 162.055 ;
        RECT 46.685 161.865 46.855 162.055 ;
        RECT 48.995 161.890 49.155 162.000 ;
        RECT 38.765 161.615 41.475 161.845 ;
        RECT 37.380 161.165 41.475 161.615 ;
        RECT 37.380 160.935 38.755 161.165 ;
        RECT 40.525 160.935 41.475 161.165 ;
        RECT 41.485 161.035 43.315 161.845 ;
        RECT 43.795 160.935 45.145 161.845 ;
        RECT 45.165 161.035 48.835 161.845 ;
        RECT 49.910 161.815 50.080 162.035 ;
        RECT 50.365 161.865 50.535 162.055 ;
        RECT 53.585 161.845 53.755 162.035 ;
        RECT 54.500 161.865 54.670 162.055 ;
        RECT 54.965 161.865 55.135 162.055 ;
        RECT 58.185 161.865 58.355 162.055 ;
        RECT 62.325 161.845 62.495 162.035 ;
        RECT 63.705 161.865 63.875 162.055 ;
        RECT 64.165 161.845 64.335 162.035 ;
        RECT 64.625 161.845 64.795 162.035 ;
        RECT 66.005 161.845 66.175 162.035 ;
        RECT 66.460 161.895 66.580 162.005 ;
        RECT 66.930 161.865 67.100 162.085 ;
        RECT 69.060 162.055 69.995 162.085 ;
        RECT 70.315 162.735 71.245 162.965 ;
        RECT 74.595 162.735 75.515 162.965 ;
        RECT 70.315 162.055 72.150 162.735 ;
        RECT 73.225 162.055 75.515 162.735 ;
        RECT 75.535 162.140 75.965 162.925 ;
        RECT 85.225 162.735 86.575 162.965 ;
        RECT 88.110 162.735 89.020 162.955 ;
        RECT 92.855 162.735 93.785 162.965 ;
        RECT 75.985 162.055 85.090 162.735 ;
        RECT 85.225 162.055 92.535 162.735 ;
        RECT 92.855 162.055 94.690 162.735 ;
        RECT 94.865 162.055 96.215 162.965 ;
        RECT 96.225 162.055 99.895 162.865 ;
        RECT 99.905 162.055 101.275 162.865 ;
        RECT 101.295 162.140 101.725 162.925 ;
        RECT 101.745 162.055 105.415 162.865 ;
        RECT 105.905 162.055 107.255 162.965 ;
        RECT 107.265 162.055 112.775 162.865 ;
        RECT 112.785 162.055 118.295 162.865 ;
        RECT 118.305 162.055 123.815 162.865 ;
        RECT 123.825 162.055 126.575 162.865 ;
        RECT 127.055 162.140 127.485 162.925 ;
        RECT 127.505 162.055 133.015 162.865 ;
        RECT 133.025 162.055 138.535 162.865 ;
        RECT 138.545 162.055 144.055 162.865 ;
        RECT 144.065 162.055 147.735 162.865 ;
        RECT 147.745 162.055 149.115 162.865 ;
        RECT 149.125 162.055 150.495 162.865 ;
        RECT 71.985 162.035 72.150 162.055 ;
        RECT 69.680 161.895 69.800 162.005 ;
        RECT 71.985 161.865 72.155 162.035 ;
        RECT 72.455 161.900 72.615 162.010 ;
        RECT 73.365 161.845 73.535 162.055 ;
        RECT 73.830 161.845 74.000 162.035 ;
        RECT 76.125 161.865 76.295 162.055 ;
        RECT 52.485 161.815 53.435 161.845 ;
        RECT 49.765 161.135 53.435 161.815 ;
        RECT 52.485 160.935 53.435 161.135 ;
        RECT 53.445 161.035 55.275 161.845 ;
        RECT 55.325 161.165 62.635 161.845 ;
        RECT 55.325 160.935 56.675 161.165 ;
        RECT 58.210 160.945 59.120 161.165 ;
        RECT 62.655 160.975 63.085 161.760 ;
        RECT 63.105 161.065 64.475 161.845 ;
        RECT 64.485 161.035 65.855 161.845 ;
        RECT 65.945 160.935 69.395 161.845 ;
        RECT 70.100 161.165 73.565 161.845 ;
        RECT 70.100 160.935 71.020 161.165 ;
        RECT 73.685 160.935 76.605 161.845 ;
        RECT 77.050 161.815 77.220 162.035 ;
        RECT 80.270 161.845 80.440 162.035 ;
        RECT 83.485 161.845 83.655 162.035 ;
        RECT 84.865 161.845 85.035 162.035 ;
        RECT 92.225 161.845 92.395 162.055 ;
        RECT 94.525 162.035 94.690 162.055 ;
        RECT 92.685 161.845 92.855 162.035 ;
        RECT 94.525 161.865 94.695 162.035 ;
        RECT 94.980 161.865 95.150 162.055 ;
        RECT 96.365 162.005 96.535 162.055 ;
        RECT 96.360 161.895 96.535 162.005 ;
        RECT 96.365 161.865 96.535 161.895 ;
        RECT 96.825 161.845 96.995 162.035 ;
        RECT 100.045 161.865 100.215 162.055 ;
        RECT 101.885 161.865 102.055 162.055 ;
        RECT 104.185 161.845 104.355 162.035 ;
        RECT 105.560 161.895 105.680 162.005 ;
        RECT 106.020 161.895 106.140 162.005 ;
        RECT 106.485 161.845 106.655 162.035 ;
        RECT 106.940 161.865 107.110 162.055 ;
        RECT 107.405 161.865 107.575 162.055 ;
        RECT 112.925 161.865 113.095 162.055 ;
        RECT 114.765 161.845 114.935 162.035 ;
        RECT 118.445 161.865 118.615 162.055 ;
        RECT 120.285 161.845 120.455 162.035 ;
        RECT 123.965 161.865 124.135 162.055 ;
        RECT 125.805 161.845 125.975 162.035 ;
        RECT 126.720 161.895 126.840 162.005 ;
        RECT 127.645 161.865 127.815 162.055 ;
        RECT 131.325 161.845 131.495 162.035 ;
        RECT 133.165 161.865 133.335 162.055 ;
        RECT 136.845 161.845 137.015 162.035 ;
        RECT 138.685 161.865 138.855 162.055 ;
        RECT 139.600 161.895 139.720 162.005 ;
        RECT 140.525 161.845 140.695 162.035 ;
        RECT 144.205 161.865 144.375 162.055 ;
        RECT 146.045 161.845 146.215 162.035 ;
        RECT 147.885 161.865 148.055 162.055 ;
        RECT 148.800 161.895 148.920 162.005 ;
        RECT 150.185 161.845 150.355 162.055 ;
        RECT 79.180 161.815 80.115 161.845 ;
        RECT 77.050 161.615 80.115 161.815 ;
        RECT 76.905 161.135 80.115 161.615 ;
        RECT 76.905 160.935 77.835 161.135 ;
        RECT 79.165 160.935 80.115 161.135 ;
        RECT 80.125 160.935 83.045 161.845 ;
        RECT 83.345 161.065 84.715 161.845 ;
        RECT 84.725 161.035 88.395 161.845 ;
        RECT 88.415 160.975 88.845 161.760 ;
        RECT 88.960 161.165 92.425 161.845 ;
        RECT 88.960 160.935 89.880 161.165 ;
        RECT 92.545 161.035 96.215 161.845 ;
        RECT 96.685 161.165 103.995 161.845 ;
        RECT 100.200 160.945 101.110 161.165 ;
        RECT 102.645 160.935 103.995 161.165 ;
        RECT 104.045 161.035 105.875 161.845 ;
        RECT 106.345 161.165 114.075 161.845 ;
        RECT 109.860 160.945 110.770 161.165 ;
        RECT 112.305 160.935 114.075 161.165 ;
        RECT 114.175 160.975 114.605 161.760 ;
        RECT 114.625 161.035 120.135 161.845 ;
        RECT 120.145 161.035 125.655 161.845 ;
        RECT 125.665 161.035 131.175 161.845 ;
        RECT 131.185 161.035 136.695 161.845 ;
        RECT 136.705 161.035 139.455 161.845 ;
        RECT 139.935 160.975 140.365 161.760 ;
        RECT 140.385 161.035 145.895 161.845 ;
        RECT 145.905 161.035 148.655 161.845 ;
        RECT 149.125 161.035 150.495 161.845 ;
      LAYER nwell ;
        RECT 10.930 157.815 150.690 160.645 ;
      LAYER pwell ;
        RECT 11.125 156.615 12.495 157.425 ;
        RECT 12.505 156.615 18.015 157.425 ;
        RECT 18.025 156.615 23.535 157.425 ;
        RECT 24.015 156.700 24.445 157.485 ;
        RECT 25.605 157.435 26.555 157.525 ;
        RECT 24.625 156.615 26.555 157.435 ;
        RECT 26.765 156.615 28.135 157.395 ;
        RECT 28.145 156.615 33.655 157.425 ;
        RECT 33.665 156.615 39.175 157.425 ;
        RECT 39.185 156.615 44.695 157.425 ;
        RECT 44.705 156.615 48.375 157.425 ;
        RECT 48.385 156.615 49.755 157.425 ;
        RECT 49.775 156.700 50.205 157.485 ;
        RECT 52.300 157.295 53.435 157.525 ;
        RECT 50.225 156.615 53.435 157.295 ;
        RECT 53.445 156.615 56.195 157.425 ;
        RECT 58.035 157.295 58.955 157.525 ;
        RECT 71.125 157.435 72.075 157.525 ;
        RECT 56.665 156.615 58.955 157.295 ;
        RECT 58.965 156.615 64.475 157.425 ;
        RECT 64.485 156.615 69.995 157.425 ;
        RECT 71.125 156.615 73.055 157.435 ;
        RECT 74.595 157.295 75.515 157.525 ;
        RECT 73.225 156.615 75.515 157.295 ;
        RECT 75.535 156.700 75.965 157.485 ;
        RECT 75.985 156.615 77.355 157.425 ;
        RECT 77.405 156.615 80.575 157.525 ;
        RECT 80.585 156.615 84.255 157.425 ;
        RECT 84.285 156.615 85.635 157.525 ;
        RECT 85.645 156.615 89.300 157.525 ;
        RECT 90.375 157.295 91.305 157.525 ;
        RECT 89.470 156.615 91.305 157.295 ;
        RECT 91.625 156.615 93.455 157.425 ;
        RECT 93.465 156.615 96.940 157.525 ;
        RECT 97.145 156.615 100.065 157.525 ;
        RECT 101.295 156.700 101.725 157.485 ;
        RECT 101.745 156.615 104.855 157.525 ;
        RECT 104.965 156.615 108.635 157.425 ;
        RECT 109.565 156.615 112.305 157.295 ;
        RECT 112.325 156.615 117.835 157.425 ;
        RECT 117.845 156.615 123.355 157.425 ;
        RECT 123.365 156.615 127.035 157.425 ;
        RECT 127.055 156.700 127.485 157.485 ;
        RECT 127.505 156.615 133.015 157.425 ;
        RECT 133.025 156.615 138.535 157.425 ;
        RECT 138.545 156.615 144.055 157.425 ;
        RECT 144.065 156.615 147.735 157.425 ;
        RECT 147.745 156.615 149.115 157.425 ;
        RECT 149.125 156.615 150.495 157.425 ;
        RECT 11.265 156.405 11.435 156.615 ;
        RECT 12.645 156.405 12.815 156.615 ;
        RECT 18.165 156.425 18.335 156.615 ;
        RECT 24.625 156.595 24.775 156.615 ;
        RECT 19.085 156.405 19.255 156.595 ;
        RECT 19.545 156.405 19.715 156.595 ;
        RECT 23.680 156.455 23.800 156.565 ;
        RECT 24.605 156.425 24.775 156.595 ;
        RECT 25.065 156.405 25.235 156.595 ;
        RECT 27.825 156.425 27.995 156.615 ;
        RECT 28.285 156.425 28.455 156.615 ;
        RECT 28.740 156.455 28.860 156.565 ;
        RECT 31.965 156.405 32.135 156.595 ;
        RECT 32.425 156.405 32.595 156.595 ;
        RECT 33.805 156.405 33.975 156.615 ;
        RECT 37.485 156.405 37.655 156.595 ;
        RECT 38.870 156.405 39.040 156.595 ;
        RECT 39.325 156.425 39.495 156.615 ;
        RECT 43.925 156.405 44.095 156.595 ;
        RECT 44.385 156.425 44.555 156.595 ;
        RECT 44.845 156.425 45.015 156.615 ;
        RECT 48.525 156.425 48.695 156.615 ;
        RECT 50.365 156.425 50.535 156.615 ;
        RECT 53.585 156.425 53.755 156.615 ;
        RECT 44.395 156.405 44.555 156.425 ;
        RECT 54.045 156.405 54.215 156.595 ;
        RECT 54.505 156.405 54.675 156.595 ;
        RECT 56.340 156.405 56.510 156.595 ;
        RECT 56.805 156.425 56.975 156.615 ;
        RECT 57.725 156.405 57.895 156.595 ;
        RECT 59.105 156.405 59.275 156.615 ;
        RECT 60.485 156.405 60.655 156.595 ;
        RECT 62.320 156.455 62.440 156.565 ;
        RECT 63.255 156.450 63.415 156.560 ;
        RECT 64.165 156.405 64.335 156.595 ;
        RECT 64.625 156.425 64.795 156.615 ;
        RECT 72.905 156.595 73.055 156.615 ;
        RECT 70.155 156.460 70.315 156.570 ;
        RECT 71.980 156.455 72.100 156.565 ;
        RECT 72.450 156.405 72.620 156.595 ;
        RECT 72.905 156.425 73.075 156.595 ;
        RECT 73.365 156.425 73.535 156.615 ;
        RECT 74.285 156.405 74.455 156.595 ;
        RECT 76.125 156.425 76.295 156.615 ;
        RECT 77.505 156.425 77.675 156.615 ;
        RECT 79.805 156.405 79.975 156.595 ;
        RECT 80.725 156.425 80.895 156.615 ;
        RECT 83.485 156.405 83.655 156.595 ;
        RECT 84.400 156.425 84.570 156.615 ;
        RECT 85.790 156.595 85.960 156.615 ;
        RECT 89.470 156.595 89.635 156.615 ;
        RECT 85.785 156.425 85.960 156.595 ;
        RECT 85.785 156.405 85.955 156.425 ;
        RECT 88.080 156.405 88.250 156.595 ;
        RECT 89.005 156.405 89.175 156.595 ;
        RECT 89.465 156.425 89.635 156.595 ;
        RECT 91.765 156.425 91.935 156.615 ;
        RECT 92.685 156.405 92.855 156.595 ;
        RECT 93.610 156.425 93.780 156.615 ;
        RECT 97.290 156.425 97.460 156.615 ;
        RECT 11.125 155.595 12.495 156.405 ;
        RECT 12.505 155.595 18.015 156.405 ;
        RECT 18.025 155.625 19.395 156.405 ;
        RECT 19.405 155.595 24.915 156.405 ;
        RECT 24.925 155.595 28.595 156.405 ;
        RECT 29.065 155.495 32.275 156.405 ;
        RECT 32.285 155.595 33.655 156.405 ;
        RECT 33.765 155.495 36.875 156.405 ;
        RECT 36.895 155.535 37.325 156.320 ;
        RECT 37.345 155.595 38.715 156.405 ;
        RECT 38.725 155.495 41.475 156.405 ;
        RECT 41.495 155.495 44.225 156.405 ;
        RECT 44.395 155.495 48.050 156.405 ;
        RECT 48.535 155.495 54.355 156.405 ;
        RECT 54.365 155.595 56.195 156.405 ;
        RECT 56.225 155.495 57.575 156.405 ;
        RECT 57.585 155.595 58.955 156.405 ;
        RECT 58.965 155.625 60.335 156.405 ;
        RECT 60.345 155.595 62.175 156.405 ;
        RECT 62.655 155.535 63.085 156.320 ;
        RECT 64.025 155.725 71.755 156.405 ;
        RECT 67.540 155.505 68.450 155.725 ;
        RECT 69.985 155.495 71.755 155.725 ;
        RECT 72.305 155.495 74.135 156.405 ;
        RECT 74.145 155.595 79.655 156.405 ;
        RECT 79.665 155.595 83.335 156.405 ;
        RECT 83.345 155.725 85.635 156.405 ;
        RECT 84.715 155.495 85.635 155.725 ;
        RECT 85.645 155.595 87.015 156.405 ;
        RECT 87.045 155.495 88.395 156.405 ;
        RECT 88.415 155.535 88.845 156.320 ;
        RECT 88.865 155.595 92.535 156.405 ;
        RECT 92.545 155.725 96.215 156.405 ;
        RECT 95.285 155.495 96.215 155.725 ;
        RECT 96.225 156.375 97.160 156.405 ;
        RECT 99.120 156.375 99.290 156.595 ;
        RECT 99.595 156.450 99.755 156.560 ;
        RECT 100.515 156.460 100.675 156.570 ;
        RECT 102.345 156.405 102.515 156.595 ;
        RECT 102.805 156.405 102.975 156.595 ;
        RECT 104.645 156.425 104.815 156.615 ;
        RECT 105.105 156.425 105.275 156.615 ;
        RECT 108.795 156.460 108.955 156.570 ;
        RECT 109.250 156.405 109.420 156.595 ;
        RECT 109.705 156.405 109.875 156.615 ;
        RECT 112.465 156.425 112.635 156.615 ;
        RECT 113.395 156.450 113.555 156.560 ;
        RECT 114.765 156.405 114.935 156.595 ;
        RECT 117.985 156.425 118.155 156.615 ;
        RECT 120.285 156.405 120.455 156.595 ;
        RECT 123.505 156.425 123.675 156.615 ;
        RECT 125.805 156.405 125.975 156.595 ;
        RECT 127.645 156.425 127.815 156.615 ;
        RECT 131.325 156.405 131.495 156.595 ;
        RECT 133.165 156.425 133.335 156.615 ;
        RECT 136.845 156.405 137.015 156.595 ;
        RECT 138.685 156.425 138.855 156.615 ;
        RECT 139.600 156.455 139.720 156.565 ;
        RECT 140.525 156.405 140.695 156.595 ;
        RECT 144.205 156.425 144.375 156.615 ;
        RECT 146.045 156.405 146.215 156.595 ;
        RECT 147.885 156.425 148.055 156.615 ;
        RECT 148.800 156.455 148.920 156.565 ;
        RECT 150.185 156.405 150.355 156.615 ;
        RECT 96.225 156.175 99.290 156.375 ;
        RECT 96.225 155.695 99.435 156.175 ;
        RECT 96.225 155.495 97.175 155.695 ;
        RECT 98.505 155.495 99.435 155.695 ;
        RECT 100.365 155.725 102.655 156.405 ;
        RECT 100.365 155.495 101.285 155.725 ;
        RECT 102.665 155.595 108.175 156.405 ;
        RECT 108.185 155.495 109.535 156.405 ;
        RECT 109.565 155.595 113.235 156.405 ;
        RECT 114.175 155.535 114.605 156.320 ;
        RECT 114.625 155.595 120.135 156.405 ;
        RECT 120.145 155.595 125.655 156.405 ;
        RECT 125.665 155.595 131.175 156.405 ;
        RECT 131.185 155.595 136.695 156.405 ;
        RECT 136.705 155.595 139.455 156.405 ;
        RECT 139.935 155.535 140.365 156.320 ;
        RECT 140.385 155.595 145.895 156.405 ;
        RECT 145.905 155.595 148.655 156.405 ;
        RECT 149.125 155.595 150.495 156.405 ;
      LAYER nwell ;
        RECT 10.930 152.375 150.690 155.205 ;
      LAYER pwell ;
        RECT 11.125 151.175 12.495 151.985 ;
        RECT 12.505 151.175 15.255 151.985 ;
        RECT 19.240 151.855 20.150 152.075 ;
        RECT 21.685 151.855 23.035 152.085 ;
        RECT 15.725 151.175 23.035 151.855 ;
        RECT 24.015 151.260 24.445 152.045 ;
        RECT 24.565 151.175 27.675 152.085 ;
        RECT 27.685 151.175 29.515 151.985 ;
        RECT 29.525 151.175 32.735 152.085 ;
        RECT 32.745 151.175 38.255 151.985 ;
        RECT 38.265 151.175 41.015 151.985 ;
        RECT 41.485 151.175 43.315 152.085 ;
        RECT 44.265 151.175 45.615 152.085 ;
        RECT 45.625 151.175 49.295 151.985 ;
        RECT 49.775 151.260 50.205 152.045 ;
        RECT 50.225 151.175 52.055 151.985 ;
        RECT 52.525 151.175 55.735 152.085 ;
        RECT 55.745 151.175 57.115 151.985 ;
        RECT 57.205 151.855 58.975 152.085 ;
        RECT 60.510 151.855 61.420 152.075 ;
        RECT 64.955 151.995 66.545 152.085 ;
        RECT 57.205 151.175 64.935 151.855 ;
        RECT 64.955 151.175 67.525 151.995 ;
        RECT 67.705 151.175 71.375 151.985 ;
        RECT 71.855 151.175 74.585 152.085 ;
        RECT 75.535 151.260 75.965 152.045 ;
        RECT 75.995 151.175 77.345 152.085 ;
        RECT 77.465 151.175 80.575 152.085 ;
        RECT 80.585 151.175 83.335 151.985 ;
        RECT 83.805 151.175 85.635 152.085 ;
        RECT 85.645 151.175 87.460 152.085 ;
        RECT 87.485 151.175 91.155 151.985 ;
        RECT 92.085 151.175 95.560 152.085 ;
        RECT 95.765 151.885 96.715 152.085 ;
        RECT 95.765 151.205 99.435 151.885 ;
        RECT 95.765 151.175 96.715 151.205 ;
        RECT 11.265 150.965 11.435 151.175 ;
        RECT 12.645 150.965 12.815 151.175 ;
        RECT 15.400 151.015 15.520 151.125 ;
        RECT 15.865 150.985 16.035 151.175 ;
        RECT 18.175 151.010 18.335 151.120 ;
        RECT 20.925 150.985 21.095 151.155 ;
        RECT 20.925 150.965 21.075 150.985 ;
        RECT 21.385 150.965 21.555 151.155 ;
        RECT 23.235 151.020 23.395 151.130 ;
        RECT 24.605 150.985 24.775 151.175 ;
        RECT 26.905 150.965 27.075 151.155 ;
        RECT 27.825 150.985 27.995 151.175 ;
        RECT 30.585 150.965 30.755 151.155 ;
        RECT 32.425 150.985 32.595 151.175 ;
        RECT 32.885 150.985 33.055 151.175 ;
        RECT 34.725 150.965 34.895 151.155 ;
        RECT 35.185 150.965 35.355 151.155 ;
        RECT 37.485 150.965 37.655 151.155 ;
        RECT 38.405 150.985 38.575 151.175 ;
        RECT 38.860 150.965 39.030 151.155 ;
        RECT 40.255 151.010 40.415 151.120 ;
        RECT 41.160 150.965 41.330 151.155 ;
        RECT 42.545 150.965 42.715 151.155 ;
        RECT 43.000 150.985 43.170 151.175 ;
        RECT 43.475 151.020 43.635 151.130 ;
        RECT 44.380 150.985 44.550 151.175 ;
        RECT 45.765 150.985 45.935 151.175 ;
        RECT 48.065 150.965 48.235 151.155 ;
        RECT 49.440 151.015 49.560 151.125 ;
        RECT 50.365 150.985 50.535 151.175 ;
        RECT 50.820 151.015 50.940 151.125 ;
        RECT 51.285 150.985 51.455 151.155 ;
        RECT 52.200 151.015 52.320 151.125 ;
        RECT 51.285 150.965 51.485 150.985 ;
        RECT 54.965 150.965 55.135 151.155 ;
        RECT 55.435 150.985 55.605 151.175 ;
        RECT 55.885 150.985 56.055 151.175 ;
        RECT 60.485 150.965 60.655 151.155 ;
        RECT 62.320 151.015 62.440 151.125 ;
        RECT 63.245 150.965 63.415 151.155 ;
        RECT 64.625 150.985 64.795 151.175 ;
        RECT 67.385 151.155 67.525 151.175 ;
        RECT 67.385 150.985 67.555 151.155 ;
        RECT 67.845 150.985 68.015 151.175 ;
        RECT 68.765 150.965 68.935 151.155 ;
        RECT 71.520 151.015 71.640 151.125 ;
        RECT 71.985 150.985 72.155 151.175 ;
        RECT 74.280 151.015 74.400 151.125 ;
        RECT 74.755 151.020 74.915 151.130 ;
        RECT 76.120 150.965 76.290 151.155 ;
        RECT 76.585 150.965 76.755 151.155 ;
        RECT 77.045 150.985 77.215 151.175 ;
        RECT 77.505 150.985 77.675 151.175 ;
        RECT 80.725 150.985 80.895 151.175 ;
        RECT 82.105 150.965 82.275 151.155 ;
        RECT 83.480 151.015 83.600 151.125 ;
        RECT 85.320 150.985 85.490 151.175 ;
        RECT 87.165 150.985 87.335 151.175 ;
        RECT 87.625 150.985 87.795 151.175 ;
        RECT 89.005 150.965 89.175 151.155 ;
        RECT 91.315 151.020 91.475 151.130 ;
        RECT 92.230 150.985 92.400 151.175 ;
        RECT 92.680 151.015 92.800 151.125 ;
        RECT 93.150 150.965 93.320 151.155 ;
        RECT 98.200 150.965 98.370 151.155 ;
        RECT 98.665 150.965 98.835 151.155 ;
        RECT 99.120 150.985 99.290 151.205 ;
        RECT 99.445 151.175 101.275 151.985 ;
        RECT 101.295 151.260 101.725 152.045 ;
        RECT 110.985 151.855 112.335 152.085 ;
        RECT 113.870 151.855 114.780 152.075 ;
        RECT 101.745 151.175 110.850 151.855 ;
        RECT 110.985 151.175 118.295 151.855 ;
        RECT 118.305 151.175 123.815 151.985 ;
        RECT 123.825 151.175 126.575 151.985 ;
        RECT 127.055 151.260 127.485 152.045 ;
        RECT 127.505 151.175 133.015 151.985 ;
        RECT 133.025 151.175 138.535 151.985 ;
        RECT 138.545 151.175 144.055 151.985 ;
        RECT 144.065 151.175 147.735 151.985 ;
        RECT 147.745 151.175 149.115 151.985 ;
        RECT 149.125 151.175 150.495 151.985 ;
        RECT 99.585 150.985 99.755 151.175 ;
        RECT 101.420 151.015 101.540 151.125 ;
        RECT 101.885 150.985 102.055 151.175 ;
        RECT 104.645 150.965 104.815 151.155 ;
        RECT 105.115 151.010 105.275 151.120 ;
        RECT 109.240 150.965 109.410 151.155 ;
        RECT 112.470 150.965 112.640 151.155 ;
        RECT 112.925 150.965 113.095 151.155 ;
        RECT 114.765 150.965 114.935 151.155 ;
        RECT 117.985 150.985 118.155 151.175 ;
        RECT 118.445 150.985 118.615 151.175 ;
        RECT 123.505 150.965 123.675 151.155 ;
        RECT 123.965 150.965 124.135 151.175 ;
        RECT 126.720 151.015 126.840 151.125 ;
        RECT 127.645 150.985 127.815 151.175 ;
        RECT 129.485 150.965 129.655 151.155 ;
        RECT 133.165 150.985 133.335 151.175 ;
        RECT 135.005 150.965 135.175 151.155 ;
        RECT 138.685 150.965 138.855 151.175 ;
        RECT 140.525 150.965 140.695 151.155 ;
        RECT 144.205 150.985 144.375 151.175 ;
        RECT 146.045 150.965 146.215 151.155 ;
        RECT 147.885 150.985 148.055 151.175 ;
        RECT 148.800 151.015 148.920 151.125 ;
        RECT 150.185 150.965 150.355 151.175 ;
        RECT 11.125 150.155 12.495 150.965 ;
        RECT 12.505 150.155 18.015 150.965 ;
        RECT 19.145 150.145 21.075 150.965 ;
        RECT 21.245 150.155 26.755 150.965 ;
        RECT 26.765 150.155 30.435 150.965 ;
        RECT 30.445 150.155 31.815 150.965 ;
        RECT 19.145 150.055 20.095 150.145 ;
        RECT 31.825 150.055 34.935 150.965 ;
        RECT 35.045 150.155 36.875 150.965 ;
        RECT 36.895 150.095 37.325 150.880 ;
        RECT 37.345 150.155 38.715 150.965 ;
        RECT 38.745 150.055 40.095 150.965 ;
        RECT 41.045 150.055 42.395 150.965 ;
        RECT 42.405 150.155 47.915 150.965 ;
        RECT 47.925 150.155 50.675 150.965 ;
        RECT 51.285 150.285 54.815 150.965 ;
        RECT 51.990 150.055 54.815 150.285 ;
        RECT 54.825 150.155 60.335 150.965 ;
        RECT 60.345 150.155 62.175 150.965 ;
        RECT 62.655 150.095 63.085 150.880 ;
        RECT 63.105 150.155 68.615 150.965 ;
        RECT 68.625 150.155 74.135 150.965 ;
        RECT 74.605 150.055 76.435 150.965 ;
        RECT 76.445 150.155 81.955 150.965 ;
        RECT 81.965 150.155 87.475 150.965 ;
        RECT 88.415 150.095 88.845 150.880 ;
        RECT 88.865 150.155 92.535 150.965 ;
        RECT 93.005 150.055 96.660 150.965 ;
        RECT 96.685 150.055 98.515 150.965 ;
        RECT 98.525 150.155 101.275 150.965 ;
        RECT 101.745 150.055 104.915 150.965 ;
        RECT 106.080 150.055 109.555 150.965 ;
        RECT 109.565 150.055 112.765 150.965 ;
        RECT 112.795 150.055 114.145 150.965 ;
        RECT 114.175 150.095 114.605 150.880 ;
        RECT 114.625 150.185 115.995 150.965 ;
        RECT 116.085 150.285 123.815 150.965 ;
        RECT 116.085 150.055 117.855 150.285 ;
        RECT 119.390 150.065 120.300 150.285 ;
        RECT 123.825 150.155 129.335 150.965 ;
        RECT 129.345 150.155 134.855 150.965 ;
        RECT 134.865 150.155 138.535 150.965 ;
        RECT 138.545 150.155 139.915 150.965 ;
        RECT 139.935 150.095 140.365 150.880 ;
        RECT 140.385 150.155 145.895 150.965 ;
        RECT 145.905 150.155 148.655 150.965 ;
        RECT 149.125 150.155 150.495 150.965 ;
      LAYER nwell ;
        RECT 10.930 146.935 150.690 149.765 ;
      LAYER pwell ;
        RECT 11.125 145.735 12.495 146.545 ;
        RECT 12.505 145.735 18.015 146.545 ;
        RECT 20.305 146.415 21.235 146.645 ;
        RECT 23.065 146.415 23.995 146.645 ;
        RECT 18.485 145.735 21.235 146.415 ;
        RECT 21.245 145.735 23.995 146.415 ;
        RECT 24.015 145.820 24.445 146.605 ;
        RECT 24.485 145.735 25.835 146.645 ;
        RECT 26.135 145.735 29.055 146.645 ;
        RECT 29.145 145.735 32.595 146.645 ;
        RECT 32.745 145.735 36.415 146.545 ;
        RECT 36.425 145.735 37.795 146.545 ;
        RECT 41.320 146.415 42.230 146.635 ;
        RECT 43.765 146.415 45.115 146.645 ;
        RECT 37.805 145.735 45.115 146.415 ;
        RECT 45.935 146.415 46.865 146.645 ;
        RECT 48.410 146.415 49.755 146.645 ;
        RECT 45.935 145.735 47.770 146.415 ;
        RECT 47.925 145.735 49.755 146.415 ;
        RECT 49.775 145.820 50.205 146.605 ;
        RECT 50.705 145.735 52.055 146.645 ;
        RECT 52.065 145.735 54.815 146.645 ;
        RECT 55.785 145.735 58.955 146.645 ;
        RECT 59.425 145.735 61.240 146.645 ;
        RECT 61.265 146.415 62.185 146.645 ;
        RECT 61.265 145.735 64.850 146.415 ;
        RECT 64.945 145.735 67.865 146.645 ;
        RECT 68.625 145.735 71.835 146.645 ;
        RECT 71.845 145.735 75.515 146.545 ;
        RECT 75.535 145.820 75.965 146.605 ;
        RECT 76.905 145.735 79.645 146.415 ;
        RECT 79.665 145.735 83.140 146.645 ;
        RECT 83.345 145.735 85.175 146.545 ;
        RECT 85.745 145.735 88.855 146.645 ;
        RECT 88.865 145.735 94.375 146.545 ;
        RECT 94.385 145.735 98.055 146.545 ;
        RECT 98.065 145.735 99.435 146.545 ;
        RECT 99.455 145.735 100.805 146.645 ;
        RECT 101.295 145.820 101.725 146.605 ;
        RECT 101.745 145.735 107.585 146.645 ;
        RECT 107.725 145.735 109.075 146.645 ;
        RECT 109.665 145.735 112.775 146.645 ;
        RECT 113.245 145.735 116.455 146.645 ;
        RECT 116.665 146.555 117.615 146.645 ;
        RECT 116.665 145.735 118.595 146.555 ;
        RECT 118.765 145.735 124.275 146.545 ;
        RECT 124.285 145.735 127.035 146.545 ;
        RECT 127.055 145.820 127.485 146.605 ;
        RECT 127.505 145.735 133.015 146.545 ;
        RECT 133.025 145.735 138.535 146.545 ;
        RECT 138.545 145.735 144.055 146.545 ;
        RECT 144.065 145.735 147.735 146.545 ;
        RECT 147.745 145.735 149.115 146.545 ;
        RECT 149.125 145.735 150.495 146.545 ;
        RECT 11.265 145.525 11.435 145.735 ;
        RECT 12.645 145.525 12.815 145.735 ;
        RECT 18.165 145.685 18.335 145.715 ;
        RECT 18.160 145.575 18.335 145.685 ;
        RECT 18.165 145.525 18.335 145.575 ;
        RECT 18.625 145.545 18.795 145.735 ;
        RECT 21.385 145.545 21.555 145.735 ;
        RECT 23.680 145.575 23.800 145.685 ;
        RECT 24.145 145.525 24.315 145.715 ;
        RECT 25.520 145.545 25.690 145.735 ;
        RECT 25.980 145.575 26.100 145.685 ;
        RECT 26.445 145.525 26.615 145.715 ;
        RECT 28.740 145.545 28.910 145.735 ;
        RECT 29.205 145.545 29.375 145.735 ;
        RECT 29.665 145.525 29.835 145.715 ;
        RECT 32.885 145.545 33.055 145.735 ;
        RECT 35.185 145.525 35.355 145.715 ;
        RECT 36.565 145.545 36.735 145.735 ;
        RECT 37.485 145.545 37.655 145.715 ;
        RECT 37.945 145.545 38.115 145.735 ;
        RECT 47.605 145.715 47.770 145.735 ;
        RECT 37.505 145.525 37.655 145.545 ;
        RECT 40.705 145.525 40.875 145.715 ;
        RECT 41.165 145.525 41.335 145.715 ;
        RECT 45.300 145.575 45.420 145.685 ;
        RECT 46.685 145.525 46.855 145.715 ;
        RECT 47.605 145.545 47.775 145.715 ;
        RECT 48.065 145.545 48.235 145.735 ;
        RECT 50.360 145.575 50.480 145.685 ;
        RECT 51.740 145.545 51.910 145.735 ;
        RECT 53.125 145.525 53.295 145.715 ;
        RECT 53.585 145.525 53.755 145.715 ;
        RECT 54.505 145.545 54.675 145.735 ;
        RECT 54.975 145.580 55.135 145.690 ;
        RECT 55.885 145.545 56.055 145.735 ;
        RECT 59.105 145.685 59.275 145.715 ;
        RECT 59.100 145.575 59.275 145.685 ;
        RECT 59.105 145.525 59.275 145.575 ;
        RECT 60.485 145.545 60.655 145.715 ;
        RECT 60.945 145.545 61.115 145.735 ;
        RECT 61.410 145.545 61.580 145.735 ;
        RECT 63.240 145.575 63.360 145.685 ;
        RECT 60.505 145.525 60.655 145.545 ;
        RECT 63.705 145.525 63.875 145.715 ;
        RECT 65.090 145.545 65.260 145.735 ;
        RECT 68.300 145.575 68.420 145.685 ;
        RECT 68.755 145.545 68.925 145.735 ;
        RECT 71.065 145.525 71.235 145.715 ;
        RECT 71.985 145.545 72.155 145.735 ;
        RECT 76.135 145.580 76.295 145.690 ;
        RECT 77.045 145.545 77.215 145.735 ;
        RECT 79.810 145.715 79.980 145.735 ;
        RECT 79.800 145.545 79.980 145.715 ;
        RECT 79.800 145.525 79.970 145.545 ;
        RECT 80.265 145.525 80.435 145.715 ;
        RECT 83.485 145.545 83.655 145.735 ;
        RECT 83.945 145.545 84.115 145.715 ;
        RECT 83.945 145.525 84.110 145.545 ;
        RECT 84.405 145.525 84.575 145.715 ;
        RECT 85.320 145.575 85.440 145.685 ;
        RECT 85.785 145.545 85.955 145.735 ;
        RECT 88.085 145.525 88.255 145.715 ;
        RECT 89.005 145.545 89.175 145.735 ;
        RECT 90.845 145.545 91.015 145.715 ;
        RECT 91.315 145.570 91.475 145.680 ;
        RECT 90.845 145.525 90.995 145.545 ;
        RECT 92.225 145.525 92.395 145.715 ;
        RECT 94.525 145.545 94.695 145.735 ;
        RECT 95.445 145.525 95.615 145.715 ;
        RECT 98.205 145.545 98.375 145.735 ;
        RECT 99.585 145.545 99.755 145.735 ;
        RECT 100.965 145.685 101.135 145.715 ;
        RECT 100.960 145.575 101.135 145.685 ;
        RECT 100.965 145.525 101.135 145.575 ;
        RECT 101.885 145.545 102.055 145.735 ;
        RECT 102.805 145.525 102.975 145.715 ;
        RECT 105.565 145.525 105.735 145.715 ;
        RECT 108.790 145.545 108.960 145.735 ;
        RECT 109.240 145.575 109.360 145.685 ;
        RECT 109.705 145.545 109.875 145.735 ;
        RECT 111.085 145.525 111.255 145.715 ;
        RECT 112.920 145.575 113.040 145.685 ;
        RECT 113.385 145.545 113.555 145.735 ;
        RECT 118.445 145.715 118.595 145.735 ;
        RECT 113.840 145.575 113.960 145.685 ;
        RECT 114.775 145.570 114.935 145.680 ;
        RECT 115.685 145.525 115.855 145.715 ;
        RECT 117.065 145.525 117.235 145.715 ;
        RECT 118.445 145.545 118.615 145.715 ;
        RECT 118.905 145.545 119.075 145.735 ;
        RECT 122.585 145.525 122.755 145.715 ;
        RECT 124.425 145.545 124.595 145.735 ;
        RECT 127.645 145.545 127.815 145.735 ;
        RECT 128.105 145.525 128.275 145.715 ;
        RECT 133.165 145.545 133.335 145.735 ;
        RECT 133.625 145.525 133.795 145.715 ;
        RECT 138.685 145.545 138.855 145.735 ;
        RECT 139.155 145.570 139.315 145.680 ;
        RECT 140.525 145.525 140.695 145.715 ;
        RECT 144.205 145.545 144.375 145.735 ;
        RECT 146.045 145.525 146.215 145.715 ;
        RECT 147.885 145.545 148.055 145.735 ;
        RECT 148.800 145.575 148.920 145.685 ;
        RECT 150.185 145.525 150.355 145.735 ;
        RECT 11.125 144.715 12.495 145.525 ;
        RECT 12.505 144.715 18.015 145.525 ;
        RECT 18.025 144.715 23.535 145.525 ;
        RECT 24.020 144.615 25.835 145.525 ;
        RECT 26.345 144.615 29.515 145.525 ;
        RECT 29.525 144.715 35.035 145.525 ;
        RECT 35.045 144.715 36.875 145.525 ;
        RECT 36.895 144.655 37.325 145.440 ;
        RECT 37.505 144.705 39.435 145.525 ;
        RECT 39.645 144.745 41.015 145.525 ;
        RECT 41.025 144.715 46.535 145.525 ;
        RECT 46.545 144.715 50.215 145.525 ;
        RECT 50.685 145.295 53.295 145.525 ;
        RECT 38.485 144.615 39.435 144.705 ;
        RECT 50.685 144.615 53.435 145.295 ;
        RECT 53.445 144.715 58.955 145.525 ;
        RECT 58.965 144.715 60.335 145.525 ;
        RECT 60.505 144.705 62.435 145.525 ;
        RECT 61.485 144.615 62.435 144.705 ;
        RECT 62.655 144.655 63.085 145.440 ;
        RECT 63.565 144.845 70.875 145.525 ;
        RECT 70.925 144.845 78.235 145.525 ;
        RECT 67.080 144.625 67.990 144.845 ;
        RECT 69.525 144.615 70.875 144.845 ;
        RECT 74.440 144.625 75.350 144.845 ;
        RECT 76.885 144.615 78.235 144.845 ;
        RECT 78.345 144.615 80.115 145.525 ;
        RECT 80.125 144.715 81.955 145.525 ;
        RECT 82.275 144.845 84.110 145.525 ;
        RECT 82.275 144.615 83.205 144.845 ;
        RECT 84.265 144.715 86.095 145.525 ;
        RECT 86.105 144.845 88.395 145.525 ;
        RECT 86.105 144.615 87.025 144.845 ;
        RECT 88.415 144.655 88.845 145.440 ;
        RECT 89.065 144.705 90.995 145.525 ;
        RECT 89.065 144.615 90.015 144.705 ;
        RECT 92.185 144.615 95.295 145.525 ;
        RECT 95.305 144.715 100.815 145.525 ;
        RECT 100.825 144.715 102.655 145.525 ;
        RECT 102.665 144.845 105.415 145.525 ;
        RECT 104.485 144.615 105.415 144.845 ;
        RECT 105.425 144.715 110.935 145.525 ;
        RECT 110.945 144.715 113.695 145.525 ;
        RECT 114.175 144.655 114.605 145.440 ;
        RECT 115.545 144.745 116.915 145.525 ;
        RECT 116.925 144.715 122.435 145.525 ;
        RECT 122.445 144.715 127.955 145.525 ;
        RECT 127.965 144.715 133.475 145.525 ;
        RECT 133.485 144.715 138.995 145.525 ;
        RECT 139.935 144.655 140.365 145.440 ;
        RECT 140.385 144.715 145.895 145.525 ;
        RECT 145.905 144.715 148.655 145.525 ;
        RECT 149.125 144.715 150.495 145.525 ;
      LAYER nwell ;
        RECT 10.930 141.495 150.690 144.325 ;
      LAYER pwell ;
        RECT 11.125 140.295 12.495 141.105 ;
        RECT 12.505 140.295 16.175 141.105 ;
        RECT 16.185 140.295 17.555 141.105 ;
        RECT 17.565 140.295 18.935 141.075 ;
        RECT 18.945 140.295 22.615 141.105 ;
        RECT 22.625 140.295 23.995 141.105 ;
        RECT 24.015 140.380 24.445 141.165 ;
        RECT 24.465 140.295 28.135 141.105 ;
        RECT 28.165 140.295 29.515 141.205 ;
        RECT 29.525 140.295 35.035 141.105 ;
        RECT 35.505 140.295 38.715 141.205 ;
        RECT 38.725 140.295 42.395 141.105 ;
        RECT 44.225 140.975 45.155 141.205 ;
        RECT 42.405 140.295 45.155 140.975 ;
        RECT 45.165 140.975 46.095 141.205 ;
        RECT 45.165 140.295 47.915 140.975 ;
        RECT 47.925 140.295 49.755 141.105 ;
        RECT 49.775 140.380 50.205 141.165 ;
        RECT 50.225 140.295 52.055 141.105 ;
        RECT 52.065 140.295 54.805 140.975 ;
        RECT 54.825 140.295 60.335 141.105 ;
        RECT 60.345 140.295 64.015 141.105 ;
        RECT 64.025 140.295 65.395 141.105 ;
        RECT 65.405 140.295 66.775 141.075 ;
        RECT 66.785 140.295 72.295 141.105 ;
        RECT 72.305 140.295 75.055 141.105 ;
        RECT 75.535 140.380 75.965 141.165 ;
        RECT 76.445 140.295 77.795 141.205 ;
        RECT 77.825 140.295 83.335 141.105 ;
        RECT 83.345 140.295 88.855 141.105 ;
        RECT 88.865 140.295 94.375 141.105 ;
        RECT 94.385 140.295 99.895 141.105 ;
        RECT 99.905 140.295 101.275 141.105 ;
        RECT 101.295 140.380 101.725 141.165 ;
        RECT 101.745 140.295 104.495 141.205 ;
        RECT 104.985 140.295 106.335 141.205 ;
        RECT 106.845 140.295 110.015 141.205 ;
        RECT 110.945 140.295 114.155 141.205 ;
        RECT 114.205 140.975 115.555 141.205 ;
        RECT 117.090 140.975 118.000 141.195 ;
        RECT 114.205 140.295 121.515 140.975 ;
        RECT 121.525 140.295 127.035 141.105 ;
        RECT 127.055 140.380 127.485 141.165 ;
        RECT 127.505 140.295 133.015 141.105 ;
        RECT 133.025 140.295 138.535 141.105 ;
        RECT 138.545 140.295 144.055 141.105 ;
        RECT 144.065 140.295 147.735 141.105 ;
        RECT 147.745 140.295 149.115 141.105 ;
        RECT 149.125 140.295 150.495 141.105 ;
        RECT 11.265 140.085 11.435 140.295 ;
        RECT 12.645 140.085 12.815 140.295 ;
        RECT 15.400 140.135 15.520 140.245 ;
        RECT 15.865 140.085 16.035 140.275 ;
        RECT 16.325 140.105 16.495 140.295 ;
        RECT 18.625 140.105 18.795 140.295 ;
        RECT 19.085 140.105 19.255 140.295 ;
        RECT 22.765 140.105 22.935 140.295 ;
        RECT 23.225 140.085 23.395 140.275 ;
        RECT 24.605 140.105 24.775 140.295 ;
        RECT 26.440 140.135 26.560 140.245 ;
        RECT 26.900 140.085 27.070 140.275 ;
        RECT 28.280 140.105 28.450 140.295 ;
        RECT 29.665 140.105 29.835 140.295 ;
        RECT 32.885 140.085 33.055 140.275 ;
        RECT 33.345 140.085 33.515 140.275 ;
        RECT 35.180 140.135 35.300 140.245 ;
        RECT 35.645 140.105 35.815 140.295 ;
        RECT 38.865 140.105 39.035 140.295 ;
        RECT 42.545 140.105 42.715 140.295 ;
        RECT 46.225 140.085 46.395 140.275 ;
        RECT 46.695 140.130 46.855 140.240 ;
        RECT 47.605 140.085 47.775 140.295 ;
        RECT 48.065 140.105 48.235 140.295 ;
        RECT 50.365 140.105 50.535 140.295 ;
        RECT 52.205 140.105 52.375 140.295 ;
        RECT 54.965 140.105 55.135 140.295 ;
        RECT 56.805 140.085 56.975 140.275 ;
        RECT 11.125 139.275 12.495 140.085 ;
        RECT 12.505 139.275 15.255 140.085 ;
        RECT 15.725 139.405 23.035 140.085 ;
        RECT 19.240 139.185 20.150 139.405 ;
        RECT 21.685 139.175 23.035 139.405 ;
        RECT 23.185 139.175 26.295 140.085 ;
        RECT 26.775 139.175 29.975 140.085 ;
        RECT 29.985 139.175 33.195 140.085 ;
        RECT 33.205 139.275 36.875 140.085 ;
        RECT 36.895 139.215 37.325 140.000 ;
        RECT 37.430 139.405 46.535 140.085 ;
        RECT 47.465 139.405 56.570 140.085 ;
        RECT 56.675 139.175 59.405 140.085 ;
        RECT 59.560 140.055 59.730 140.275 ;
        RECT 60.485 140.105 60.655 140.295 ;
        RECT 61.875 140.130 62.035 140.240 ;
        RECT 63.245 140.085 63.415 140.275 ;
        RECT 64.165 140.105 64.335 140.295 ;
        RECT 65.085 140.085 65.255 140.275 ;
        RECT 66.465 140.105 66.635 140.295 ;
        RECT 66.925 140.105 67.095 140.295 ;
        RECT 67.845 140.085 68.015 140.275 ;
        RECT 71.525 140.085 71.695 140.275 ;
        RECT 72.445 140.105 72.615 140.295 ;
        RECT 72.905 140.085 73.075 140.275 ;
        RECT 75.200 140.135 75.320 140.245 ;
        RECT 76.120 140.135 76.240 140.245 ;
        RECT 77.510 140.105 77.680 140.295 ;
        RECT 77.965 140.105 78.135 140.295 ;
        RECT 78.420 140.135 78.540 140.245 ;
        RECT 77.965 140.085 78.130 140.105 ;
        RECT 78.890 140.085 79.060 140.275 ;
        RECT 82.565 140.085 82.735 140.275 ;
        RECT 83.485 140.105 83.655 140.295 ;
        RECT 89.005 140.275 89.175 140.295 ;
        RECT 84.405 140.105 84.575 140.275 ;
        RECT 84.425 140.085 84.575 140.105 ;
        RECT 87.620 140.085 87.790 140.275 ;
        RECT 88.080 140.135 88.200 140.245 ;
        RECT 89.005 140.105 89.180 140.275 ;
        RECT 89.010 140.085 89.180 140.105 ;
        RECT 90.385 140.085 90.555 140.275 ;
        RECT 94.525 140.105 94.695 140.295 ;
        RECT 98.665 140.085 98.835 140.275 ;
        RECT 99.125 140.085 99.295 140.275 ;
        RECT 100.045 140.105 100.215 140.295 ;
        RECT 100.510 140.085 100.680 140.275 ;
        RECT 101.885 140.105 102.055 140.295 ;
        RECT 103.725 140.085 103.895 140.275 ;
        RECT 104.640 140.135 104.760 140.245 ;
        RECT 106.020 140.105 106.190 140.295 ;
        RECT 106.485 140.245 106.655 140.275 ;
        RECT 106.480 140.135 106.655 140.245 ;
        RECT 106.485 140.085 106.655 140.135 ;
        RECT 106.945 140.105 107.115 140.295 ;
        RECT 108.325 140.085 108.495 140.275 ;
        RECT 110.175 140.140 110.335 140.250 ;
        RECT 111.085 140.105 111.255 140.295 ;
        RECT 113.840 140.135 113.960 140.245 ;
        RECT 114.765 140.105 114.935 140.275 ;
        RECT 114.785 140.085 114.935 140.105 ;
        RECT 117.065 140.085 117.235 140.275 ;
        RECT 121.205 140.105 121.375 140.295 ;
        RECT 121.665 140.105 121.835 140.295 ;
        RECT 122.585 140.085 122.755 140.275 ;
        RECT 127.645 140.105 127.815 140.295 ;
        RECT 128.105 140.085 128.275 140.275 ;
        RECT 133.165 140.105 133.335 140.295 ;
        RECT 133.625 140.085 133.795 140.275 ;
        RECT 138.685 140.105 138.855 140.295 ;
        RECT 139.155 140.130 139.315 140.240 ;
        RECT 140.525 140.085 140.695 140.275 ;
        RECT 144.205 140.105 144.375 140.295 ;
        RECT 146.045 140.085 146.215 140.275 ;
        RECT 147.885 140.105 148.055 140.295 ;
        RECT 148.800 140.135 148.920 140.245 ;
        RECT 150.185 140.085 150.355 140.295 ;
        RECT 60.760 140.055 61.715 140.085 ;
        RECT 59.435 139.375 61.715 140.055 ;
        RECT 60.760 139.175 61.715 139.375 ;
        RECT 62.655 139.215 63.085 140.000 ;
        RECT 63.105 139.275 64.935 140.085 ;
        RECT 64.945 139.405 67.685 140.085 ;
        RECT 67.705 139.275 71.375 140.085 ;
        RECT 71.385 139.275 72.755 140.085 ;
        RECT 72.865 139.175 75.975 140.085 ;
        RECT 76.295 139.405 78.130 140.085 ;
        RECT 76.295 139.175 77.225 139.405 ;
        RECT 78.745 139.175 82.415 140.085 ;
        RECT 82.425 139.275 84.255 140.085 ;
        RECT 84.425 139.265 86.355 140.085 ;
        RECT 85.405 139.175 86.355 139.265 ;
        RECT 86.585 139.175 87.935 140.085 ;
        RECT 88.415 139.215 88.845 140.000 ;
        RECT 88.865 139.175 90.215 140.085 ;
        RECT 90.245 139.275 91.615 140.085 ;
        RECT 91.665 139.405 98.975 140.085 ;
        RECT 91.665 139.175 93.015 139.405 ;
        RECT 94.550 139.185 95.460 139.405 ;
        RECT 98.985 139.275 100.355 140.085 ;
        RECT 100.365 139.175 103.285 140.085 ;
        RECT 103.585 139.405 106.335 140.085 ;
        RECT 105.405 139.175 106.335 139.405 ;
        RECT 106.360 139.175 108.175 140.085 ;
        RECT 108.185 139.275 113.695 140.085 ;
        RECT 114.175 139.215 114.605 140.000 ;
        RECT 114.785 139.265 116.715 140.085 ;
        RECT 116.925 139.275 122.435 140.085 ;
        RECT 122.445 139.275 127.955 140.085 ;
        RECT 127.965 139.275 133.475 140.085 ;
        RECT 133.485 139.275 138.995 140.085 ;
        RECT 115.765 139.175 116.715 139.265 ;
        RECT 139.935 139.215 140.365 140.000 ;
        RECT 140.385 139.275 145.895 140.085 ;
        RECT 145.905 139.275 148.655 140.085 ;
        RECT 149.125 139.275 150.495 140.085 ;
      LAYER nwell ;
        RECT 10.930 136.055 150.690 138.885 ;
      LAYER pwell ;
        RECT 18.685 135.675 19.635 135.765 ;
        RECT 11.125 134.855 12.495 135.665 ;
        RECT 12.505 134.855 18.015 135.665 ;
        RECT 18.685 134.855 20.615 135.675 ;
        RECT 20.785 134.855 23.535 135.665 ;
        RECT 24.015 134.940 24.445 135.725 ;
        RECT 24.465 134.855 26.295 135.665 ;
        RECT 26.405 134.855 29.515 135.765 ;
        RECT 29.525 134.855 35.035 135.665 ;
        RECT 35.045 134.855 36.875 135.665 ;
        RECT 37.345 134.855 40.515 135.765 ;
        RECT 41.495 134.855 44.225 135.765 ;
        RECT 46.965 135.565 47.915 135.765 ;
        RECT 44.245 134.885 47.915 135.565 ;
        RECT 11.265 134.645 11.435 134.855 ;
        RECT 12.645 134.645 12.815 134.855 ;
        RECT 20.465 134.835 20.615 134.855 ;
        RECT 18.165 134.805 18.335 134.835 ;
        RECT 18.160 134.695 18.335 134.805 ;
        RECT 18.165 134.645 18.335 134.695 ;
        RECT 20.465 134.665 20.635 134.835 ;
        RECT 20.925 134.665 21.095 134.855 ;
        RECT 23.685 134.805 23.855 134.835 ;
        RECT 23.680 134.695 23.855 134.805 ;
        RECT 23.685 134.645 23.855 134.695 ;
        RECT 24.605 134.665 24.775 134.855 ;
        RECT 26.445 134.665 26.615 134.855 ;
        RECT 29.205 134.645 29.375 134.835 ;
        RECT 29.665 134.665 29.835 134.855 ;
        RECT 31.040 134.695 31.160 134.805 ;
        RECT 32.425 134.645 32.595 134.835 ;
        RECT 32.885 134.645 33.055 134.835 ;
        RECT 35.185 134.665 35.355 134.855 ;
        RECT 36.570 134.645 36.740 134.835 ;
        RECT 37.020 134.695 37.140 134.805 ;
        RECT 37.490 134.645 37.660 134.835 ;
        RECT 40.245 134.665 40.415 134.855 ;
        RECT 40.715 134.700 40.875 134.810 ;
        RECT 41.160 134.695 41.280 134.805 ;
        RECT 42.540 134.645 42.710 134.835 ;
        RECT 43.925 134.665 44.095 134.855 ;
        RECT 44.390 134.665 44.560 134.885 ;
        RECT 46.965 134.855 47.915 134.885 ;
        RECT 47.925 134.855 49.275 135.765 ;
        RECT 49.775 134.940 50.205 135.725 ;
        RECT 50.725 134.855 53.895 135.765 ;
        RECT 53.905 134.855 56.655 135.665 ;
        RECT 57.145 134.855 58.495 135.765 ;
        RECT 58.505 135.565 59.450 135.765 ;
        RECT 58.505 134.885 61.255 135.565 ;
        RECT 61.265 135.535 62.185 135.765 ;
        RECT 68.000 135.535 68.910 135.755 ;
        RECT 70.445 135.535 72.215 135.765 ;
        RECT 58.505 134.855 59.450 134.885 ;
        RECT 45.765 134.645 45.935 134.835 ;
        RECT 48.070 134.665 48.240 134.855 ;
        RECT 48.525 134.645 48.695 134.835 ;
        RECT 48.985 134.645 49.155 134.835 ;
        RECT 49.440 134.695 49.560 134.805 ;
        RECT 50.360 134.695 50.480 134.805 ;
        RECT 50.825 134.665 50.995 134.855 ;
        RECT 51.740 134.695 51.860 134.805 ;
        RECT 11.125 133.835 12.495 134.645 ;
        RECT 12.505 133.835 18.015 134.645 ;
        RECT 18.025 133.835 23.535 134.645 ;
        RECT 23.545 133.835 29.055 134.645 ;
        RECT 29.065 133.835 30.895 134.645 ;
        RECT 31.375 133.735 32.725 134.645 ;
        RECT 32.745 133.835 35.495 134.645 ;
        RECT 35.505 133.735 36.855 134.645 ;
        RECT 36.895 133.775 37.325 134.560 ;
        RECT 37.345 133.735 40.820 134.645 ;
        RECT 41.505 133.735 42.855 134.645 ;
        RECT 42.865 133.735 46.035 134.645 ;
        RECT 46.095 133.735 48.825 134.645 ;
        RECT 48.845 133.835 51.595 134.645 ;
        RECT 52.210 134.615 52.380 134.835 ;
        RECT 54.045 134.665 54.215 134.855 ;
        RECT 54.965 134.645 55.135 134.835 ;
        RECT 56.800 134.695 56.920 134.805 ;
        RECT 57.260 134.665 57.430 134.855 ;
        RECT 60.485 134.645 60.655 134.835 ;
        RECT 60.940 134.665 61.110 134.885 ;
        RECT 61.265 134.855 63.555 135.535 ;
        RECT 64.485 134.855 72.215 135.535 ;
        RECT 72.305 135.535 73.225 135.765 ;
        RECT 72.305 134.855 74.595 135.535 ;
        RECT 75.535 134.940 75.965 135.725 ;
        RECT 75.985 135.535 76.905 135.765 ;
        RECT 75.985 134.855 78.275 135.535 ;
        RECT 78.285 134.855 81.955 135.665 ;
        RECT 81.965 134.855 83.780 135.765 ;
        RECT 83.805 134.855 85.155 135.765 ;
        RECT 85.185 134.855 87.015 135.665 ;
        RECT 87.525 134.855 90.695 135.765 ;
        RECT 90.705 134.855 92.075 135.665 ;
        RECT 92.085 134.855 95.295 135.765 ;
        RECT 96.445 135.675 97.395 135.765 ;
        RECT 95.465 134.855 97.395 135.675 ;
        RECT 97.605 134.855 98.975 135.635 ;
        RECT 98.985 134.855 100.815 135.665 ;
        RECT 101.295 134.940 101.725 135.725 ;
        RECT 101.745 134.855 107.255 135.665 ;
        RECT 107.265 134.855 112.775 135.665 ;
        RECT 112.785 134.855 118.295 135.665 ;
        RECT 118.305 134.855 123.815 135.665 ;
        RECT 123.825 134.855 126.575 135.665 ;
        RECT 127.055 134.940 127.485 135.725 ;
        RECT 127.505 134.855 133.015 135.665 ;
        RECT 133.025 134.855 138.535 135.665 ;
        RECT 138.545 134.855 144.055 135.665 ;
        RECT 144.065 134.855 147.735 135.665 ;
        RECT 147.745 134.855 149.115 135.665 ;
        RECT 149.125 134.855 150.495 135.665 ;
        RECT 62.320 134.695 62.440 134.805 ;
        RECT 63.245 134.645 63.415 134.855 ;
        RECT 63.715 134.700 63.875 134.810 ;
        RECT 64.625 134.665 64.795 134.855 ;
        RECT 65.080 134.695 65.200 134.805 ;
        RECT 66.470 134.645 66.640 134.835 ;
        RECT 66.935 134.690 67.095 134.800 ;
        RECT 67.845 134.645 68.015 134.835 ;
        RECT 70.605 134.645 70.775 134.835 ;
        RECT 74.285 134.665 74.455 134.855 ;
        RECT 74.755 134.700 74.915 134.810 ;
        RECT 76.125 134.645 76.295 134.835 ;
        RECT 77.965 134.665 78.135 134.855 ;
        RECT 78.425 134.665 78.595 134.855 ;
        RECT 81.645 134.645 81.815 134.835 ;
        RECT 83.485 134.665 83.655 134.855 ;
        RECT 84.870 134.665 85.040 134.855 ;
        RECT 85.325 134.665 85.495 134.855 ;
        RECT 87.165 134.805 87.335 134.835 ;
        RECT 87.160 134.695 87.335 134.805 ;
        RECT 87.165 134.645 87.335 134.695 ;
        RECT 87.625 134.665 87.795 134.855 ;
        RECT 89.005 134.645 89.175 134.835 ;
        RECT 90.845 134.665 91.015 134.855 ;
        RECT 92.225 134.665 92.395 134.855 ;
        RECT 95.465 134.835 95.615 134.855 ;
        RECT 94.525 134.645 94.695 134.835 ;
        RECT 95.445 134.665 95.615 134.835 ;
        RECT 98.665 134.665 98.835 134.855 ;
        RECT 99.125 134.665 99.295 134.855 ;
        RECT 100.045 134.645 100.215 134.835 ;
        RECT 100.960 134.695 101.080 134.805 ;
        RECT 101.425 134.645 101.595 134.835 ;
        RECT 101.885 134.665 102.055 134.855 ;
        RECT 104.645 134.645 104.815 134.835 ;
        RECT 106.020 134.695 106.140 134.805 ;
        RECT 106.485 134.645 106.655 134.835 ;
        RECT 107.405 134.665 107.575 134.855 ;
        RECT 109.705 134.665 109.875 134.835 ;
        RECT 109.725 134.645 109.875 134.665 ;
        RECT 112.005 134.645 112.175 134.835 ;
        RECT 112.925 134.665 113.095 134.855 ;
        RECT 113.395 134.690 113.555 134.800 ;
        RECT 114.765 134.645 114.935 134.835 ;
        RECT 118.445 134.665 118.615 134.855 ;
        RECT 120.285 134.645 120.455 134.835 ;
        RECT 123.965 134.665 124.135 134.855 ;
        RECT 125.805 134.645 125.975 134.835 ;
        RECT 126.720 134.695 126.840 134.805 ;
        RECT 127.645 134.665 127.815 134.855 ;
        RECT 131.325 134.645 131.495 134.835 ;
        RECT 133.165 134.665 133.335 134.855 ;
        RECT 136.845 134.645 137.015 134.835 ;
        RECT 138.685 134.665 138.855 134.855 ;
        RECT 139.600 134.695 139.720 134.805 ;
        RECT 140.525 134.645 140.695 134.835 ;
        RECT 144.205 134.665 144.375 134.855 ;
        RECT 146.045 134.645 146.215 134.835 ;
        RECT 147.885 134.665 148.055 134.855 ;
        RECT 148.800 134.695 148.920 134.805 ;
        RECT 150.185 134.645 150.355 134.855 ;
        RECT 53.870 134.615 54.815 134.645 ;
        RECT 52.065 133.935 54.815 134.615 ;
        RECT 53.870 133.735 54.815 133.935 ;
        RECT 54.825 133.835 60.335 134.645 ;
        RECT 60.345 133.835 62.175 134.645 ;
        RECT 62.655 133.775 63.085 134.560 ;
        RECT 63.105 133.835 64.935 134.645 ;
        RECT 65.405 133.735 66.755 134.645 ;
        RECT 67.705 133.735 70.455 134.645 ;
        RECT 70.465 133.835 75.975 134.645 ;
        RECT 75.985 133.835 81.495 134.645 ;
        RECT 81.505 133.835 87.015 134.645 ;
        RECT 87.025 133.835 88.395 134.645 ;
        RECT 88.415 133.775 88.845 134.560 ;
        RECT 88.865 133.835 94.375 134.645 ;
        RECT 94.385 133.835 99.895 134.645 ;
        RECT 99.905 133.835 101.275 134.645 ;
        RECT 101.385 133.735 104.495 134.645 ;
        RECT 104.515 133.735 105.865 134.645 ;
        RECT 106.345 133.735 109.555 134.645 ;
        RECT 109.725 133.825 111.655 134.645 ;
        RECT 111.865 133.865 113.235 134.645 ;
        RECT 110.705 133.735 111.655 133.825 ;
        RECT 114.175 133.775 114.605 134.560 ;
        RECT 114.625 133.835 120.135 134.645 ;
        RECT 120.145 133.835 125.655 134.645 ;
        RECT 125.665 133.835 131.175 134.645 ;
        RECT 131.185 133.835 136.695 134.645 ;
        RECT 136.705 133.835 139.455 134.645 ;
        RECT 139.935 133.775 140.365 134.560 ;
        RECT 140.385 133.835 145.895 134.645 ;
        RECT 145.905 133.835 148.655 134.645 ;
        RECT 149.125 133.835 150.495 134.645 ;
      LAYER nwell ;
        RECT 10.930 130.615 150.690 133.445 ;
      LAYER pwell ;
        RECT 11.125 129.415 12.495 130.225 ;
        RECT 12.505 129.415 18.015 130.225 ;
        RECT 18.025 129.415 23.535 130.225 ;
        RECT 24.015 129.500 24.445 130.285 ;
        RECT 24.465 129.415 27.215 130.225 ;
        RECT 27.265 130.095 28.615 130.325 ;
        RECT 30.150 130.095 31.060 130.315 ;
        RECT 27.265 129.415 34.575 130.095 ;
        RECT 34.585 129.415 40.095 130.225 ;
        RECT 40.105 129.415 41.935 130.225 ;
        RECT 41.945 129.415 45.155 130.325 ;
        RECT 45.165 129.415 48.835 130.225 ;
        RECT 49.775 129.500 50.205 130.285 ;
        RECT 50.225 129.415 52.055 130.225 ;
        RECT 52.540 129.415 54.355 130.325 ;
        RECT 54.365 129.415 57.285 130.325 ;
        RECT 58.505 130.125 59.435 130.325 ;
        RECT 60.770 130.125 61.715 130.325 ;
        RECT 58.505 129.645 61.715 130.125 ;
        RECT 58.645 129.445 61.715 129.645 ;
        RECT 11.265 129.205 11.435 129.415 ;
        RECT 12.645 129.205 12.815 129.415 ;
        RECT 18.165 129.205 18.335 129.415 ;
        RECT 23.685 129.365 23.855 129.395 ;
        RECT 23.680 129.255 23.855 129.365 ;
        RECT 23.685 129.205 23.855 129.255 ;
        RECT 24.605 129.225 24.775 129.415 ;
        RECT 29.205 129.205 29.375 129.395 ;
        RECT 34.265 129.225 34.435 129.415 ;
        RECT 34.725 129.205 34.895 129.415 ;
        RECT 36.560 129.255 36.680 129.365 ;
        RECT 37.485 129.205 37.655 129.395 ;
        RECT 40.245 129.225 40.415 129.415 ;
        RECT 41.175 129.250 41.335 129.360 ;
        RECT 42.085 129.225 42.255 129.415 ;
        RECT 42.090 129.205 42.255 129.225 ;
        RECT 44.385 129.205 44.555 129.395 ;
        RECT 45.305 129.225 45.475 129.415 ;
        RECT 45.765 129.205 45.935 129.395 ;
        RECT 48.520 129.255 48.640 129.365 ;
        RECT 48.995 129.260 49.155 129.370 ;
        RECT 49.900 129.205 50.070 129.395 ;
        RECT 50.365 129.365 50.535 129.415 ;
        RECT 50.360 129.255 50.535 129.365 ;
        RECT 50.365 129.225 50.535 129.255 ;
        RECT 50.830 129.205 51.000 129.395 ;
        RECT 52.200 129.255 52.320 129.365 ;
        RECT 52.665 129.225 52.835 129.415 ;
        RECT 54.510 129.395 54.680 129.415 ;
        RECT 54.505 129.225 54.680 129.395 ;
        RECT 57.735 129.260 57.895 129.370 ;
        RECT 58.195 129.250 58.355 129.360 ;
        RECT 58.645 129.225 58.815 129.445 ;
        RECT 60.770 129.415 61.715 129.445 ;
        RECT 61.725 129.415 67.235 130.225 ;
        RECT 67.555 130.095 68.485 130.325 ;
        RECT 67.555 129.415 69.390 130.095 ;
        RECT 69.545 129.415 73.215 130.225 ;
        RECT 73.700 129.415 75.515 130.325 ;
        RECT 75.535 129.500 75.965 130.285 ;
        RECT 75.985 130.095 76.910 130.325 ;
        RECT 80.715 130.095 81.645 130.325 ;
        RECT 75.985 129.415 79.655 130.095 ;
        RECT 79.810 129.415 81.645 130.095 ;
        RECT 81.965 129.415 83.335 130.225 ;
        RECT 85.420 130.095 86.555 130.325 ;
        RECT 83.345 129.415 86.555 130.095 ;
        RECT 86.565 129.415 89.775 130.325 ;
        RECT 89.785 129.415 95.295 130.225 ;
        RECT 95.305 129.415 97.135 130.225 ;
        RECT 97.645 129.415 100.815 130.325 ;
        RECT 101.295 129.500 101.725 130.285 ;
        RECT 101.745 129.415 105.415 130.225 ;
        RECT 105.425 129.415 106.795 130.225 ;
        RECT 106.885 130.095 108.655 130.325 ;
        RECT 110.190 130.095 111.100 130.315 ;
        RECT 106.885 129.415 114.615 130.095 ;
        RECT 114.625 129.415 120.135 130.225 ;
        RECT 120.145 129.415 125.655 130.225 ;
        RECT 125.665 129.415 127.035 130.225 ;
        RECT 127.055 129.500 127.485 130.285 ;
        RECT 127.505 129.415 133.015 130.225 ;
        RECT 133.025 129.415 138.535 130.225 ;
        RECT 138.545 129.415 144.055 130.225 ;
        RECT 144.065 129.415 147.735 130.225 ;
        RECT 147.745 129.415 149.115 130.225 ;
        RECT 149.125 129.415 150.495 130.225 ;
        RECT 54.505 129.205 54.675 129.225 ;
        RECT 59.105 129.205 59.275 129.395 ;
        RECT 60.940 129.205 61.110 129.395 ;
        RECT 61.865 129.225 62.035 129.415 ;
        RECT 69.225 129.395 69.390 129.415 ;
        RECT 62.320 129.255 62.440 129.365 ;
        RECT 66.465 129.205 66.635 129.395 ;
        RECT 66.925 129.205 67.095 129.395 ;
        RECT 69.225 129.225 69.395 129.395 ;
        RECT 69.685 129.225 69.855 129.415 ;
        RECT 73.360 129.255 73.480 129.365 ;
        RECT 73.825 129.225 73.995 129.415 ;
        RECT 74.285 129.205 74.455 129.395 ;
        RECT 76.130 129.225 76.300 129.415 ;
        RECT 79.810 129.395 79.975 129.415 ;
        RECT 78.425 129.205 78.595 129.395 ;
        RECT 78.885 129.205 79.055 129.395 ;
        RECT 79.805 129.225 79.975 129.395 ;
        RECT 80.720 129.255 80.840 129.365 ;
        RECT 81.180 129.205 81.350 129.395 ;
        RECT 82.105 129.225 82.275 129.415 ;
        RECT 82.565 129.225 82.735 129.395 ;
        RECT 83.485 129.225 83.655 129.415 ;
        RECT 84.860 129.255 84.980 129.365 ;
        RECT 86.705 129.225 86.875 129.415 ;
        RECT 82.570 129.205 82.735 129.225 ;
        RECT 11.125 128.395 12.495 129.205 ;
        RECT 12.505 128.395 18.015 129.205 ;
        RECT 18.025 128.395 23.535 129.205 ;
        RECT 23.545 128.395 29.055 129.205 ;
        RECT 29.065 128.395 34.575 129.205 ;
        RECT 34.585 128.395 36.415 129.205 ;
        RECT 36.895 128.335 37.325 129.120 ;
        RECT 37.345 128.395 41.015 129.205 ;
        RECT 42.090 128.525 43.925 129.205 ;
        RECT 42.995 128.295 43.925 128.525 ;
        RECT 44.245 128.425 45.615 129.205 ;
        RECT 45.625 128.395 48.375 129.205 ;
        RECT 48.865 128.295 50.215 129.205 ;
        RECT 50.685 128.525 54.355 129.205 ;
        RECT 50.685 128.295 51.610 128.525 ;
        RECT 54.365 128.395 58.035 129.205 ;
        RECT 58.980 128.295 60.795 129.205 ;
        RECT 60.825 128.295 62.175 129.205 ;
        RECT 62.655 128.335 63.085 129.120 ;
        RECT 63.200 128.525 66.665 129.205 ;
        RECT 66.785 128.525 74.095 129.205 ;
        RECT 63.200 128.295 64.120 128.525 ;
        RECT 70.300 128.305 71.210 128.525 ;
        RECT 72.745 128.295 74.095 128.525 ;
        RECT 74.145 128.395 75.515 129.205 ;
        RECT 75.525 128.295 78.635 129.205 ;
        RECT 78.745 128.395 80.575 129.205 ;
        RECT 81.065 128.295 82.415 129.205 ;
        RECT 82.570 128.525 84.405 129.205 ;
        RECT 83.475 128.295 84.405 128.525 ;
        RECT 85.185 129.175 86.130 129.205 ;
        RECT 88.085 129.175 88.255 129.395 ;
        RECT 89.925 129.225 90.095 129.415 ;
        RECT 90.385 129.205 90.555 129.395 ;
        RECT 95.445 129.225 95.615 129.415 ;
        RECT 97.280 129.255 97.400 129.365 ;
        RECT 97.745 129.225 97.915 129.415 ;
        RECT 98.205 129.205 98.375 129.395 ;
        RECT 98.665 129.205 98.835 129.395 ;
        RECT 100.960 129.255 101.080 129.365 ;
        RECT 101.885 129.225 102.055 129.415 ;
        RECT 104.185 129.205 104.355 129.395 ;
        RECT 105.565 129.225 105.735 129.415 ;
        RECT 109.705 129.205 109.875 129.395 ;
        RECT 113.395 129.250 113.555 129.360 ;
        RECT 114.305 129.225 114.475 129.415 ;
        RECT 114.765 129.205 114.935 129.415 ;
        RECT 120.285 129.205 120.455 129.415 ;
        RECT 125.805 129.205 125.975 129.415 ;
        RECT 127.645 129.225 127.815 129.415 ;
        RECT 131.325 129.205 131.495 129.395 ;
        RECT 133.165 129.225 133.335 129.415 ;
        RECT 136.845 129.205 137.015 129.395 ;
        RECT 138.685 129.225 138.855 129.415 ;
        RECT 139.600 129.255 139.720 129.365 ;
        RECT 140.525 129.205 140.695 129.395 ;
        RECT 144.205 129.225 144.375 129.415 ;
        RECT 146.045 129.205 146.215 129.395 ;
        RECT 147.885 129.225 148.055 129.415 ;
        RECT 148.800 129.255 148.920 129.365 ;
        RECT 150.185 129.205 150.355 129.415 ;
        RECT 85.185 128.975 88.255 129.175 ;
        RECT 85.185 128.495 88.395 128.975 ;
        RECT 85.185 128.295 86.130 128.495 ;
        RECT 87.465 128.295 88.395 128.495 ;
        RECT 88.415 128.335 88.845 129.120 ;
        RECT 88.865 128.295 90.680 129.205 ;
        RECT 90.785 128.525 98.515 129.205 ;
        RECT 90.785 128.295 92.555 128.525 ;
        RECT 94.090 128.305 95.000 128.525 ;
        RECT 98.525 128.395 104.035 129.205 ;
        RECT 104.045 128.395 109.555 129.205 ;
        RECT 109.565 128.395 113.235 129.205 ;
        RECT 114.175 128.335 114.605 129.120 ;
        RECT 114.625 128.395 120.135 129.205 ;
        RECT 120.145 128.395 125.655 129.205 ;
        RECT 125.665 128.395 131.175 129.205 ;
        RECT 131.185 128.395 136.695 129.205 ;
        RECT 136.705 128.395 139.455 129.205 ;
        RECT 139.935 128.335 140.365 129.120 ;
        RECT 140.385 128.395 145.895 129.205 ;
        RECT 145.905 128.395 148.655 129.205 ;
        RECT 149.125 128.395 150.495 129.205 ;
      LAYER nwell ;
        RECT 10.930 125.175 150.690 128.005 ;
      LAYER pwell ;
        RECT 11.125 123.975 12.495 124.785 ;
        RECT 12.505 123.975 18.015 124.785 ;
        RECT 18.025 123.975 23.535 124.785 ;
        RECT 24.015 124.060 24.445 124.845 ;
        RECT 24.465 123.975 29.975 124.785 ;
        RECT 29.985 123.975 35.495 124.785 ;
        RECT 35.505 123.975 39.175 124.785 ;
        RECT 39.265 124.655 41.035 124.885 ;
        RECT 42.570 124.655 43.480 124.875 ;
        RECT 39.265 123.975 46.995 124.655 ;
        RECT 47.005 123.975 49.755 124.785 ;
        RECT 49.775 124.060 50.205 124.845 ;
        RECT 50.225 123.975 55.735 124.785 ;
        RECT 55.745 123.975 57.575 124.785 ;
        RECT 61.100 124.655 62.010 124.875 ;
        RECT 63.545 124.655 65.315 124.885 ;
        RECT 57.585 123.975 65.315 124.655 ;
        RECT 65.405 123.975 66.775 124.755 ;
        RECT 66.785 123.975 72.295 124.785 ;
        RECT 72.305 123.975 75.055 124.785 ;
        RECT 75.535 124.060 75.965 124.845 ;
        RECT 75.985 123.975 81.495 124.785 ;
        RECT 81.505 123.975 87.015 124.785 ;
        RECT 87.025 123.975 90.695 124.785 ;
        RECT 94.280 124.655 95.200 124.885 ;
        RECT 91.735 123.975 95.200 124.655 ;
        RECT 95.305 123.975 96.655 124.885 ;
        RECT 96.685 123.975 100.355 124.785 ;
        RECT 101.295 124.060 101.725 124.845 ;
        RECT 101.745 123.975 107.255 124.785 ;
        RECT 107.265 123.975 112.775 124.785 ;
        RECT 112.785 123.975 118.295 124.785 ;
        RECT 118.305 123.975 123.815 124.785 ;
        RECT 123.825 123.975 126.575 124.785 ;
        RECT 127.055 124.060 127.485 124.845 ;
        RECT 127.505 123.975 133.015 124.785 ;
        RECT 133.025 123.975 138.535 124.785 ;
        RECT 138.545 123.975 144.055 124.785 ;
        RECT 144.065 123.975 147.735 124.785 ;
        RECT 147.745 123.975 149.115 124.785 ;
        RECT 149.125 123.975 150.495 124.785 ;
        RECT 11.265 123.765 11.435 123.975 ;
        RECT 12.645 123.765 12.815 123.975 ;
        RECT 18.165 123.765 18.335 123.975 ;
        RECT 23.685 123.925 23.855 123.955 ;
        RECT 23.680 123.815 23.855 123.925 ;
        RECT 23.685 123.765 23.855 123.815 ;
        RECT 24.605 123.785 24.775 123.975 ;
        RECT 29.205 123.765 29.375 123.955 ;
        RECT 30.125 123.785 30.295 123.975 ;
        RECT 34.725 123.765 34.895 123.955 ;
        RECT 35.645 123.785 35.815 123.975 ;
        RECT 36.560 123.815 36.680 123.925 ;
        RECT 37.485 123.765 37.655 123.955 ;
        RECT 43.005 123.765 43.175 123.955 ;
        RECT 46.685 123.785 46.855 123.975 ;
        RECT 47.145 123.785 47.315 123.975 ;
        RECT 47.605 123.765 47.775 123.955 ;
        RECT 50.365 123.785 50.535 123.975 ;
        RECT 55.425 123.765 55.595 123.955 ;
        RECT 55.885 123.785 56.055 123.975 ;
        RECT 57.725 123.785 57.895 123.975 ;
        RECT 60.945 123.765 61.115 123.955 ;
        RECT 63.245 123.765 63.415 123.955 ;
        RECT 65.545 123.785 65.715 123.975 ;
        RECT 66.925 123.785 67.095 123.975 ;
        RECT 68.765 123.765 68.935 123.955 ;
        RECT 72.445 123.785 72.615 123.975 ;
        RECT 74.285 123.765 74.455 123.955 ;
        RECT 75.200 123.815 75.320 123.925 ;
        RECT 76.125 123.785 76.295 123.975 ;
        RECT 79.805 123.765 79.975 123.955 ;
        RECT 81.645 123.785 81.815 123.975 ;
        RECT 85.325 123.765 85.495 123.955 ;
        RECT 87.165 123.785 87.335 123.975 ;
        RECT 88.080 123.815 88.200 123.925 ;
        RECT 89.005 123.765 89.175 123.955 ;
        RECT 90.855 123.820 91.015 123.930 ;
        RECT 91.765 123.785 91.935 123.975 ;
        RECT 94.525 123.765 94.695 123.955 ;
        RECT 96.370 123.785 96.540 123.975 ;
        RECT 96.825 123.785 96.995 123.975 ;
        RECT 100.045 123.765 100.215 123.955 ;
        RECT 100.515 123.820 100.675 123.930 ;
        RECT 101.885 123.785 102.055 123.975 ;
        RECT 105.565 123.765 105.735 123.955 ;
        RECT 107.405 123.785 107.575 123.975 ;
        RECT 111.085 123.765 111.255 123.955 ;
        RECT 112.925 123.785 113.095 123.975 ;
        RECT 113.840 123.815 113.960 123.925 ;
        RECT 114.765 123.765 114.935 123.955 ;
        RECT 118.445 123.785 118.615 123.975 ;
        RECT 120.285 123.765 120.455 123.955 ;
        RECT 123.965 123.785 124.135 123.975 ;
        RECT 125.805 123.765 125.975 123.955 ;
        RECT 126.720 123.815 126.840 123.925 ;
        RECT 127.645 123.785 127.815 123.975 ;
        RECT 131.325 123.765 131.495 123.955 ;
        RECT 133.165 123.785 133.335 123.975 ;
        RECT 136.845 123.765 137.015 123.955 ;
        RECT 138.685 123.785 138.855 123.975 ;
        RECT 139.600 123.815 139.720 123.925 ;
        RECT 140.525 123.765 140.695 123.955 ;
        RECT 144.205 123.785 144.375 123.975 ;
        RECT 146.045 123.765 146.215 123.955 ;
        RECT 147.885 123.785 148.055 123.975 ;
        RECT 148.800 123.815 148.920 123.925 ;
        RECT 150.185 123.765 150.355 123.975 ;
        RECT 11.125 122.955 12.495 123.765 ;
        RECT 12.505 122.955 18.015 123.765 ;
        RECT 18.025 122.955 23.535 123.765 ;
        RECT 23.545 122.955 29.055 123.765 ;
        RECT 29.065 122.955 34.575 123.765 ;
        RECT 34.585 122.955 36.415 123.765 ;
        RECT 36.895 122.895 37.325 123.680 ;
        RECT 37.345 122.955 42.855 123.765 ;
        RECT 42.865 122.955 46.535 123.765 ;
        RECT 47.465 123.085 55.195 123.765 ;
        RECT 50.980 122.865 51.890 123.085 ;
        RECT 53.425 122.855 55.195 123.085 ;
        RECT 55.285 122.955 60.795 123.765 ;
        RECT 60.805 122.955 62.635 123.765 ;
        RECT 62.655 122.895 63.085 123.680 ;
        RECT 63.105 122.955 68.615 123.765 ;
        RECT 68.625 122.955 74.135 123.765 ;
        RECT 74.145 122.955 79.655 123.765 ;
        RECT 79.665 122.955 85.175 123.765 ;
        RECT 85.185 122.955 87.935 123.765 ;
        RECT 88.415 122.895 88.845 123.680 ;
        RECT 88.865 122.955 94.375 123.765 ;
        RECT 94.385 122.955 99.895 123.765 ;
        RECT 99.905 122.955 105.415 123.765 ;
        RECT 105.425 122.955 110.935 123.765 ;
        RECT 110.945 122.955 113.695 123.765 ;
        RECT 114.175 122.895 114.605 123.680 ;
        RECT 114.625 122.955 120.135 123.765 ;
        RECT 120.145 122.955 125.655 123.765 ;
        RECT 125.665 122.955 131.175 123.765 ;
        RECT 131.185 122.955 136.695 123.765 ;
        RECT 136.705 122.955 139.455 123.765 ;
        RECT 139.935 122.895 140.365 123.680 ;
        RECT 140.385 122.955 145.895 123.765 ;
        RECT 145.905 122.955 148.655 123.765 ;
        RECT 149.125 122.955 150.495 123.765 ;
      LAYER nwell ;
        RECT 10.930 119.735 150.690 122.565 ;
      LAYER pwell ;
        RECT 11.125 118.535 12.495 119.345 ;
        RECT 12.505 118.535 18.015 119.345 ;
        RECT 18.025 118.535 23.535 119.345 ;
        RECT 24.015 118.620 24.445 119.405 ;
        RECT 24.465 118.535 29.975 119.345 ;
        RECT 29.985 118.535 35.495 119.345 ;
        RECT 35.505 118.535 41.015 119.345 ;
        RECT 41.025 118.535 46.535 119.345 ;
        RECT 46.545 118.535 49.295 119.345 ;
        RECT 49.775 118.620 50.205 119.405 ;
        RECT 50.225 118.535 55.735 119.345 ;
        RECT 55.745 118.535 61.255 119.345 ;
        RECT 61.265 118.535 66.775 119.345 ;
        RECT 66.785 118.535 72.295 119.345 ;
        RECT 72.305 118.535 75.055 119.345 ;
        RECT 75.535 118.620 75.965 119.405 ;
        RECT 75.985 118.535 81.495 119.345 ;
        RECT 81.505 118.535 87.015 119.345 ;
        RECT 87.025 118.535 92.535 119.345 ;
        RECT 92.545 118.535 98.055 119.345 ;
        RECT 98.065 118.535 100.815 119.345 ;
        RECT 101.295 118.620 101.725 119.405 ;
        RECT 101.745 118.535 107.255 119.345 ;
        RECT 107.265 118.535 112.775 119.345 ;
        RECT 112.785 118.535 118.295 119.345 ;
        RECT 118.305 118.535 123.815 119.345 ;
        RECT 123.825 118.535 126.575 119.345 ;
        RECT 127.055 118.620 127.485 119.405 ;
        RECT 127.505 118.535 133.015 119.345 ;
        RECT 133.025 118.535 138.535 119.345 ;
        RECT 138.545 118.535 144.055 119.345 ;
        RECT 144.065 118.535 147.735 119.345 ;
        RECT 147.745 118.535 149.115 119.345 ;
        RECT 149.125 118.535 150.495 119.345 ;
        RECT 11.265 118.325 11.435 118.535 ;
        RECT 12.645 118.325 12.815 118.535 ;
        RECT 18.165 118.325 18.335 118.535 ;
        RECT 23.685 118.485 23.855 118.515 ;
        RECT 23.680 118.375 23.855 118.485 ;
        RECT 23.685 118.325 23.855 118.375 ;
        RECT 24.605 118.345 24.775 118.535 ;
        RECT 29.205 118.325 29.375 118.515 ;
        RECT 30.125 118.345 30.295 118.535 ;
        RECT 34.725 118.325 34.895 118.515 ;
        RECT 35.645 118.345 35.815 118.535 ;
        RECT 36.560 118.375 36.680 118.485 ;
        RECT 37.485 118.325 37.655 118.515 ;
        RECT 41.165 118.345 41.335 118.535 ;
        RECT 43.005 118.325 43.175 118.515 ;
        RECT 46.685 118.345 46.855 118.535 ;
        RECT 48.525 118.325 48.695 118.515 ;
        RECT 49.440 118.375 49.560 118.485 ;
        RECT 50.365 118.345 50.535 118.535 ;
        RECT 54.045 118.325 54.215 118.515 ;
        RECT 55.885 118.345 56.055 118.535 ;
        RECT 59.565 118.325 59.735 118.515 ;
        RECT 61.405 118.345 61.575 118.535 ;
        RECT 62.320 118.375 62.440 118.485 ;
        RECT 63.245 118.325 63.415 118.515 ;
        RECT 66.925 118.345 67.095 118.535 ;
        RECT 68.765 118.325 68.935 118.515 ;
        RECT 72.445 118.345 72.615 118.535 ;
        RECT 74.285 118.325 74.455 118.515 ;
        RECT 75.200 118.375 75.320 118.485 ;
        RECT 76.125 118.345 76.295 118.535 ;
        RECT 79.805 118.325 79.975 118.515 ;
        RECT 81.645 118.345 81.815 118.535 ;
        RECT 85.325 118.325 85.495 118.515 ;
        RECT 87.165 118.345 87.335 118.535 ;
        RECT 88.080 118.375 88.200 118.485 ;
        RECT 89.005 118.325 89.175 118.515 ;
        RECT 92.685 118.345 92.855 118.535 ;
        RECT 94.525 118.325 94.695 118.515 ;
        RECT 98.205 118.345 98.375 118.535 ;
        RECT 100.045 118.325 100.215 118.515 ;
        RECT 100.960 118.375 101.080 118.485 ;
        RECT 101.885 118.345 102.055 118.535 ;
        RECT 105.565 118.325 105.735 118.515 ;
        RECT 107.405 118.345 107.575 118.535 ;
        RECT 111.085 118.325 111.255 118.515 ;
        RECT 112.925 118.345 113.095 118.535 ;
        RECT 113.840 118.375 113.960 118.485 ;
        RECT 114.765 118.325 114.935 118.515 ;
        RECT 118.445 118.345 118.615 118.535 ;
        RECT 120.285 118.325 120.455 118.515 ;
        RECT 123.965 118.345 124.135 118.535 ;
        RECT 125.805 118.325 125.975 118.515 ;
        RECT 126.720 118.375 126.840 118.485 ;
        RECT 127.645 118.345 127.815 118.535 ;
        RECT 131.325 118.325 131.495 118.515 ;
        RECT 133.165 118.345 133.335 118.535 ;
        RECT 136.845 118.325 137.015 118.515 ;
        RECT 138.685 118.345 138.855 118.535 ;
        RECT 139.600 118.375 139.720 118.485 ;
        RECT 140.525 118.325 140.695 118.515 ;
        RECT 144.205 118.345 144.375 118.535 ;
        RECT 146.045 118.325 146.215 118.515 ;
        RECT 147.885 118.345 148.055 118.535 ;
        RECT 148.800 118.375 148.920 118.485 ;
        RECT 150.185 118.325 150.355 118.535 ;
        RECT 11.125 117.515 12.495 118.325 ;
        RECT 12.505 117.515 18.015 118.325 ;
        RECT 18.025 117.515 23.535 118.325 ;
        RECT 23.545 117.515 29.055 118.325 ;
        RECT 29.065 117.515 34.575 118.325 ;
        RECT 34.585 117.515 36.415 118.325 ;
        RECT 36.895 117.455 37.325 118.240 ;
        RECT 37.345 117.515 42.855 118.325 ;
        RECT 42.865 117.515 48.375 118.325 ;
        RECT 48.385 117.515 53.895 118.325 ;
        RECT 53.905 117.515 59.415 118.325 ;
        RECT 59.425 117.515 62.175 118.325 ;
        RECT 62.655 117.455 63.085 118.240 ;
        RECT 63.105 117.515 68.615 118.325 ;
        RECT 68.625 117.515 74.135 118.325 ;
        RECT 74.145 117.515 79.655 118.325 ;
        RECT 79.665 117.515 85.175 118.325 ;
        RECT 85.185 117.515 87.935 118.325 ;
        RECT 88.415 117.455 88.845 118.240 ;
        RECT 88.865 117.515 94.375 118.325 ;
        RECT 94.385 117.515 99.895 118.325 ;
        RECT 99.905 117.515 105.415 118.325 ;
        RECT 105.425 117.515 110.935 118.325 ;
        RECT 110.945 117.515 113.695 118.325 ;
        RECT 114.175 117.455 114.605 118.240 ;
        RECT 114.625 117.515 120.135 118.325 ;
        RECT 120.145 117.515 125.655 118.325 ;
        RECT 125.665 117.515 131.175 118.325 ;
        RECT 131.185 117.515 136.695 118.325 ;
        RECT 136.705 117.515 139.455 118.325 ;
        RECT 139.935 117.455 140.365 118.240 ;
        RECT 140.385 117.515 145.895 118.325 ;
        RECT 145.905 117.515 148.655 118.325 ;
        RECT 149.125 117.515 150.495 118.325 ;
      LAYER nwell ;
        RECT 10.930 114.295 150.690 117.125 ;
      LAYER pwell ;
        RECT 11.125 113.095 12.495 113.905 ;
        RECT 12.505 113.095 18.015 113.905 ;
        RECT 18.025 113.095 23.535 113.905 ;
        RECT 24.015 113.180 24.445 113.965 ;
        RECT 24.465 113.095 29.975 113.905 ;
        RECT 29.985 113.095 35.495 113.905 ;
        RECT 35.505 113.095 41.015 113.905 ;
        RECT 41.025 113.095 46.535 113.905 ;
        RECT 46.545 113.095 49.295 113.905 ;
        RECT 49.775 113.180 50.205 113.965 ;
        RECT 50.225 113.095 55.735 113.905 ;
        RECT 55.745 113.095 61.255 113.905 ;
        RECT 61.265 113.095 66.775 113.905 ;
        RECT 66.785 113.095 72.295 113.905 ;
        RECT 72.305 113.095 75.055 113.905 ;
        RECT 75.535 113.180 75.965 113.965 ;
        RECT 75.985 113.095 81.495 113.905 ;
        RECT 81.505 113.095 87.015 113.905 ;
        RECT 87.025 113.095 92.535 113.905 ;
        RECT 92.545 113.095 98.055 113.905 ;
        RECT 98.065 113.095 100.815 113.905 ;
        RECT 101.295 113.180 101.725 113.965 ;
        RECT 101.745 113.095 107.255 113.905 ;
        RECT 107.265 113.095 112.775 113.905 ;
        RECT 112.785 113.095 118.295 113.905 ;
        RECT 118.305 113.095 123.815 113.905 ;
        RECT 123.825 113.095 126.575 113.905 ;
        RECT 127.055 113.180 127.485 113.965 ;
        RECT 127.505 113.095 133.015 113.905 ;
        RECT 133.025 113.095 138.535 113.905 ;
        RECT 138.545 113.095 144.055 113.905 ;
        RECT 144.065 113.095 147.735 113.905 ;
        RECT 147.745 113.095 149.115 113.905 ;
        RECT 149.125 113.095 150.495 113.905 ;
        RECT 11.265 112.885 11.435 113.095 ;
        RECT 12.645 112.885 12.815 113.095 ;
        RECT 18.165 112.885 18.335 113.095 ;
        RECT 23.685 113.045 23.855 113.075 ;
        RECT 23.680 112.935 23.855 113.045 ;
        RECT 23.685 112.885 23.855 112.935 ;
        RECT 24.605 112.905 24.775 113.095 ;
        RECT 29.205 112.885 29.375 113.075 ;
        RECT 30.125 112.905 30.295 113.095 ;
        RECT 34.725 112.885 34.895 113.075 ;
        RECT 35.645 112.905 35.815 113.095 ;
        RECT 36.560 112.935 36.680 113.045 ;
        RECT 37.485 112.885 37.655 113.075 ;
        RECT 41.165 112.905 41.335 113.095 ;
        RECT 43.005 112.885 43.175 113.075 ;
        RECT 46.685 112.905 46.855 113.095 ;
        RECT 48.525 112.885 48.695 113.075 ;
        RECT 49.440 112.935 49.560 113.045 ;
        RECT 50.365 112.905 50.535 113.095 ;
        RECT 54.045 112.885 54.215 113.075 ;
        RECT 55.885 112.905 56.055 113.095 ;
        RECT 59.565 112.885 59.735 113.075 ;
        RECT 61.405 112.905 61.575 113.095 ;
        RECT 62.320 112.935 62.440 113.045 ;
        RECT 63.245 112.885 63.415 113.075 ;
        RECT 66.925 112.905 67.095 113.095 ;
        RECT 68.765 112.885 68.935 113.075 ;
        RECT 72.445 112.905 72.615 113.095 ;
        RECT 74.285 112.885 74.455 113.075 ;
        RECT 75.200 112.935 75.320 113.045 ;
        RECT 76.125 112.905 76.295 113.095 ;
        RECT 79.805 112.885 79.975 113.075 ;
        RECT 81.645 112.905 81.815 113.095 ;
        RECT 85.325 112.885 85.495 113.075 ;
        RECT 87.165 112.905 87.335 113.095 ;
        RECT 88.080 112.935 88.200 113.045 ;
        RECT 89.005 112.885 89.175 113.075 ;
        RECT 92.685 112.905 92.855 113.095 ;
        RECT 94.525 112.885 94.695 113.075 ;
        RECT 98.205 112.905 98.375 113.095 ;
        RECT 100.045 112.885 100.215 113.075 ;
        RECT 100.960 112.935 101.080 113.045 ;
        RECT 101.885 112.905 102.055 113.095 ;
        RECT 105.565 112.885 105.735 113.075 ;
        RECT 107.405 112.905 107.575 113.095 ;
        RECT 111.085 112.885 111.255 113.075 ;
        RECT 112.925 112.905 113.095 113.095 ;
        RECT 113.840 112.935 113.960 113.045 ;
        RECT 114.765 112.885 114.935 113.075 ;
        RECT 118.445 112.905 118.615 113.095 ;
        RECT 120.285 112.885 120.455 113.075 ;
        RECT 123.965 112.905 124.135 113.095 ;
        RECT 125.805 112.885 125.975 113.075 ;
        RECT 126.720 112.935 126.840 113.045 ;
        RECT 127.645 112.905 127.815 113.095 ;
        RECT 131.325 112.885 131.495 113.075 ;
        RECT 133.165 112.905 133.335 113.095 ;
        RECT 136.845 112.885 137.015 113.075 ;
        RECT 138.685 112.905 138.855 113.095 ;
        RECT 139.600 112.935 139.720 113.045 ;
        RECT 140.525 112.885 140.695 113.075 ;
        RECT 144.205 112.905 144.375 113.095 ;
        RECT 146.045 112.885 146.215 113.075 ;
        RECT 147.885 112.905 148.055 113.095 ;
        RECT 148.800 112.935 148.920 113.045 ;
        RECT 150.185 112.885 150.355 113.095 ;
        RECT 11.125 112.075 12.495 112.885 ;
        RECT 12.505 112.075 18.015 112.885 ;
        RECT 18.025 112.075 23.535 112.885 ;
        RECT 23.545 112.075 29.055 112.885 ;
        RECT 29.065 112.075 34.575 112.885 ;
        RECT 34.585 112.075 36.415 112.885 ;
        RECT 36.895 112.015 37.325 112.800 ;
        RECT 37.345 112.075 42.855 112.885 ;
        RECT 42.865 112.075 48.375 112.885 ;
        RECT 48.385 112.075 53.895 112.885 ;
        RECT 53.905 112.075 59.415 112.885 ;
        RECT 59.425 112.075 62.175 112.885 ;
        RECT 62.655 112.015 63.085 112.800 ;
        RECT 63.105 112.075 68.615 112.885 ;
        RECT 68.625 112.075 74.135 112.885 ;
        RECT 74.145 112.075 79.655 112.885 ;
        RECT 79.665 112.075 85.175 112.885 ;
        RECT 85.185 112.075 87.935 112.885 ;
        RECT 88.415 112.015 88.845 112.800 ;
        RECT 88.865 112.075 94.375 112.885 ;
        RECT 94.385 112.075 99.895 112.885 ;
        RECT 99.905 112.075 105.415 112.885 ;
        RECT 105.425 112.075 110.935 112.885 ;
        RECT 110.945 112.075 113.695 112.885 ;
        RECT 114.175 112.015 114.605 112.800 ;
        RECT 114.625 112.075 120.135 112.885 ;
        RECT 120.145 112.075 125.655 112.885 ;
        RECT 125.665 112.075 131.175 112.885 ;
        RECT 131.185 112.075 136.695 112.885 ;
        RECT 136.705 112.075 139.455 112.885 ;
        RECT 139.935 112.015 140.365 112.800 ;
        RECT 140.385 112.075 145.895 112.885 ;
        RECT 145.905 112.075 148.655 112.885 ;
        RECT 149.125 112.075 150.495 112.885 ;
      LAYER nwell ;
        RECT 10.930 108.855 150.690 111.685 ;
      LAYER pwell ;
        RECT 11.125 107.655 12.495 108.465 ;
        RECT 12.505 107.655 18.015 108.465 ;
        RECT 18.025 107.655 23.535 108.465 ;
        RECT 24.015 107.740 24.445 108.525 ;
        RECT 24.465 107.655 29.975 108.465 ;
        RECT 29.985 107.655 35.495 108.465 ;
        RECT 35.505 107.655 41.015 108.465 ;
        RECT 41.025 107.655 46.535 108.465 ;
        RECT 46.545 107.655 49.295 108.465 ;
        RECT 49.775 107.740 50.205 108.525 ;
        RECT 50.225 107.655 55.735 108.465 ;
        RECT 55.745 107.655 61.255 108.465 ;
        RECT 61.265 107.655 66.775 108.465 ;
        RECT 66.785 107.655 72.295 108.465 ;
        RECT 72.305 107.655 75.055 108.465 ;
        RECT 75.535 107.740 75.965 108.525 ;
        RECT 75.985 107.655 81.495 108.465 ;
        RECT 81.505 107.655 87.015 108.465 ;
        RECT 87.025 107.655 92.535 108.465 ;
        RECT 92.545 107.655 98.055 108.465 ;
        RECT 98.065 107.655 100.815 108.465 ;
        RECT 101.295 107.740 101.725 108.525 ;
        RECT 101.745 107.655 107.255 108.465 ;
        RECT 107.265 107.655 112.775 108.465 ;
        RECT 112.785 107.655 118.295 108.465 ;
        RECT 118.305 107.655 123.815 108.465 ;
        RECT 123.825 107.655 126.575 108.465 ;
        RECT 127.055 107.740 127.485 108.525 ;
        RECT 127.505 107.655 133.015 108.465 ;
        RECT 133.025 107.655 138.535 108.465 ;
        RECT 138.545 107.655 144.055 108.465 ;
        RECT 144.065 107.655 147.735 108.465 ;
        RECT 147.745 107.655 149.115 108.465 ;
        RECT 149.125 107.655 150.495 108.465 ;
        RECT 11.265 107.445 11.435 107.655 ;
        RECT 12.645 107.445 12.815 107.655 ;
        RECT 18.165 107.445 18.335 107.655 ;
        RECT 23.685 107.605 23.855 107.635 ;
        RECT 23.680 107.495 23.855 107.605 ;
        RECT 23.685 107.445 23.855 107.495 ;
        RECT 24.605 107.465 24.775 107.655 ;
        RECT 29.205 107.445 29.375 107.635 ;
        RECT 30.125 107.465 30.295 107.655 ;
        RECT 34.725 107.445 34.895 107.635 ;
        RECT 35.645 107.465 35.815 107.655 ;
        RECT 36.560 107.495 36.680 107.605 ;
        RECT 37.485 107.445 37.655 107.635 ;
        RECT 41.165 107.465 41.335 107.655 ;
        RECT 43.005 107.445 43.175 107.635 ;
        RECT 46.685 107.465 46.855 107.655 ;
        RECT 48.525 107.445 48.695 107.635 ;
        RECT 49.440 107.495 49.560 107.605 ;
        RECT 50.365 107.465 50.535 107.655 ;
        RECT 54.045 107.445 54.215 107.635 ;
        RECT 55.885 107.465 56.055 107.655 ;
        RECT 59.565 107.445 59.735 107.635 ;
        RECT 61.405 107.465 61.575 107.655 ;
        RECT 62.320 107.495 62.440 107.605 ;
        RECT 63.245 107.445 63.415 107.635 ;
        RECT 66.925 107.465 67.095 107.655 ;
        RECT 68.765 107.445 68.935 107.635 ;
        RECT 72.445 107.465 72.615 107.655 ;
        RECT 74.285 107.445 74.455 107.635 ;
        RECT 75.200 107.495 75.320 107.605 ;
        RECT 76.125 107.465 76.295 107.655 ;
        RECT 79.805 107.445 79.975 107.635 ;
        RECT 81.645 107.465 81.815 107.655 ;
        RECT 85.325 107.445 85.495 107.635 ;
        RECT 87.165 107.465 87.335 107.655 ;
        RECT 88.080 107.495 88.200 107.605 ;
        RECT 89.005 107.445 89.175 107.635 ;
        RECT 92.685 107.465 92.855 107.655 ;
        RECT 94.525 107.445 94.695 107.635 ;
        RECT 98.205 107.465 98.375 107.655 ;
        RECT 100.045 107.445 100.215 107.635 ;
        RECT 100.960 107.495 101.080 107.605 ;
        RECT 101.885 107.465 102.055 107.655 ;
        RECT 105.565 107.445 105.735 107.635 ;
        RECT 107.405 107.465 107.575 107.655 ;
        RECT 111.085 107.445 111.255 107.635 ;
        RECT 112.925 107.465 113.095 107.655 ;
        RECT 113.840 107.495 113.960 107.605 ;
        RECT 114.765 107.445 114.935 107.635 ;
        RECT 118.445 107.465 118.615 107.655 ;
        RECT 120.285 107.445 120.455 107.635 ;
        RECT 123.965 107.465 124.135 107.655 ;
        RECT 125.805 107.445 125.975 107.635 ;
        RECT 126.720 107.495 126.840 107.605 ;
        RECT 127.645 107.465 127.815 107.655 ;
        RECT 131.325 107.445 131.495 107.635 ;
        RECT 133.165 107.465 133.335 107.655 ;
        RECT 136.845 107.445 137.015 107.635 ;
        RECT 138.685 107.465 138.855 107.655 ;
        RECT 139.600 107.495 139.720 107.605 ;
        RECT 140.525 107.445 140.695 107.635 ;
        RECT 144.205 107.465 144.375 107.655 ;
        RECT 146.045 107.445 146.215 107.635 ;
        RECT 147.885 107.465 148.055 107.655 ;
        RECT 148.800 107.495 148.920 107.605 ;
        RECT 150.185 107.445 150.355 107.655 ;
        RECT 11.125 106.635 12.495 107.445 ;
        RECT 12.505 106.635 18.015 107.445 ;
        RECT 18.025 106.635 23.535 107.445 ;
        RECT 23.545 106.635 29.055 107.445 ;
        RECT 29.065 106.635 34.575 107.445 ;
        RECT 34.585 106.635 36.415 107.445 ;
        RECT 36.895 106.575 37.325 107.360 ;
        RECT 37.345 106.635 42.855 107.445 ;
        RECT 42.865 106.635 48.375 107.445 ;
        RECT 48.385 106.635 53.895 107.445 ;
        RECT 53.905 106.635 59.415 107.445 ;
        RECT 59.425 106.635 62.175 107.445 ;
        RECT 62.655 106.575 63.085 107.360 ;
        RECT 63.105 106.635 68.615 107.445 ;
        RECT 68.625 106.635 74.135 107.445 ;
        RECT 74.145 106.635 79.655 107.445 ;
        RECT 79.665 106.635 85.175 107.445 ;
        RECT 85.185 106.635 87.935 107.445 ;
        RECT 88.415 106.575 88.845 107.360 ;
        RECT 88.865 106.635 94.375 107.445 ;
        RECT 94.385 106.635 99.895 107.445 ;
        RECT 99.905 106.635 105.415 107.445 ;
        RECT 105.425 106.635 110.935 107.445 ;
        RECT 110.945 106.635 113.695 107.445 ;
        RECT 114.175 106.575 114.605 107.360 ;
        RECT 114.625 106.635 120.135 107.445 ;
        RECT 120.145 106.635 125.655 107.445 ;
        RECT 125.665 106.635 131.175 107.445 ;
        RECT 131.185 106.635 136.695 107.445 ;
        RECT 136.705 106.635 139.455 107.445 ;
        RECT 139.935 106.575 140.365 107.360 ;
        RECT 140.385 106.635 145.895 107.445 ;
        RECT 145.905 106.635 148.655 107.445 ;
        RECT 149.125 106.635 150.495 107.445 ;
      LAYER nwell ;
        RECT 10.930 103.415 150.690 106.245 ;
      LAYER pwell ;
        RECT 11.125 102.215 12.495 103.025 ;
        RECT 12.505 102.215 18.015 103.025 ;
        RECT 18.025 102.215 23.535 103.025 ;
        RECT 24.015 102.300 24.445 103.085 ;
        RECT 24.465 102.215 29.975 103.025 ;
        RECT 29.985 102.215 35.495 103.025 ;
        RECT 35.505 102.215 41.015 103.025 ;
        RECT 41.025 102.215 46.535 103.025 ;
        RECT 46.545 102.215 49.295 103.025 ;
        RECT 49.775 102.300 50.205 103.085 ;
        RECT 50.225 102.215 55.735 103.025 ;
        RECT 55.745 102.215 61.255 103.025 ;
        RECT 61.265 102.215 66.775 103.025 ;
        RECT 66.785 102.215 72.295 103.025 ;
        RECT 72.305 102.215 75.055 103.025 ;
        RECT 75.535 102.300 75.965 103.085 ;
        RECT 75.985 102.215 81.495 103.025 ;
        RECT 81.505 102.215 87.015 103.025 ;
        RECT 87.025 102.215 92.535 103.025 ;
        RECT 92.545 102.215 98.055 103.025 ;
        RECT 98.065 102.215 100.815 103.025 ;
        RECT 101.295 102.300 101.725 103.085 ;
        RECT 101.745 102.215 107.255 103.025 ;
        RECT 107.265 102.215 112.775 103.025 ;
        RECT 112.785 102.215 118.295 103.025 ;
        RECT 118.305 102.215 123.815 103.025 ;
        RECT 123.825 102.215 126.575 103.025 ;
        RECT 127.055 102.300 127.485 103.085 ;
        RECT 127.505 102.215 133.015 103.025 ;
        RECT 133.025 102.215 138.535 103.025 ;
        RECT 138.545 102.215 144.055 103.025 ;
        RECT 144.065 102.215 147.735 103.025 ;
        RECT 147.745 102.215 149.115 103.025 ;
        RECT 149.125 102.215 150.495 103.025 ;
        RECT 11.265 102.005 11.435 102.215 ;
        RECT 12.645 102.005 12.815 102.215 ;
        RECT 18.165 102.005 18.335 102.215 ;
        RECT 23.685 102.165 23.855 102.195 ;
        RECT 23.680 102.055 23.855 102.165 ;
        RECT 23.685 102.005 23.855 102.055 ;
        RECT 24.605 102.025 24.775 102.215 ;
        RECT 29.205 102.005 29.375 102.195 ;
        RECT 30.125 102.025 30.295 102.215 ;
        RECT 34.725 102.005 34.895 102.195 ;
        RECT 35.645 102.025 35.815 102.215 ;
        RECT 36.560 102.055 36.680 102.165 ;
        RECT 37.485 102.005 37.655 102.195 ;
        RECT 41.165 102.025 41.335 102.215 ;
        RECT 43.005 102.005 43.175 102.195 ;
        RECT 46.685 102.025 46.855 102.215 ;
        RECT 48.525 102.005 48.695 102.195 ;
        RECT 49.440 102.055 49.560 102.165 ;
        RECT 50.365 102.025 50.535 102.215 ;
        RECT 54.045 102.005 54.215 102.195 ;
        RECT 55.885 102.025 56.055 102.215 ;
        RECT 59.565 102.005 59.735 102.195 ;
        RECT 61.405 102.025 61.575 102.215 ;
        RECT 62.320 102.055 62.440 102.165 ;
        RECT 63.245 102.005 63.415 102.195 ;
        RECT 66.925 102.025 67.095 102.215 ;
        RECT 68.765 102.005 68.935 102.195 ;
        RECT 72.445 102.025 72.615 102.215 ;
        RECT 74.285 102.005 74.455 102.195 ;
        RECT 75.200 102.055 75.320 102.165 ;
        RECT 76.125 102.025 76.295 102.215 ;
        RECT 79.805 102.005 79.975 102.195 ;
        RECT 81.645 102.025 81.815 102.215 ;
        RECT 85.325 102.005 85.495 102.195 ;
        RECT 87.165 102.025 87.335 102.215 ;
        RECT 88.080 102.055 88.200 102.165 ;
        RECT 89.005 102.005 89.175 102.195 ;
        RECT 92.685 102.025 92.855 102.215 ;
        RECT 94.525 102.005 94.695 102.195 ;
        RECT 98.205 102.025 98.375 102.215 ;
        RECT 100.045 102.005 100.215 102.195 ;
        RECT 100.960 102.055 101.080 102.165 ;
        RECT 101.885 102.025 102.055 102.215 ;
        RECT 105.565 102.005 105.735 102.195 ;
        RECT 107.405 102.025 107.575 102.215 ;
        RECT 111.085 102.005 111.255 102.195 ;
        RECT 112.925 102.025 113.095 102.215 ;
        RECT 113.840 102.055 113.960 102.165 ;
        RECT 114.765 102.005 114.935 102.195 ;
        RECT 118.445 102.025 118.615 102.215 ;
        RECT 120.285 102.005 120.455 102.195 ;
        RECT 123.965 102.025 124.135 102.215 ;
        RECT 125.805 102.005 125.975 102.195 ;
        RECT 126.720 102.055 126.840 102.165 ;
        RECT 127.645 102.025 127.815 102.215 ;
        RECT 131.325 102.005 131.495 102.195 ;
        RECT 133.165 102.025 133.335 102.215 ;
        RECT 136.845 102.005 137.015 102.195 ;
        RECT 138.685 102.025 138.855 102.215 ;
        RECT 139.600 102.055 139.720 102.165 ;
        RECT 140.525 102.005 140.695 102.195 ;
        RECT 144.205 102.025 144.375 102.215 ;
        RECT 146.045 102.005 146.215 102.195 ;
        RECT 147.885 102.025 148.055 102.215 ;
        RECT 148.800 102.055 148.920 102.165 ;
        RECT 150.185 102.005 150.355 102.215 ;
        RECT 11.125 101.195 12.495 102.005 ;
        RECT 12.505 101.195 18.015 102.005 ;
        RECT 18.025 101.195 23.535 102.005 ;
        RECT 23.545 101.195 29.055 102.005 ;
        RECT 29.065 101.195 34.575 102.005 ;
        RECT 34.585 101.195 36.415 102.005 ;
        RECT 36.895 101.135 37.325 101.920 ;
        RECT 37.345 101.195 42.855 102.005 ;
        RECT 42.865 101.195 48.375 102.005 ;
        RECT 48.385 101.195 53.895 102.005 ;
        RECT 53.905 101.195 59.415 102.005 ;
        RECT 59.425 101.195 62.175 102.005 ;
        RECT 62.655 101.135 63.085 101.920 ;
        RECT 63.105 101.195 68.615 102.005 ;
        RECT 68.625 101.195 74.135 102.005 ;
        RECT 74.145 101.195 79.655 102.005 ;
        RECT 79.665 101.195 85.175 102.005 ;
        RECT 85.185 101.195 87.935 102.005 ;
        RECT 88.415 101.135 88.845 101.920 ;
        RECT 88.865 101.195 94.375 102.005 ;
        RECT 94.385 101.195 99.895 102.005 ;
        RECT 99.905 101.195 105.415 102.005 ;
        RECT 105.425 101.195 110.935 102.005 ;
        RECT 110.945 101.195 113.695 102.005 ;
        RECT 114.175 101.135 114.605 101.920 ;
        RECT 114.625 101.195 120.135 102.005 ;
        RECT 120.145 101.195 125.655 102.005 ;
        RECT 125.665 101.195 131.175 102.005 ;
        RECT 131.185 101.195 136.695 102.005 ;
        RECT 136.705 101.195 139.455 102.005 ;
        RECT 139.935 101.135 140.365 101.920 ;
        RECT 140.385 101.195 145.895 102.005 ;
        RECT 145.905 101.195 148.655 102.005 ;
        RECT 149.125 101.195 150.495 102.005 ;
      LAYER nwell ;
        RECT 10.930 97.975 150.690 100.805 ;
      LAYER pwell ;
        RECT 11.125 96.775 12.495 97.585 ;
        RECT 12.505 96.775 18.015 97.585 ;
        RECT 18.025 96.775 23.535 97.585 ;
        RECT 24.015 96.860 24.445 97.645 ;
        RECT 24.465 96.775 29.975 97.585 ;
        RECT 29.985 96.775 35.495 97.585 ;
        RECT 35.505 96.775 41.015 97.585 ;
        RECT 41.025 96.775 46.535 97.585 ;
        RECT 46.545 96.775 49.295 97.585 ;
        RECT 49.775 96.860 50.205 97.645 ;
        RECT 50.225 96.775 55.735 97.585 ;
        RECT 55.745 96.775 61.255 97.585 ;
        RECT 61.265 96.775 66.775 97.585 ;
        RECT 66.785 96.775 72.295 97.585 ;
        RECT 72.305 96.775 75.055 97.585 ;
        RECT 75.535 96.860 75.965 97.645 ;
        RECT 75.985 96.775 81.495 97.585 ;
        RECT 81.505 96.775 87.015 97.585 ;
        RECT 87.025 96.775 92.535 97.585 ;
        RECT 92.545 96.775 98.055 97.585 ;
        RECT 98.065 96.775 100.815 97.585 ;
        RECT 101.295 96.860 101.725 97.645 ;
        RECT 101.745 96.775 107.255 97.585 ;
        RECT 107.265 96.775 112.775 97.585 ;
        RECT 112.785 96.775 118.295 97.585 ;
        RECT 118.305 96.775 123.815 97.585 ;
        RECT 123.825 96.775 126.575 97.585 ;
        RECT 127.055 96.860 127.485 97.645 ;
        RECT 127.505 96.775 133.015 97.585 ;
        RECT 133.025 96.775 138.535 97.585 ;
        RECT 138.545 96.775 144.055 97.585 ;
        RECT 144.065 96.775 147.735 97.585 ;
        RECT 147.745 96.775 149.115 97.585 ;
        RECT 149.125 96.775 150.495 97.585 ;
        RECT 11.265 96.565 11.435 96.775 ;
        RECT 12.645 96.565 12.815 96.775 ;
        RECT 18.165 96.565 18.335 96.775 ;
        RECT 23.685 96.725 23.855 96.755 ;
        RECT 23.680 96.615 23.855 96.725 ;
        RECT 23.685 96.565 23.855 96.615 ;
        RECT 24.605 96.585 24.775 96.775 ;
        RECT 29.205 96.565 29.375 96.755 ;
        RECT 30.125 96.585 30.295 96.775 ;
        RECT 34.725 96.565 34.895 96.755 ;
        RECT 35.645 96.585 35.815 96.775 ;
        RECT 36.560 96.615 36.680 96.725 ;
        RECT 37.485 96.565 37.655 96.755 ;
        RECT 41.165 96.585 41.335 96.775 ;
        RECT 43.005 96.565 43.175 96.755 ;
        RECT 46.685 96.585 46.855 96.775 ;
        RECT 48.525 96.565 48.695 96.755 ;
        RECT 49.440 96.615 49.560 96.725 ;
        RECT 50.365 96.585 50.535 96.775 ;
        RECT 54.045 96.565 54.215 96.755 ;
        RECT 55.885 96.585 56.055 96.775 ;
        RECT 59.565 96.565 59.735 96.755 ;
        RECT 61.405 96.585 61.575 96.775 ;
        RECT 62.320 96.615 62.440 96.725 ;
        RECT 63.245 96.565 63.415 96.755 ;
        RECT 66.925 96.585 67.095 96.775 ;
        RECT 68.765 96.565 68.935 96.755 ;
        RECT 72.445 96.585 72.615 96.775 ;
        RECT 74.285 96.565 74.455 96.755 ;
        RECT 75.200 96.615 75.320 96.725 ;
        RECT 76.125 96.585 76.295 96.775 ;
        RECT 79.805 96.565 79.975 96.755 ;
        RECT 81.645 96.585 81.815 96.775 ;
        RECT 85.325 96.565 85.495 96.755 ;
        RECT 87.165 96.585 87.335 96.775 ;
        RECT 88.080 96.615 88.200 96.725 ;
        RECT 89.005 96.565 89.175 96.755 ;
        RECT 92.685 96.585 92.855 96.775 ;
        RECT 94.525 96.565 94.695 96.755 ;
        RECT 98.205 96.585 98.375 96.775 ;
        RECT 100.045 96.565 100.215 96.755 ;
        RECT 100.960 96.615 101.080 96.725 ;
        RECT 101.885 96.585 102.055 96.775 ;
        RECT 105.565 96.565 105.735 96.755 ;
        RECT 107.405 96.585 107.575 96.775 ;
        RECT 111.085 96.565 111.255 96.755 ;
        RECT 112.925 96.585 113.095 96.775 ;
        RECT 113.840 96.615 113.960 96.725 ;
        RECT 114.765 96.565 114.935 96.755 ;
        RECT 118.445 96.585 118.615 96.775 ;
        RECT 120.285 96.565 120.455 96.755 ;
        RECT 123.965 96.585 124.135 96.775 ;
        RECT 125.805 96.565 125.975 96.755 ;
        RECT 126.720 96.615 126.840 96.725 ;
        RECT 127.645 96.585 127.815 96.775 ;
        RECT 131.325 96.565 131.495 96.755 ;
        RECT 133.165 96.585 133.335 96.775 ;
        RECT 136.845 96.565 137.015 96.755 ;
        RECT 138.685 96.585 138.855 96.775 ;
        RECT 139.600 96.615 139.720 96.725 ;
        RECT 140.525 96.565 140.695 96.755 ;
        RECT 144.205 96.585 144.375 96.775 ;
        RECT 146.045 96.565 146.215 96.755 ;
        RECT 147.885 96.585 148.055 96.775 ;
        RECT 148.800 96.615 148.920 96.725 ;
        RECT 150.185 96.565 150.355 96.775 ;
        RECT 11.125 95.755 12.495 96.565 ;
        RECT 12.505 95.755 18.015 96.565 ;
        RECT 18.025 95.755 23.535 96.565 ;
        RECT 23.545 95.755 29.055 96.565 ;
        RECT 29.065 95.755 34.575 96.565 ;
        RECT 34.585 95.755 36.415 96.565 ;
        RECT 36.895 95.695 37.325 96.480 ;
        RECT 37.345 95.755 42.855 96.565 ;
        RECT 42.865 95.755 48.375 96.565 ;
        RECT 48.385 95.755 53.895 96.565 ;
        RECT 53.905 95.755 59.415 96.565 ;
        RECT 59.425 95.755 62.175 96.565 ;
        RECT 62.655 95.695 63.085 96.480 ;
        RECT 63.105 95.755 68.615 96.565 ;
        RECT 68.625 95.755 74.135 96.565 ;
        RECT 74.145 95.755 79.655 96.565 ;
        RECT 79.665 95.755 85.175 96.565 ;
        RECT 85.185 95.755 87.935 96.565 ;
        RECT 88.415 95.695 88.845 96.480 ;
        RECT 88.865 95.755 94.375 96.565 ;
        RECT 94.385 95.755 99.895 96.565 ;
        RECT 99.905 95.755 105.415 96.565 ;
        RECT 105.425 95.755 110.935 96.565 ;
        RECT 110.945 95.755 113.695 96.565 ;
        RECT 114.175 95.695 114.605 96.480 ;
        RECT 114.625 95.755 120.135 96.565 ;
        RECT 120.145 95.755 125.655 96.565 ;
        RECT 125.665 95.755 131.175 96.565 ;
        RECT 131.185 95.755 136.695 96.565 ;
        RECT 136.705 95.755 139.455 96.565 ;
        RECT 139.935 95.695 140.365 96.480 ;
        RECT 140.385 95.755 145.895 96.565 ;
        RECT 145.905 95.755 148.655 96.565 ;
        RECT 149.125 95.755 150.495 96.565 ;
      LAYER nwell ;
        RECT 10.930 92.535 150.690 95.365 ;
      LAYER pwell ;
        RECT 11.125 91.335 12.495 92.145 ;
        RECT 12.505 91.335 18.015 92.145 ;
        RECT 18.025 91.335 23.535 92.145 ;
        RECT 24.015 91.420 24.445 92.205 ;
        RECT 24.465 91.335 29.975 92.145 ;
        RECT 29.985 91.335 35.495 92.145 ;
        RECT 35.505 91.335 41.015 92.145 ;
        RECT 41.025 91.335 46.535 92.145 ;
        RECT 46.545 91.335 49.295 92.145 ;
        RECT 49.775 91.420 50.205 92.205 ;
        RECT 50.225 91.335 55.735 92.145 ;
        RECT 55.745 91.335 61.255 92.145 ;
        RECT 61.265 91.335 66.775 92.145 ;
        RECT 66.785 91.335 72.295 92.145 ;
        RECT 72.305 91.335 75.055 92.145 ;
        RECT 75.535 91.420 75.965 92.205 ;
        RECT 75.985 91.335 81.495 92.145 ;
        RECT 81.505 91.335 87.015 92.145 ;
        RECT 87.025 91.335 92.535 92.145 ;
        RECT 92.545 91.335 98.055 92.145 ;
        RECT 98.065 91.335 100.815 92.145 ;
        RECT 101.295 91.420 101.725 92.205 ;
        RECT 101.745 91.335 107.255 92.145 ;
        RECT 107.265 91.335 112.775 92.145 ;
        RECT 112.785 91.335 118.295 92.145 ;
        RECT 118.305 91.335 123.815 92.145 ;
        RECT 123.825 91.335 126.575 92.145 ;
        RECT 127.055 91.420 127.485 92.205 ;
        RECT 127.505 91.335 133.015 92.145 ;
        RECT 133.025 91.335 138.535 92.145 ;
        RECT 138.545 91.335 144.055 92.145 ;
        RECT 144.065 91.335 147.735 92.145 ;
        RECT 147.745 91.335 149.115 92.145 ;
        RECT 149.125 91.335 150.495 92.145 ;
        RECT 11.265 91.125 11.435 91.335 ;
        RECT 12.645 91.125 12.815 91.335 ;
        RECT 18.165 91.125 18.335 91.335 ;
        RECT 23.685 91.285 23.855 91.315 ;
        RECT 23.680 91.175 23.855 91.285 ;
        RECT 23.685 91.125 23.855 91.175 ;
        RECT 24.605 91.145 24.775 91.335 ;
        RECT 29.205 91.125 29.375 91.315 ;
        RECT 30.125 91.145 30.295 91.335 ;
        RECT 34.725 91.125 34.895 91.315 ;
        RECT 35.645 91.145 35.815 91.335 ;
        RECT 36.560 91.175 36.680 91.285 ;
        RECT 37.485 91.125 37.655 91.315 ;
        RECT 41.165 91.145 41.335 91.335 ;
        RECT 43.005 91.125 43.175 91.315 ;
        RECT 46.685 91.145 46.855 91.335 ;
        RECT 48.525 91.125 48.695 91.315 ;
        RECT 49.440 91.175 49.560 91.285 ;
        RECT 50.365 91.145 50.535 91.335 ;
        RECT 54.045 91.125 54.215 91.315 ;
        RECT 55.885 91.145 56.055 91.335 ;
        RECT 59.565 91.125 59.735 91.315 ;
        RECT 61.405 91.145 61.575 91.335 ;
        RECT 62.320 91.175 62.440 91.285 ;
        RECT 63.245 91.125 63.415 91.315 ;
        RECT 66.925 91.145 67.095 91.335 ;
        RECT 68.765 91.125 68.935 91.315 ;
        RECT 72.445 91.145 72.615 91.335 ;
        RECT 74.285 91.125 74.455 91.315 ;
        RECT 75.200 91.175 75.320 91.285 ;
        RECT 76.125 91.145 76.295 91.335 ;
        RECT 79.805 91.125 79.975 91.315 ;
        RECT 81.645 91.145 81.815 91.335 ;
        RECT 85.325 91.125 85.495 91.315 ;
        RECT 87.165 91.145 87.335 91.335 ;
        RECT 88.080 91.175 88.200 91.285 ;
        RECT 89.005 91.125 89.175 91.315 ;
        RECT 92.685 91.145 92.855 91.335 ;
        RECT 94.525 91.125 94.695 91.315 ;
        RECT 98.205 91.145 98.375 91.335 ;
        RECT 100.045 91.125 100.215 91.315 ;
        RECT 100.960 91.175 101.080 91.285 ;
        RECT 101.885 91.145 102.055 91.335 ;
        RECT 105.565 91.125 105.735 91.315 ;
        RECT 107.405 91.145 107.575 91.335 ;
        RECT 111.085 91.125 111.255 91.315 ;
        RECT 112.925 91.145 113.095 91.335 ;
        RECT 113.840 91.175 113.960 91.285 ;
        RECT 114.765 91.125 114.935 91.315 ;
        RECT 118.445 91.145 118.615 91.335 ;
        RECT 120.285 91.125 120.455 91.315 ;
        RECT 123.965 91.145 124.135 91.335 ;
        RECT 125.805 91.125 125.975 91.315 ;
        RECT 126.720 91.175 126.840 91.285 ;
        RECT 127.645 91.145 127.815 91.335 ;
        RECT 131.325 91.125 131.495 91.315 ;
        RECT 133.165 91.145 133.335 91.335 ;
        RECT 136.845 91.125 137.015 91.315 ;
        RECT 138.685 91.145 138.855 91.335 ;
        RECT 139.600 91.175 139.720 91.285 ;
        RECT 140.525 91.125 140.695 91.315 ;
        RECT 144.205 91.145 144.375 91.335 ;
        RECT 146.045 91.125 146.215 91.315 ;
        RECT 147.885 91.145 148.055 91.335 ;
        RECT 148.800 91.175 148.920 91.285 ;
        RECT 150.185 91.125 150.355 91.335 ;
        RECT 11.125 90.315 12.495 91.125 ;
        RECT 12.505 90.315 18.015 91.125 ;
        RECT 18.025 90.315 23.535 91.125 ;
        RECT 23.545 90.315 29.055 91.125 ;
        RECT 29.065 90.315 34.575 91.125 ;
        RECT 34.585 90.315 36.415 91.125 ;
        RECT 36.895 90.255 37.325 91.040 ;
        RECT 37.345 90.315 42.855 91.125 ;
        RECT 42.865 90.315 48.375 91.125 ;
        RECT 48.385 90.315 53.895 91.125 ;
        RECT 53.905 90.315 59.415 91.125 ;
        RECT 59.425 90.315 62.175 91.125 ;
        RECT 62.655 90.255 63.085 91.040 ;
        RECT 63.105 90.315 68.615 91.125 ;
        RECT 68.625 90.315 74.135 91.125 ;
        RECT 74.145 90.315 79.655 91.125 ;
        RECT 79.665 90.315 85.175 91.125 ;
        RECT 85.185 90.315 87.935 91.125 ;
        RECT 88.415 90.255 88.845 91.040 ;
        RECT 88.865 90.315 94.375 91.125 ;
        RECT 94.385 90.315 99.895 91.125 ;
        RECT 99.905 90.315 105.415 91.125 ;
        RECT 105.425 90.315 110.935 91.125 ;
        RECT 110.945 90.315 113.695 91.125 ;
        RECT 114.175 90.255 114.605 91.040 ;
        RECT 114.625 90.315 120.135 91.125 ;
        RECT 120.145 90.315 125.655 91.125 ;
        RECT 125.665 90.315 131.175 91.125 ;
        RECT 131.185 90.315 136.695 91.125 ;
        RECT 136.705 90.315 139.455 91.125 ;
        RECT 139.935 90.255 140.365 91.040 ;
        RECT 140.385 90.315 145.895 91.125 ;
        RECT 145.905 90.315 148.655 91.125 ;
        RECT 149.125 90.315 150.495 91.125 ;
      LAYER nwell ;
        RECT 10.930 87.095 150.690 89.925 ;
      LAYER pwell ;
        RECT 11.125 85.895 12.495 86.705 ;
        RECT 12.505 85.895 18.015 86.705 ;
        RECT 18.025 85.895 23.535 86.705 ;
        RECT 24.015 85.980 24.445 86.765 ;
        RECT 24.465 85.895 29.975 86.705 ;
        RECT 29.985 85.895 35.495 86.705 ;
        RECT 35.505 85.895 41.015 86.705 ;
        RECT 41.025 85.895 46.535 86.705 ;
        RECT 46.545 85.895 49.295 86.705 ;
        RECT 49.775 85.980 50.205 86.765 ;
        RECT 50.225 85.895 55.735 86.705 ;
        RECT 55.745 85.895 61.255 86.705 ;
        RECT 61.265 85.895 66.775 86.705 ;
        RECT 66.785 85.895 72.295 86.705 ;
        RECT 72.305 85.895 75.055 86.705 ;
        RECT 75.535 85.980 75.965 86.765 ;
        RECT 75.985 85.895 81.495 86.705 ;
        RECT 81.505 85.895 87.015 86.705 ;
        RECT 87.025 85.895 92.535 86.705 ;
        RECT 92.545 85.895 98.055 86.705 ;
        RECT 98.065 85.895 100.815 86.705 ;
        RECT 101.295 85.980 101.725 86.765 ;
        RECT 101.745 85.895 107.255 86.705 ;
        RECT 107.265 85.895 112.775 86.705 ;
        RECT 112.785 85.895 118.295 86.705 ;
        RECT 118.305 85.895 123.815 86.705 ;
        RECT 123.825 85.895 126.575 86.705 ;
        RECT 127.055 85.980 127.485 86.765 ;
        RECT 127.505 85.895 133.015 86.705 ;
        RECT 133.025 85.895 138.535 86.705 ;
        RECT 138.545 85.895 144.055 86.705 ;
        RECT 144.065 85.895 147.735 86.705 ;
        RECT 147.745 85.895 149.115 86.705 ;
        RECT 149.125 85.895 150.495 86.705 ;
        RECT 11.265 85.685 11.435 85.895 ;
        RECT 12.645 85.685 12.815 85.895 ;
        RECT 18.165 85.685 18.335 85.895 ;
        RECT 23.685 85.845 23.855 85.875 ;
        RECT 23.680 85.735 23.855 85.845 ;
        RECT 23.685 85.685 23.855 85.735 ;
        RECT 24.605 85.705 24.775 85.895 ;
        RECT 29.205 85.685 29.375 85.875 ;
        RECT 30.125 85.705 30.295 85.895 ;
        RECT 34.725 85.685 34.895 85.875 ;
        RECT 35.645 85.705 35.815 85.895 ;
        RECT 36.560 85.735 36.680 85.845 ;
        RECT 37.485 85.685 37.655 85.875 ;
        RECT 41.165 85.705 41.335 85.895 ;
        RECT 43.005 85.685 43.175 85.875 ;
        RECT 46.685 85.705 46.855 85.895 ;
        RECT 48.525 85.685 48.695 85.875 ;
        RECT 49.440 85.735 49.560 85.845 ;
        RECT 50.365 85.705 50.535 85.895 ;
        RECT 54.045 85.685 54.215 85.875 ;
        RECT 55.885 85.705 56.055 85.895 ;
        RECT 59.565 85.685 59.735 85.875 ;
        RECT 61.405 85.705 61.575 85.895 ;
        RECT 62.320 85.735 62.440 85.845 ;
        RECT 63.245 85.685 63.415 85.875 ;
        RECT 66.925 85.705 67.095 85.895 ;
        RECT 68.765 85.685 68.935 85.875 ;
        RECT 72.445 85.705 72.615 85.895 ;
        RECT 74.285 85.685 74.455 85.875 ;
        RECT 75.200 85.735 75.320 85.845 ;
        RECT 76.125 85.705 76.295 85.895 ;
        RECT 79.805 85.685 79.975 85.875 ;
        RECT 81.645 85.705 81.815 85.895 ;
        RECT 85.325 85.685 85.495 85.875 ;
        RECT 87.165 85.705 87.335 85.895 ;
        RECT 88.080 85.735 88.200 85.845 ;
        RECT 89.005 85.685 89.175 85.875 ;
        RECT 92.685 85.705 92.855 85.895 ;
        RECT 94.525 85.685 94.695 85.875 ;
        RECT 98.205 85.705 98.375 85.895 ;
        RECT 100.045 85.685 100.215 85.875 ;
        RECT 100.960 85.735 101.080 85.845 ;
        RECT 101.885 85.705 102.055 85.895 ;
        RECT 105.565 85.685 105.735 85.875 ;
        RECT 107.405 85.705 107.575 85.895 ;
        RECT 111.085 85.685 111.255 85.875 ;
        RECT 112.925 85.705 113.095 85.895 ;
        RECT 113.840 85.735 113.960 85.845 ;
        RECT 114.765 85.685 114.935 85.875 ;
        RECT 118.445 85.705 118.615 85.895 ;
        RECT 120.285 85.685 120.455 85.875 ;
        RECT 123.965 85.705 124.135 85.895 ;
        RECT 125.805 85.685 125.975 85.875 ;
        RECT 126.720 85.735 126.840 85.845 ;
        RECT 127.645 85.705 127.815 85.895 ;
        RECT 131.325 85.685 131.495 85.875 ;
        RECT 133.165 85.705 133.335 85.895 ;
        RECT 136.845 85.685 137.015 85.875 ;
        RECT 138.685 85.705 138.855 85.895 ;
        RECT 139.600 85.735 139.720 85.845 ;
        RECT 140.525 85.685 140.695 85.875 ;
        RECT 144.205 85.705 144.375 85.895 ;
        RECT 146.045 85.685 146.215 85.875 ;
        RECT 147.885 85.705 148.055 85.895 ;
        RECT 148.800 85.735 148.920 85.845 ;
        RECT 150.185 85.685 150.355 85.895 ;
        RECT 11.125 84.875 12.495 85.685 ;
        RECT 12.505 84.875 18.015 85.685 ;
        RECT 18.025 84.875 23.535 85.685 ;
        RECT 23.545 84.875 29.055 85.685 ;
        RECT 29.065 84.875 34.575 85.685 ;
        RECT 34.585 84.875 36.415 85.685 ;
        RECT 36.895 84.815 37.325 85.600 ;
        RECT 37.345 84.875 42.855 85.685 ;
        RECT 42.865 84.875 48.375 85.685 ;
        RECT 48.385 84.875 53.895 85.685 ;
        RECT 53.905 84.875 59.415 85.685 ;
        RECT 59.425 84.875 62.175 85.685 ;
        RECT 62.655 84.815 63.085 85.600 ;
        RECT 63.105 84.875 68.615 85.685 ;
        RECT 68.625 84.875 74.135 85.685 ;
        RECT 74.145 84.875 79.655 85.685 ;
        RECT 79.665 84.875 85.175 85.685 ;
        RECT 85.185 84.875 87.935 85.685 ;
        RECT 88.415 84.815 88.845 85.600 ;
        RECT 88.865 84.875 94.375 85.685 ;
        RECT 94.385 84.875 99.895 85.685 ;
        RECT 99.905 84.875 105.415 85.685 ;
        RECT 105.425 84.875 110.935 85.685 ;
        RECT 110.945 84.875 113.695 85.685 ;
        RECT 114.175 84.815 114.605 85.600 ;
        RECT 114.625 84.875 120.135 85.685 ;
        RECT 120.145 84.875 125.655 85.685 ;
        RECT 125.665 84.875 131.175 85.685 ;
        RECT 131.185 84.875 136.695 85.685 ;
        RECT 136.705 84.875 139.455 85.685 ;
        RECT 139.935 84.815 140.365 85.600 ;
        RECT 140.385 84.875 145.895 85.685 ;
        RECT 145.905 84.875 148.655 85.685 ;
        RECT 149.125 84.875 150.495 85.685 ;
      LAYER nwell ;
        RECT 10.930 81.655 150.690 84.485 ;
      LAYER pwell ;
        RECT 11.125 80.455 12.495 81.265 ;
        RECT 12.505 80.455 18.015 81.265 ;
        RECT 18.025 80.455 23.535 81.265 ;
        RECT 24.015 80.540 24.445 81.325 ;
        RECT 24.465 80.455 29.975 81.265 ;
        RECT 29.985 80.455 35.495 81.265 ;
        RECT 35.505 80.455 41.015 81.265 ;
        RECT 41.025 80.455 46.535 81.265 ;
        RECT 46.545 80.455 49.295 81.265 ;
        RECT 49.775 80.540 50.205 81.325 ;
        RECT 50.225 80.455 55.735 81.265 ;
        RECT 55.745 80.455 61.255 81.265 ;
        RECT 61.265 80.455 66.775 81.265 ;
        RECT 66.785 80.455 72.295 81.265 ;
        RECT 72.305 80.455 75.055 81.265 ;
        RECT 75.535 80.540 75.965 81.325 ;
        RECT 75.985 80.455 81.495 81.265 ;
        RECT 81.505 80.455 87.015 81.265 ;
        RECT 87.025 80.455 92.535 81.265 ;
        RECT 92.545 80.455 98.055 81.265 ;
        RECT 98.065 80.455 100.815 81.265 ;
        RECT 101.295 80.540 101.725 81.325 ;
        RECT 101.745 80.455 107.255 81.265 ;
        RECT 107.265 80.455 112.775 81.265 ;
        RECT 112.785 80.455 118.295 81.265 ;
        RECT 118.305 80.455 123.815 81.265 ;
        RECT 123.825 80.455 126.575 81.265 ;
        RECT 127.055 80.540 127.485 81.325 ;
        RECT 127.505 80.455 133.015 81.265 ;
        RECT 133.025 80.455 138.535 81.265 ;
        RECT 138.545 80.455 144.055 81.265 ;
        RECT 144.065 80.455 147.735 81.265 ;
        RECT 147.745 80.455 149.115 81.265 ;
        RECT 149.125 80.455 150.495 81.265 ;
        RECT 11.265 80.245 11.435 80.455 ;
        RECT 12.645 80.245 12.815 80.455 ;
        RECT 18.165 80.245 18.335 80.455 ;
        RECT 23.685 80.405 23.855 80.435 ;
        RECT 23.680 80.295 23.855 80.405 ;
        RECT 23.685 80.245 23.855 80.295 ;
        RECT 24.605 80.265 24.775 80.455 ;
        RECT 29.205 80.245 29.375 80.435 ;
        RECT 30.125 80.265 30.295 80.455 ;
        RECT 34.725 80.245 34.895 80.435 ;
        RECT 35.645 80.265 35.815 80.455 ;
        RECT 36.560 80.295 36.680 80.405 ;
        RECT 37.485 80.245 37.655 80.435 ;
        RECT 41.165 80.265 41.335 80.455 ;
        RECT 43.005 80.245 43.175 80.435 ;
        RECT 46.685 80.265 46.855 80.455 ;
        RECT 48.525 80.245 48.695 80.435 ;
        RECT 49.440 80.295 49.560 80.405 ;
        RECT 50.365 80.265 50.535 80.455 ;
        RECT 54.045 80.245 54.215 80.435 ;
        RECT 55.885 80.265 56.055 80.455 ;
        RECT 59.565 80.245 59.735 80.435 ;
        RECT 61.405 80.265 61.575 80.455 ;
        RECT 62.320 80.295 62.440 80.405 ;
        RECT 63.245 80.245 63.415 80.435 ;
        RECT 66.925 80.265 67.095 80.455 ;
        RECT 68.765 80.245 68.935 80.435 ;
        RECT 72.445 80.265 72.615 80.455 ;
        RECT 74.285 80.245 74.455 80.435 ;
        RECT 75.200 80.295 75.320 80.405 ;
        RECT 76.125 80.265 76.295 80.455 ;
        RECT 79.805 80.245 79.975 80.435 ;
        RECT 81.645 80.265 81.815 80.455 ;
        RECT 85.325 80.245 85.495 80.435 ;
        RECT 87.165 80.265 87.335 80.455 ;
        RECT 88.080 80.295 88.200 80.405 ;
        RECT 89.005 80.245 89.175 80.435 ;
        RECT 92.685 80.265 92.855 80.455 ;
        RECT 94.525 80.245 94.695 80.435 ;
        RECT 98.205 80.265 98.375 80.455 ;
        RECT 100.045 80.245 100.215 80.435 ;
        RECT 100.960 80.295 101.080 80.405 ;
        RECT 101.885 80.265 102.055 80.455 ;
        RECT 105.565 80.245 105.735 80.435 ;
        RECT 107.405 80.265 107.575 80.455 ;
        RECT 111.085 80.245 111.255 80.435 ;
        RECT 112.925 80.265 113.095 80.455 ;
        RECT 113.840 80.295 113.960 80.405 ;
        RECT 114.765 80.245 114.935 80.435 ;
        RECT 118.445 80.265 118.615 80.455 ;
        RECT 120.285 80.245 120.455 80.435 ;
        RECT 123.965 80.265 124.135 80.455 ;
        RECT 125.805 80.245 125.975 80.435 ;
        RECT 126.720 80.295 126.840 80.405 ;
        RECT 127.645 80.265 127.815 80.455 ;
        RECT 131.325 80.245 131.495 80.435 ;
        RECT 133.165 80.265 133.335 80.455 ;
        RECT 136.845 80.245 137.015 80.435 ;
        RECT 138.685 80.265 138.855 80.455 ;
        RECT 139.600 80.295 139.720 80.405 ;
        RECT 140.525 80.245 140.695 80.435 ;
        RECT 144.205 80.265 144.375 80.455 ;
        RECT 146.045 80.245 146.215 80.435 ;
        RECT 147.885 80.265 148.055 80.455 ;
        RECT 148.800 80.295 148.920 80.405 ;
        RECT 150.185 80.245 150.355 80.455 ;
        RECT 11.125 79.435 12.495 80.245 ;
        RECT 12.505 79.435 18.015 80.245 ;
        RECT 18.025 79.435 23.535 80.245 ;
        RECT 23.545 79.435 29.055 80.245 ;
        RECT 29.065 79.435 34.575 80.245 ;
        RECT 34.585 79.435 36.415 80.245 ;
        RECT 36.895 79.375 37.325 80.160 ;
        RECT 37.345 79.435 42.855 80.245 ;
        RECT 42.865 79.435 48.375 80.245 ;
        RECT 48.385 79.435 53.895 80.245 ;
        RECT 53.905 79.435 59.415 80.245 ;
        RECT 59.425 79.435 62.175 80.245 ;
        RECT 62.655 79.375 63.085 80.160 ;
        RECT 63.105 79.435 68.615 80.245 ;
        RECT 68.625 79.435 74.135 80.245 ;
        RECT 74.145 79.435 79.655 80.245 ;
        RECT 79.665 79.435 85.175 80.245 ;
        RECT 85.185 79.435 87.935 80.245 ;
        RECT 88.415 79.375 88.845 80.160 ;
        RECT 88.865 79.435 94.375 80.245 ;
        RECT 94.385 79.435 99.895 80.245 ;
        RECT 99.905 79.435 105.415 80.245 ;
        RECT 105.425 79.435 110.935 80.245 ;
        RECT 110.945 79.435 113.695 80.245 ;
        RECT 114.175 79.375 114.605 80.160 ;
        RECT 114.625 79.435 120.135 80.245 ;
        RECT 120.145 79.435 125.655 80.245 ;
        RECT 125.665 79.435 131.175 80.245 ;
        RECT 131.185 79.435 136.695 80.245 ;
        RECT 136.705 79.435 139.455 80.245 ;
        RECT 139.935 79.375 140.365 80.160 ;
        RECT 140.385 79.435 145.895 80.245 ;
        RECT 145.905 79.435 148.655 80.245 ;
        RECT 149.125 79.435 150.495 80.245 ;
      LAYER nwell ;
        RECT 10.930 76.215 150.690 79.045 ;
      LAYER pwell ;
        RECT 11.125 75.015 12.495 75.825 ;
        RECT 12.505 75.015 18.015 75.825 ;
        RECT 18.025 75.015 23.535 75.825 ;
        RECT 24.015 75.100 24.445 75.885 ;
        RECT 24.465 75.015 29.975 75.825 ;
        RECT 29.985 75.015 35.495 75.825 ;
        RECT 35.505 75.015 36.875 75.825 ;
        RECT 36.895 75.100 37.325 75.885 ;
        RECT 37.345 75.015 42.855 75.825 ;
        RECT 42.865 75.015 48.375 75.825 ;
        RECT 48.385 75.015 49.755 75.825 ;
        RECT 49.775 75.100 50.205 75.885 ;
        RECT 50.225 75.015 55.735 75.825 ;
        RECT 55.745 75.015 61.255 75.825 ;
        RECT 61.265 75.015 62.635 75.825 ;
        RECT 62.655 75.100 63.085 75.885 ;
        RECT 63.105 75.015 68.615 75.825 ;
        RECT 68.625 75.015 74.135 75.825 ;
        RECT 74.145 75.015 75.515 75.825 ;
        RECT 75.535 75.100 75.965 75.885 ;
        RECT 75.985 75.015 81.495 75.825 ;
        RECT 81.505 75.015 87.015 75.825 ;
        RECT 87.025 75.015 88.395 75.825 ;
        RECT 88.415 75.100 88.845 75.885 ;
        RECT 88.865 75.015 94.375 75.825 ;
        RECT 94.385 75.015 99.895 75.825 ;
        RECT 99.905 75.015 101.275 75.825 ;
        RECT 101.295 75.100 101.725 75.885 ;
        RECT 101.745 75.015 107.255 75.825 ;
        RECT 107.265 75.015 112.775 75.825 ;
        RECT 112.785 75.015 114.155 75.825 ;
        RECT 114.175 75.100 114.605 75.885 ;
        RECT 114.625 75.015 120.135 75.825 ;
        RECT 120.145 75.015 125.655 75.825 ;
        RECT 125.665 75.015 127.035 75.825 ;
        RECT 127.055 75.100 127.485 75.885 ;
        RECT 127.505 75.015 133.015 75.825 ;
        RECT 133.025 75.015 138.535 75.825 ;
        RECT 138.545 75.015 139.915 75.825 ;
        RECT 139.935 75.100 140.365 75.885 ;
        RECT 140.385 75.015 145.895 75.825 ;
        RECT 145.905 75.015 148.655 75.825 ;
        RECT 149.125 75.015 150.495 75.825 ;
        RECT 11.265 74.825 11.435 75.015 ;
        RECT 12.645 74.825 12.815 75.015 ;
        RECT 18.165 74.825 18.335 75.015 ;
        RECT 23.680 74.855 23.800 74.965 ;
        RECT 24.605 74.825 24.775 75.015 ;
        RECT 30.125 74.825 30.295 75.015 ;
        RECT 35.645 74.825 35.815 75.015 ;
        RECT 37.485 74.825 37.655 75.015 ;
        RECT 43.005 74.825 43.175 75.015 ;
        RECT 48.525 74.825 48.695 75.015 ;
        RECT 50.365 74.825 50.535 75.015 ;
        RECT 55.885 74.825 56.055 75.015 ;
        RECT 61.405 74.825 61.575 75.015 ;
        RECT 63.245 74.825 63.415 75.015 ;
        RECT 68.765 74.825 68.935 75.015 ;
        RECT 74.285 74.825 74.455 75.015 ;
        RECT 76.125 74.825 76.295 75.015 ;
        RECT 81.645 74.825 81.815 75.015 ;
        RECT 87.165 74.825 87.335 75.015 ;
        RECT 89.005 74.825 89.175 75.015 ;
        RECT 94.525 74.825 94.695 75.015 ;
        RECT 100.045 74.825 100.215 75.015 ;
        RECT 101.885 74.825 102.055 75.015 ;
        RECT 107.405 74.825 107.575 75.015 ;
        RECT 112.925 74.825 113.095 75.015 ;
        RECT 114.765 74.825 114.935 75.015 ;
        RECT 120.285 74.825 120.455 75.015 ;
        RECT 125.805 74.825 125.975 75.015 ;
        RECT 127.645 74.825 127.815 75.015 ;
        RECT 133.165 74.825 133.335 75.015 ;
        RECT 138.685 74.825 138.855 75.015 ;
        RECT 140.525 74.825 140.695 75.015 ;
        RECT 146.045 74.825 146.215 75.015 ;
        RECT 148.800 74.855 148.920 74.965 ;
        RECT 150.185 74.825 150.355 75.015 ;
      LAYER nwell ;
        RECT 60.880 34.830 66.730 50.240 ;
      LAYER pwell ;
        RECT 61.590 29.860 65.980 34.460 ;
        RECT 54.850 24.420 65.680 27.520 ;
        RECT 72.510 25.370 75.610 43.070 ;
      LAYER nwell ;
        RECT 77.650 32.760 80.840 50.230 ;
      LAYER pwell ;
        RECT 99.400 41.360 101.410 49.980 ;
        RECT 94.790 37.040 105.620 40.140 ;
      LAYER nwell ;
        RECT 123.110 34.430 128.960 49.840 ;
      LAYER pwell ;
        RECT 123.820 29.460 128.210 34.060 ;
        RECT 117.080 24.020 127.910 27.120 ;
        RECT 134.740 24.970 137.840 42.670 ;
      LAYER nwell ;
        RECT 139.880 32.360 143.070 49.830 ;
      LAYER li1 ;
        RECT 11.120 213.545 150.500 213.715 ;
        RECT 11.205 212.455 12.415 213.545 ;
        RECT 12.585 213.110 17.930 213.545 ;
        RECT 18.105 213.110 23.450 213.545 ;
        RECT 11.205 211.745 11.725 212.285 ;
        RECT 11.895 211.915 12.415 212.455 ;
        RECT 11.205 210.995 12.415 211.745 ;
        RECT 14.170 211.540 14.510 212.370 ;
        RECT 15.990 211.860 16.340 213.110 ;
        RECT 19.690 211.540 20.030 212.370 ;
        RECT 21.510 211.860 21.860 213.110 ;
        RECT 24.085 212.380 24.375 213.545 ;
        RECT 24.545 213.110 29.890 213.545 ;
        RECT 30.065 213.110 35.410 213.545 ;
        RECT 12.585 210.995 17.930 211.540 ;
        RECT 18.105 210.995 23.450 211.540 ;
        RECT 24.085 210.995 24.375 211.720 ;
        RECT 26.130 211.540 26.470 212.370 ;
        RECT 27.950 211.860 28.300 213.110 ;
        RECT 31.650 211.540 31.990 212.370 ;
        RECT 33.470 211.860 33.820 213.110 ;
        RECT 35.585 212.455 36.795 213.545 ;
        RECT 35.585 211.745 36.105 212.285 ;
        RECT 36.275 211.915 36.795 212.455 ;
        RECT 36.965 212.380 37.255 213.545 ;
        RECT 37.425 213.110 42.770 213.545 ;
        RECT 42.945 213.110 48.290 213.545 ;
        RECT 24.545 210.995 29.890 211.540 ;
        RECT 30.065 210.995 35.410 211.540 ;
        RECT 35.585 210.995 36.795 211.745 ;
        RECT 36.965 210.995 37.255 211.720 ;
        RECT 39.010 211.540 39.350 212.370 ;
        RECT 40.830 211.860 41.180 213.110 ;
        RECT 44.530 211.540 44.870 212.370 ;
        RECT 46.350 211.860 46.700 213.110 ;
        RECT 48.465 212.455 49.675 213.545 ;
        RECT 48.465 211.745 48.985 212.285 ;
        RECT 49.155 211.915 49.675 212.455 ;
        RECT 49.845 212.380 50.135 213.545 ;
        RECT 50.305 213.110 55.650 213.545 ;
        RECT 55.825 213.110 61.170 213.545 ;
        RECT 37.425 210.995 42.770 211.540 ;
        RECT 42.945 210.995 48.290 211.540 ;
        RECT 48.465 210.995 49.675 211.745 ;
        RECT 49.845 210.995 50.135 211.720 ;
        RECT 51.890 211.540 52.230 212.370 ;
        RECT 53.710 211.860 54.060 213.110 ;
        RECT 57.410 211.540 57.750 212.370 ;
        RECT 59.230 211.860 59.580 213.110 ;
        RECT 61.345 212.455 62.555 213.545 ;
        RECT 61.345 211.745 61.865 212.285 ;
        RECT 62.035 211.915 62.555 212.455 ;
        RECT 62.725 212.380 63.015 213.545 ;
        RECT 64.195 212.615 64.365 213.375 ;
        RECT 64.580 212.785 64.910 213.545 ;
        RECT 64.195 212.445 64.910 212.615 ;
        RECT 65.080 212.470 65.335 213.375 ;
        RECT 64.105 211.895 64.460 212.265 ;
        RECT 64.740 212.235 64.910 212.445 ;
        RECT 64.740 211.905 64.995 212.235 ;
        RECT 50.305 210.995 55.650 211.540 ;
        RECT 55.825 210.995 61.170 211.540 ;
        RECT 61.345 210.995 62.555 211.745 ;
        RECT 62.725 210.995 63.015 211.720 ;
        RECT 64.740 211.715 64.910 211.905 ;
        RECT 65.165 211.740 65.335 212.470 ;
        RECT 65.510 212.395 65.770 213.545 ;
        RECT 65.945 213.110 71.290 213.545 ;
        RECT 64.195 211.545 64.910 211.715 ;
        RECT 64.195 211.165 64.365 211.545 ;
        RECT 64.580 210.995 64.910 211.375 ;
        RECT 65.080 211.165 65.335 211.740 ;
        RECT 65.510 210.995 65.770 211.835 ;
        RECT 67.530 211.540 67.870 212.370 ;
        RECT 69.350 211.860 69.700 213.110 ;
        RECT 71.465 212.455 74.975 213.545 ;
        RECT 71.465 211.765 73.115 212.285 ;
        RECT 73.285 211.935 74.975 212.455 ;
        RECT 75.605 212.380 75.895 213.545 ;
        RECT 76.065 213.110 81.410 213.545 ;
        RECT 65.945 210.995 71.290 211.540 ;
        RECT 71.465 210.995 74.975 211.765 ;
        RECT 75.605 210.995 75.895 211.720 ;
        RECT 77.650 211.540 77.990 212.370 ;
        RECT 79.470 211.860 79.820 213.110 ;
        RECT 81.585 212.455 85.095 213.545 ;
        RECT 85.265 212.455 86.475 213.545 ;
        RECT 81.585 211.765 83.235 212.285 ;
        RECT 83.405 211.935 85.095 212.455 ;
        RECT 76.065 210.995 81.410 211.540 ;
        RECT 81.585 210.995 85.095 211.765 ;
        RECT 85.265 211.745 85.785 212.285 ;
        RECT 85.955 211.915 86.475 212.455 ;
        RECT 86.735 212.615 86.905 213.375 ;
        RECT 87.085 212.785 87.415 213.545 ;
        RECT 86.735 212.445 87.400 212.615 ;
        RECT 87.585 212.470 87.855 213.375 ;
        RECT 87.230 212.300 87.400 212.445 ;
        RECT 86.665 211.895 86.995 212.265 ;
        RECT 87.230 211.970 87.515 212.300 ;
        RECT 85.265 210.995 86.475 211.745 ;
        RECT 87.230 211.715 87.400 211.970 ;
        RECT 86.735 211.545 87.400 211.715 ;
        RECT 87.685 211.670 87.855 212.470 ;
        RECT 88.485 212.380 88.775 213.545 ;
        RECT 88.945 213.110 94.290 213.545 ;
        RECT 86.735 211.165 86.905 211.545 ;
        RECT 87.085 210.995 87.415 211.375 ;
        RECT 87.595 211.165 87.855 211.670 ;
        RECT 88.485 210.995 88.775 211.720 ;
        RECT 90.530 211.540 90.870 212.370 ;
        RECT 92.350 211.860 92.700 213.110 ;
        RECT 94.465 212.455 96.135 213.545 ;
        RECT 94.465 211.765 95.215 212.285 ;
        RECT 95.385 211.935 96.135 212.455 ;
        RECT 96.395 212.615 96.565 213.375 ;
        RECT 96.745 212.785 97.075 213.545 ;
        RECT 96.395 212.445 97.060 212.615 ;
        RECT 97.245 212.470 97.515 213.375 ;
        RECT 96.890 212.300 97.060 212.445 ;
        RECT 96.325 211.895 96.655 212.265 ;
        RECT 96.890 211.970 97.175 212.300 ;
        RECT 88.945 210.995 94.290 211.540 ;
        RECT 94.465 210.995 96.135 211.765 ;
        RECT 96.890 211.715 97.060 211.970 ;
        RECT 96.395 211.545 97.060 211.715 ;
        RECT 97.345 211.670 97.515 212.470 ;
        RECT 97.685 212.455 101.195 213.545 ;
        RECT 96.395 211.165 96.565 211.545 ;
        RECT 96.745 210.995 97.075 211.375 ;
        RECT 97.255 211.165 97.515 211.670 ;
        RECT 97.685 211.765 99.335 212.285 ;
        RECT 99.505 211.935 101.195 212.455 ;
        RECT 101.365 212.380 101.655 213.545 ;
        RECT 101.825 212.455 104.415 213.545 ;
        RECT 104.700 212.915 104.985 213.375 ;
        RECT 105.155 213.085 105.425 213.545 ;
        RECT 104.700 212.695 105.655 212.915 ;
        RECT 101.825 211.765 103.035 212.285 ;
        RECT 103.205 211.935 104.415 212.455 ;
        RECT 104.585 211.965 105.275 212.525 ;
        RECT 105.445 211.795 105.655 212.695 ;
        RECT 97.685 210.995 101.195 211.765 ;
        RECT 101.365 210.995 101.655 211.720 ;
        RECT 101.825 210.995 104.415 211.765 ;
        RECT 104.700 211.625 105.655 211.795 ;
        RECT 105.825 212.525 106.225 213.375 ;
        RECT 106.415 212.915 106.695 213.375 ;
        RECT 107.215 213.085 107.540 213.545 ;
        RECT 106.415 212.695 107.540 212.915 ;
        RECT 105.825 211.965 106.920 212.525 ;
        RECT 107.090 212.235 107.540 212.695 ;
        RECT 107.710 212.405 108.095 213.375 ;
        RECT 108.325 212.405 108.535 213.545 ;
        RECT 104.700 211.165 104.985 211.625 ;
        RECT 105.155 210.995 105.425 211.455 ;
        RECT 105.825 211.165 106.225 211.965 ;
        RECT 107.090 211.905 107.645 212.235 ;
        RECT 107.090 211.795 107.540 211.905 ;
        RECT 106.415 211.625 107.540 211.795 ;
        RECT 107.815 211.735 108.095 212.405 ;
        RECT 108.705 212.395 109.035 213.375 ;
        RECT 109.205 212.405 109.435 213.545 ;
        RECT 109.645 212.470 109.915 213.375 ;
        RECT 110.085 212.785 110.415 213.545 ;
        RECT 110.595 212.615 110.765 213.375 ;
        RECT 106.415 211.165 106.695 211.625 ;
        RECT 107.215 210.995 107.540 211.455 ;
        RECT 107.710 211.165 108.095 211.735 ;
        RECT 108.325 210.995 108.535 211.815 ;
        RECT 108.705 211.795 108.955 212.395 ;
        RECT 109.125 211.985 109.455 212.235 ;
        RECT 108.705 211.165 109.035 211.795 ;
        RECT 109.205 210.995 109.435 211.815 ;
        RECT 109.645 211.670 109.815 212.470 ;
        RECT 110.100 212.445 110.765 212.615 ;
        RECT 111.025 212.455 113.615 213.545 ;
        RECT 110.100 212.300 110.270 212.445 ;
        RECT 109.985 211.970 110.270 212.300 ;
        RECT 110.100 211.715 110.270 211.970 ;
        RECT 110.505 211.895 110.835 212.265 ;
        RECT 111.025 211.765 112.235 212.285 ;
        RECT 112.405 211.935 113.615 212.455 ;
        RECT 114.245 212.380 114.535 213.545 ;
        RECT 114.705 212.455 116.375 213.545 ;
        RECT 114.705 211.765 115.455 212.285 ;
        RECT 115.625 211.935 116.375 212.455 ;
        RECT 116.545 212.470 116.815 213.375 ;
        RECT 116.985 212.785 117.315 213.545 ;
        RECT 117.495 212.615 117.665 213.375 ;
        RECT 117.925 213.110 123.270 213.545 ;
        RECT 109.645 211.165 109.905 211.670 ;
        RECT 110.100 211.545 110.765 211.715 ;
        RECT 110.085 210.995 110.415 211.375 ;
        RECT 110.595 211.165 110.765 211.545 ;
        RECT 111.025 210.995 113.615 211.765 ;
        RECT 114.245 210.995 114.535 211.720 ;
        RECT 114.705 210.995 116.375 211.765 ;
        RECT 116.545 211.670 116.715 212.470 ;
        RECT 117.000 212.445 117.665 212.615 ;
        RECT 117.000 212.300 117.170 212.445 ;
        RECT 116.885 211.970 117.170 212.300 ;
        RECT 117.000 211.715 117.170 211.970 ;
        RECT 117.405 211.895 117.735 212.265 ;
        RECT 116.545 211.165 116.805 211.670 ;
        RECT 117.000 211.545 117.665 211.715 ;
        RECT 116.985 210.995 117.315 211.375 ;
        RECT 117.495 211.165 117.665 211.545 ;
        RECT 119.510 211.540 119.850 212.370 ;
        RECT 121.330 211.860 121.680 213.110 ;
        RECT 123.445 212.455 126.955 213.545 ;
        RECT 123.445 211.765 125.095 212.285 ;
        RECT 125.265 211.935 126.955 212.455 ;
        RECT 127.125 212.380 127.415 213.545 ;
        RECT 127.585 212.470 127.855 213.375 ;
        RECT 128.025 212.785 128.355 213.545 ;
        RECT 128.535 212.615 128.705 213.375 ;
        RECT 128.965 213.110 134.310 213.545 ;
        RECT 117.925 210.995 123.270 211.540 ;
        RECT 123.445 210.995 126.955 211.765 ;
        RECT 127.125 210.995 127.415 211.720 ;
        RECT 127.585 211.670 127.755 212.470 ;
        RECT 128.040 212.445 128.705 212.615 ;
        RECT 128.040 212.300 128.210 212.445 ;
        RECT 127.925 211.970 128.210 212.300 ;
        RECT 128.040 211.715 128.210 211.970 ;
        RECT 128.445 211.895 128.775 212.265 ;
        RECT 127.585 211.165 127.845 211.670 ;
        RECT 128.040 211.545 128.705 211.715 ;
        RECT 128.025 210.995 128.355 211.375 ;
        RECT 128.535 211.165 128.705 211.545 ;
        RECT 130.550 211.540 130.890 212.370 ;
        RECT 132.370 211.860 132.720 213.110 ;
        RECT 134.485 212.455 136.155 213.545 ;
        RECT 134.485 211.765 135.235 212.285 ;
        RECT 135.405 211.935 136.155 212.455 ;
        RECT 136.785 212.575 137.095 213.375 ;
        RECT 137.265 212.745 137.575 213.545 ;
        RECT 137.745 212.915 138.005 213.375 ;
        RECT 138.175 213.085 138.430 213.545 ;
        RECT 138.605 212.915 138.865 213.375 ;
        RECT 137.745 212.745 138.865 212.915 ;
        RECT 136.785 212.405 137.815 212.575 ;
        RECT 128.965 210.995 134.310 211.540 ;
        RECT 134.485 210.995 136.155 211.765 ;
        RECT 136.785 211.495 136.955 212.405 ;
        RECT 137.125 211.665 137.475 212.235 ;
        RECT 137.645 212.155 137.815 212.405 ;
        RECT 138.605 212.495 138.865 212.745 ;
        RECT 139.035 212.675 139.320 213.545 ;
        RECT 138.605 212.325 139.360 212.495 ;
        RECT 140.005 212.380 140.295 213.545 ;
        RECT 140.465 213.110 145.810 213.545 ;
        RECT 137.645 211.985 138.785 212.155 ;
        RECT 138.955 211.815 139.360 212.325 ;
        RECT 137.710 211.645 139.360 211.815 ;
        RECT 136.785 211.165 137.085 211.495 ;
        RECT 137.255 210.995 137.530 211.475 ;
        RECT 137.710 211.255 138.005 211.645 ;
        RECT 138.175 210.995 138.430 211.475 ;
        RECT 138.605 211.255 138.865 211.645 ;
        RECT 139.035 210.995 139.315 211.475 ;
        RECT 140.005 210.995 140.295 211.720 ;
        RECT 142.050 211.540 142.390 212.370 ;
        RECT 143.870 211.860 144.220 213.110 ;
        RECT 145.985 212.455 148.575 213.545 ;
        RECT 145.985 211.765 147.195 212.285 ;
        RECT 147.365 211.935 148.575 212.455 ;
        RECT 149.205 212.455 150.415 213.545 ;
        RECT 149.205 211.915 149.725 212.455 ;
        RECT 140.465 210.995 145.810 211.540 ;
        RECT 145.985 210.995 148.575 211.765 ;
        RECT 149.895 211.745 150.415 212.285 ;
        RECT 149.205 210.995 150.415 211.745 ;
        RECT 11.120 210.825 150.500 210.995 ;
        RECT 11.205 210.075 12.415 210.825 ;
        RECT 11.205 209.535 11.725 210.075 ;
        RECT 12.585 210.055 15.175 210.825 ;
        RECT 15.405 210.345 15.685 210.825 ;
        RECT 15.855 210.175 16.115 210.565 ;
        RECT 16.290 210.345 16.545 210.825 ;
        RECT 16.715 210.175 17.010 210.565 ;
        RECT 17.190 210.345 17.465 210.825 ;
        RECT 17.635 210.325 17.935 210.655 ;
        RECT 11.895 209.365 12.415 209.905 ;
        RECT 12.585 209.535 13.795 210.055 ;
        RECT 15.360 210.005 17.010 210.175 ;
        RECT 13.965 209.365 15.175 209.885 ;
        RECT 11.205 208.275 12.415 209.365 ;
        RECT 12.585 208.275 15.175 209.365 ;
        RECT 15.360 209.495 15.765 210.005 ;
        RECT 15.935 209.665 17.075 209.835 ;
        RECT 15.360 209.325 16.115 209.495 ;
        RECT 15.400 208.275 15.685 209.145 ;
        RECT 15.855 209.075 16.115 209.325 ;
        RECT 16.905 209.415 17.075 209.665 ;
        RECT 17.245 209.585 17.595 210.155 ;
        RECT 17.765 209.415 17.935 210.325 ;
        RECT 18.105 210.055 19.775 210.825 ;
        RECT 20.035 210.275 20.205 210.565 ;
        RECT 20.375 210.445 20.705 210.825 ;
        RECT 20.035 210.105 20.700 210.275 ;
        RECT 18.105 209.535 18.855 210.055 ;
        RECT 16.905 209.245 17.935 209.415 ;
        RECT 19.025 209.365 19.775 209.885 ;
        RECT 15.855 208.905 16.975 209.075 ;
        RECT 15.855 208.445 16.115 208.905 ;
        RECT 16.290 208.275 16.545 208.735 ;
        RECT 16.715 208.445 16.975 208.905 ;
        RECT 17.145 208.275 17.455 209.075 ;
        RECT 17.625 208.445 17.935 209.245 ;
        RECT 18.105 208.275 19.775 209.365 ;
        RECT 19.950 209.285 20.300 209.935 ;
        RECT 20.470 209.115 20.700 210.105 ;
        RECT 20.035 208.945 20.700 209.115 ;
        RECT 20.035 208.445 20.205 208.945 ;
        RECT 20.375 208.275 20.705 208.775 ;
        RECT 20.875 208.445 21.060 210.565 ;
        RECT 21.315 210.365 21.565 210.825 ;
        RECT 21.735 210.375 22.070 210.545 ;
        RECT 22.265 210.375 22.940 210.545 ;
        RECT 21.735 210.235 21.905 210.375 ;
        RECT 21.230 209.245 21.510 210.195 ;
        RECT 21.680 210.105 21.905 210.235 ;
        RECT 21.680 209.000 21.850 210.105 ;
        RECT 22.075 209.955 22.600 210.175 ;
        RECT 22.020 209.190 22.260 209.785 ;
        RECT 22.430 209.255 22.600 209.955 ;
        RECT 22.770 209.595 22.940 210.375 ;
        RECT 23.260 210.325 23.630 210.825 ;
        RECT 23.810 210.375 24.215 210.545 ;
        RECT 24.385 210.375 25.170 210.545 ;
        RECT 23.810 210.145 23.980 210.375 ;
        RECT 23.150 209.845 23.980 210.145 ;
        RECT 24.365 209.875 24.830 210.205 ;
        RECT 23.150 209.815 23.350 209.845 ;
        RECT 23.470 209.595 23.640 209.665 ;
        RECT 22.770 209.425 23.640 209.595 ;
        RECT 23.130 209.335 23.640 209.425 ;
        RECT 21.680 208.870 21.985 209.000 ;
        RECT 22.430 208.890 22.960 209.255 ;
        RECT 21.300 208.275 21.565 208.735 ;
        RECT 21.735 208.445 21.985 208.870 ;
        RECT 23.130 208.720 23.300 209.335 ;
        RECT 22.195 208.550 23.300 208.720 ;
        RECT 23.470 208.275 23.640 209.075 ;
        RECT 23.810 208.775 23.980 209.845 ;
        RECT 24.150 208.945 24.340 209.665 ;
        RECT 24.510 208.915 24.830 209.875 ;
        RECT 25.000 209.915 25.170 210.375 ;
        RECT 25.445 210.295 25.655 210.825 ;
        RECT 25.915 210.085 26.245 210.610 ;
        RECT 26.415 210.215 26.585 210.825 ;
        RECT 26.755 210.170 27.085 210.605 ;
        RECT 27.365 210.345 27.645 210.825 ;
        RECT 27.815 210.175 28.075 210.565 ;
        RECT 28.250 210.345 28.505 210.825 ;
        RECT 28.675 210.175 28.970 210.565 ;
        RECT 29.150 210.345 29.425 210.825 ;
        RECT 29.595 210.325 29.895 210.655 ;
        RECT 26.755 210.085 27.135 210.170 ;
        RECT 26.045 209.915 26.245 210.085 ;
        RECT 26.910 210.045 27.135 210.085 ;
        RECT 25.000 209.585 25.875 209.915 ;
        RECT 26.045 209.585 26.795 209.915 ;
        RECT 23.810 208.445 24.060 208.775 ;
        RECT 25.000 208.745 25.170 209.585 ;
        RECT 26.045 209.380 26.235 209.585 ;
        RECT 26.965 209.465 27.135 210.045 ;
        RECT 26.920 209.415 27.135 209.465 ;
        RECT 25.340 209.005 26.235 209.380 ;
        RECT 26.745 209.335 27.135 209.415 ;
        RECT 27.320 210.005 28.970 210.175 ;
        RECT 27.320 209.495 27.725 210.005 ;
        RECT 27.895 209.665 29.035 209.835 ;
        RECT 24.285 208.575 25.170 208.745 ;
        RECT 25.350 208.275 25.665 208.775 ;
        RECT 25.895 208.445 26.235 209.005 ;
        RECT 26.405 208.275 26.575 209.285 ;
        RECT 26.745 208.490 27.075 209.335 ;
        RECT 27.320 209.325 28.075 209.495 ;
        RECT 27.360 208.275 27.645 209.145 ;
        RECT 27.815 209.075 28.075 209.325 ;
        RECT 28.865 209.415 29.035 209.665 ;
        RECT 29.205 209.585 29.555 210.155 ;
        RECT 29.725 209.415 29.895 210.325 ;
        RECT 28.865 209.245 29.895 209.415 ;
        RECT 27.815 208.905 28.935 209.075 ;
        RECT 27.815 208.445 28.075 208.905 ;
        RECT 28.250 208.275 28.505 208.735 ;
        RECT 28.675 208.445 28.935 208.905 ;
        RECT 29.105 208.275 29.415 209.075 ;
        RECT 29.585 208.445 29.895 209.245 ;
        RECT 30.560 210.085 31.175 210.655 ;
        RECT 31.345 210.315 31.560 210.825 ;
        RECT 31.790 210.315 32.070 210.645 ;
        RECT 32.250 210.315 32.490 210.825 ;
        RECT 30.560 209.065 30.875 210.085 ;
        RECT 31.045 209.415 31.215 209.915 ;
        RECT 31.465 209.585 31.730 210.145 ;
        RECT 31.900 209.415 32.070 210.315 ;
        RECT 32.240 209.585 32.595 210.145 ;
        RECT 32.825 210.025 33.520 210.655 ;
        RECT 33.725 210.025 34.035 210.825 ;
        RECT 34.265 210.345 34.545 210.825 ;
        RECT 34.715 210.175 34.975 210.565 ;
        RECT 35.150 210.345 35.405 210.825 ;
        RECT 35.575 210.175 35.870 210.565 ;
        RECT 36.050 210.345 36.325 210.825 ;
        RECT 36.495 210.325 36.795 210.655 ;
        RECT 32.845 209.585 33.180 209.835 ;
        RECT 33.350 209.425 33.520 210.025 ;
        RECT 34.220 210.005 35.870 210.175 ;
        RECT 33.690 209.585 34.025 209.855 ;
        RECT 34.220 209.495 34.625 210.005 ;
        RECT 34.795 209.665 35.935 209.835 ;
        RECT 31.045 209.245 32.470 209.415 ;
        RECT 30.560 208.445 31.095 209.065 ;
        RECT 31.265 208.275 31.595 209.075 ;
        RECT 32.080 209.070 32.470 209.245 ;
        RECT 32.825 208.275 33.085 209.415 ;
        RECT 33.255 208.445 33.585 209.425 ;
        RECT 33.755 208.275 34.035 209.415 ;
        RECT 34.220 209.325 34.975 209.495 ;
        RECT 34.260 208.275 34.545 209.145 ;
        RECT 34.715 209.075 34.975 209.325 ;
        RECT 35.765 209.415 35.935 209.665 ;
        RECT 36.105 209.585 36.455 210.155 ;
        RECT 36.625 209.415 36.795 210.325 ;
        RECT 36.965 210.100 37.255 210.825 ;
        RECT 37.425 210.150 37.685 210.655 ;
        RECT 37.865 210.445 38.195 210.825 ;
        RECT 38.375 210.275 38.545 210.655 ;
        RECT 35.765 209.245 36.795 209.415 ;
        RECT 34.715 208.905 35.835 209.075 ;
        RECT 34.715 208.445 34.975 208.905 ;
        RECT 35.150 208.275 35.405 208.735 ;
        RECT 35.575 208.445 35.835 208.905 ;
        RECT 36.005 208.275 36.315 209.075 ;
        RECT 36.485 208.445 36.795 209.245 ;
        RECT 36.965 208.275 37.255 209.440 ;
        RECT 37.425 209.350 37.595 210.150 ;
        RECT 37.880 210.105 38.545 210.275 ;
        RECT 37.880 209.850 38.050 210.105 ;
        RECT 39.265 210.085 39.730 210.630 ;
        RECT 37.765 209.520 38.050 209.850 ;
        RECT 38.285 209.555 38.615 209.925 ;
        RECT 37.880 209.375 38.050 209.520 ;
        RECT 37.425 208.445 37.695 209.350 ;
        RECT 37.880 209.205 38.545 209.375 ;
        RECT 37.865 208.275 38.195 209.035 ;
        RECT 38.375 208.445 38.545 209.205 ;
        RECT 39.265 209.125 39.435 210.085 ;
        RECT 40.235 210.005 40.405 210.825 ;
        RECT 40.575 210.175 40.905 210.655 ;
        RECT 41.075 210.435 41.425 210.825 ;
        RECT 41.595 210.255 41.825 210.655 ;
        RECT 41.315 210.175 41.825 210.255 ;
        RECT 40.575 210.085 41.825 210.175 ;
        RECT 41.995 210.085 42.315 210.565 ;
        RECT 42.545 210.345 42.825 210.825 ;
        RECT 42.995 210.175 43.255 210.565 ;
        RECT 43.430 210.345 43.685 210.825 ;
        RECT 43.855 210.175 44.150 210.565 ;
        RECT 44.330 210.345 44.605 210.825 ;
        RECT 44.775 210.325 45.075 210.655 ;
        RECT 40.575 210.005 41.485 210.085 ;
        RECT 39.605 209.465 39.850 209.915 ;
        RECT 40.110 209.635 40.805 209.835 ;
        RECT 40.975 209.665 41.575 209.835 ;
        RECT 40.975 209.465 41.145 209.665 ;
        RECT 41.805 209.495 41.975 209.915 ;
        RECT 39.605 209.295 41.145 209.465 ;
        RECT 41.315 209.325 41.975 209.495 ;
        RECT 41.315 209.125 41.485 209.325 ;
        RECT 42.145 209.155 42.315 210.085 ;
        RECT 42.500 210.005 44.150 210.175 ;
        RECT 42.500 209.495 42.905 210.005 ;
        RECT 43.075 209.665 44.215 209.835 ;
        RECT 42.500 209.325 43.255 209.495 ;
        RECT 39.265 208.955 41.485 209.125 ;
        RECT 41.655 208.955 42.315 209.155 ;
        RECT 39.265 208.275 39.565 208.785 ;
        RECT 39.735 208.445 40.065 208.955 ;
        RECT 41.655 208.785 41.825 208.955 ;
        RECT 40.235 208.275 40.865 208.785 ;
        RECT 41.445 208.615 41.825 208.785 ;
        RECT 41.995 208.275 42.295 208.785 ;
        RECT 42.540 208.275 42.825 209.145 ;
        RECT 42.995 209.075 43.255 209.325 ;
        RECT 44.045 209.415 44.215 209.665 ;
        RECT 44.385 209.585 44.735 210.155 ;
        RECT 44.905 209.415 45.075 210.325 ;
        RECT 44.045 209.245 45.075 209.415 ;
        RECT 43.465 209.075 43.635 209.125 ;
        RECT 42.995 208.905 44.115 209.075 ;
        RECT 42.995 208.445 43.255 208.905 ;
        RECT 43.430 208.275 43.685 208.735 ;
        RECT 43.855 208.445 44.115 208.905 ;
        RECT 44.285 208.275 44.595 209.075 ;
        RECT 44.765 208.445 45.075 209.245 ;
        RECT 45.245 210.085 45.710 210.630 ;
        RECT 45.245 209.125 45.415 210.085 ;
        RECT 46.215 210.005 46.385 210.825 ;
        RECT 46.555 210.175 46.885 210.655 ;
        RECT 47.055 210.435 47.405 210.825 ;
        RECT 47.575 210.255 47.805 210.655 ;
        RECT 47.295 210.175 47.805 210.255 ;
        RECT 46.555 210.085 47.805 210.175 ;
        RECT 47.975 210.085 48.295 210.565 ;
        RECT 48.515 210.435 48.845 210.825 ;
        RECT 49.015 210.255 49.185 210.575 ;
        RECT 49.355 210.435 49.685 210.825 ;
        RECT 50.100 210.425 51.055 210.595 ;
        RECT 46.555 210.005 47.465 210.085 ;
        RECT 45.585 209.465 45.830 209.915 ;
        RECT 46.090 209.635 46.785 209.835 ;
        RECT 46.955 209.665 47.555 209.835 ;
        RECT 46.955 209.465 47.125 209.665 ;
        RECT 47.785 209.495 47.955 209.915 ;
        RECT 45.585 209.295 47.125 209.465 ;
        RECT 47.295 209.325 47.955 209.495 ;
        RECT 47.295 209.125 47.465 209.325 ;
        RECT 48.125 209.155 48.295 210.085 ;
        RECT 45.245 208.955 47.465 209.125 ;
        RECT 47.635 208.955 48.295 209.155 ;
        RECT 48.465 210.085 50.715 210.255 ;
        RECT 48.465 209.125 48.635 210.085 ;
        RECT 48.805 209.465 49.050 209.915 ;
        RECT 49.220 209.635 49.770 209.835 ;
        RECT 49.940 209.665 50.315 209.835 ;
        RECT 49.940 209.465 50.110 209.665 ;
        RECT 50.485 209.585 50.715 210.085 ;
        RECT 48.805 209.295 50.110 209.465 ;
        RECT 50.885 209.545 51.055 210.425 ;
        RECT 51.225 209.990 51.515 210.825 ;
        RECT 52.145 210.085 52.610 210.630 ;
        RECT 50.885 209.375 51.515 209.545 ;
        RECT 45.245 208.275 45.545 208.785 ;
        RECT 45.715 208.445 46.045 208.955 ;
        RECT 47.635 208.785 47.805 208.955 ;
        RECT 46.215 208.275 46.845 208.785 ;
        RECT 47.425 208.615 47.805 208.785 ;
        RECT 47.975 208.275 48.275 208.785 ;
        RECT 48.465 208.445 48.845 209.125 ;
        RECT 49.435 208.275 49.605 209.125 ;
        RECT 49.775 208.955 51.015 209.125 ;
        RECT 49.775 208.445 50.105 208.955 ;
        RECT 50.275 208.275 50.445 208.785 ;
        RECT 50.615 208.445 51.015 208.955 ;
        RECT 51.195 208.445 51.515 209.375 ;
        RECT 52.145 209.125 52.315 210.085 ;
        RECT 53.115 210.005 53.285 210.825 ;
        RECT 53.455 210.175 53.785 210.655 ;
        RECT 53.955 210.435 54.305 210.825 ;
        RECT 54.475 210.255 54.705 210.655 ;
        RECT 54.195 210.175 54.705 210.255 ;
        RECT 53.455 210.085 54.705 210.175 ;
        RECT 54.875 210.085 55.195 210.565 ;
        RECT 55.455 210.275 55.625 210.565 ;
        RECT 55.795 210.445 56.125 210.825 ;
        RECT 55.455 210.105 56.120 210.275 ;
        RECT 53.455 210.005 54.365 210.085 ;
        RECT 52.485 209.465 52.730 209.915 ;
        RECT 52.990 209.635 53.685 209.835 ;
        RECT 53.855 209.665 54.455 209.835 ;
        RECT 53.855 209.465 54.025 209.665 ;
        RECT 54.685 209.495 54.855 209.915 ;
        RECT 52.485 209.295 54.025 209.465 ;
        RECT 54.195 209.325 54.855 209.495 ;
        RECT 54.195 209.125 54.365 209.325 ;
        RECT 55.025 209.155 55.195 210.085 ;
        RECT 55.370 209.285 55.720 209.935 ;
        RECT 52.145 208.955 54.365 209.125 ;
        RECT 54.535 208.955 55.195 209.155 ;
        RECT 55.890 209.115 56.120 210.105 ;
        RECT 52.145 208.275 52.445 208.785 ;
        RECT 52.615 208.445 52.945 208.955 ;
        RECT 54.535 208.785 54.705 208.955 ;
        RECT 55.455 208.945 56.120 209.115 ;
        RECT 53.115 208.275 53.745 208.785 ;
        RECT 54.325 208.615 54.705 208.785 ;
        RECT 54.875 208.275 55.175 208.785 ;
        RECT 55.455 208.445 55.625 208.945 ;
        RECT 55.795 208.275 56.125 208.775 ;
        RECT 56.295 208.445 56.480 210.565 ;
        RECT 56.735 210.365 56.985 210.825 ;
        RECT 57.155 210.375 57.490 210.545 ;
        RECT 57.685 210.375 58.360 210.545 ;
        RECT 57.155 210.235 57.325 210.375 ;
        RECT 56.650 209.245 56.930 210.195 ;
        RECT 57.100 210.105 57.325 210.235 ;
        RECT 57.100 209.000 57.270 210.105 ;
        RECT 57.495 209.955 58.020 210.175 ;
        RECT 57.440 209.190 57.680 209.785 ;
        RECT 57.850 209.255 58.020 209.955 ;
        RECT 58.190 209.595 58.360 210.375 ;
        RECT 58.680 210.325 59.050 210.825 ;
        RECT 59.230 210.375 59.635 210.545 ;
        RECT 59.805 210.375 60.590 210.545 ;
        RECT 59.230 210.145 59.400 210.375 ;
        RECT 58.570 209.845 59.400 210.145 ;
        RECT 59.785 209.875 60.250 210.205 ;
        RECT 58.570 209.815 58.770 209.845 ;
        RECT 58.890 209.595 59.060 209.665 ;
        RECT 58.190 209.425 59.060 209.595 ;
        RECT 58.550 209.335 59.060 209.425 ;
        RECT 57.100 208.870 57.405 209.000 ;
        RECT 57.850 208.890 58.380 209.255 ;
        RECT 56.720 208.275 56.985 208.735 ;
        RECT 57.155 208.445 57.405 208.870 ;
        RECT 58.550 208.720 58.720 209.335 ;
        RECT 57.615 208.550 58.720 208.720 ;
        RECT 58.890 208.275 59.060 209.075 ;
        RECT 59.230 208.775 59.400 209.845 ;
        RECT 59.570 208.945 59.760 209.665 ;
        RECT 59.930 208.915 60.250 209.875 ;
        RECT 60.420 209.915 60.590 210.375 ;
        RECT 60.865 210.295 61.075 210.825 ;
        RECT 61.335 210.085 61.665 210.610 ;
        RECT 61.835 210.215 62.005 210.825 ;
        RECT 62.175 210.170 62.505 210.605 ;
        RECT 62.175 210.085 62.555 210.170 ;
        RECT 62.725 210.100 63.015 210.825 ;
        RECT 64.195 210.275 64.365 210.565 ;
        RECT 64.535 210.445 64.865 210.825 ;
        RECT 64.195 210.105 64.860 210.275 ;
        RECT 61.465 209.915 61.665 210.085 ;
        RECT 62.330 210.045 62.555 210.085 ;
        RECT 60.420 209.585 61.295 209.915 ;
        RECT 61.465 209.585 62.215 209.915 ;
        RECT 59.230 208.445 59.480 208.775 ;
        RECT 60.420 208.745 60.590 209.585 ;
        RECT 61.465 209.380 61.655 209.585 ;
        RECT 62.385 209.465 62.555 210.045 ;
        RECT 62.340 209.415 62.555 209.465 ;
        RECT 60.760 209.005 61.655 209.380 ;
        RECT 62.165 209.335 62.555 209.415 ;
        RECT 59.705 208.575 60.590 208.745 ;
        RECT 60.770 208.275 61.085 208.775 ;
        RECT 61.315 208.445 61.655 209.005 ;
        RECT 61.825 208.275 61.995 209.285 ;
        RECT 62.165 208.490 62.495 209.335 ;
        RECT 62.725 208.275 63.015 209.440 ;
        RECT 64.110 209.285 64.460 209.935 ;
        RECT 64.630 209.115 64.860 210.105 ;
        RECT 64.195 208.945 64.860 209.115 ;
        RECT 64.195 208.445 64.365 208.945 ;
        RECT 64.535 208.275 64.865 208.775 ;
        RECT 65.035 208.445 65.220 210.565 ;
        RECT 65.475 210.365 65.725 210.825 ;
        RECT 65.895 210.375 66.230 210.545 ;
        RECT 66.425 210.375 67.100 210.545 ;
        RECT 65.895 210.235 66.065 210.375 ;
        RECT 65.390 209.245 65.670 210.195 ;
        RECT 65.840 210.105 66.065 210.235 ;
        RECT 65.840 209.000 66.010 210.105 ;
        RECT 66.235 209.955 66.760 210.175 ;
        RECT 66.180 209.190 66.420 209.785 ;
        RECT 66.590 209.255 66.760 209.955 ;
        RECT 66.930 209.595 67.100 210.375 ;
        RECT 67.420 210.325 67.790 210.825 ;
        RECT 67.970 210.375 68.375 210.545 ;
        RECT 68.545 210.375 69.330 210.545 ;
        RECT 67.970 210.145 68.140 210.375 ;
        RECT 67.310 209.845 68.140 210.145 ;
        RECT 68.525 209.875 68.990 210.205 ;
        RECT 67.310 209.815 67.510 209.845 ;
        RECT 67.630 209.595 67.800 209.665 ;
        RECT 66.930 209.425 67.800 209.595 ;
        RECT 67.290 209.335 67.800 209.425 ;
        RECT 65.840 208.870 66.145 209.000 ;
        RECT 66.590 208.890 67.120 209.255 ;
        RECT 65.460 208.275 65.725 208.735 ;
        RECT 65.895 208.445 66.145 208.870 ;
        RECT 67.290 208.720 67.460 209.335 ;
        RECT 66.355 208.550 67.460 208.720 ;
        RECT 67.630 208.275 67.800 209.075 ;
        RECT 67.970 208.775 68.140 209.845 ;
        RECT 68.310 208.945 68.500 209.665 ;
        RECT 68.670 208.915 68.990 209.875 ;
        RECT 69.160 209.915 69.330 210.375 ;
        RECT 69.605 210.295 69.815 210.825 ;
        RECT 70.075 210.085 70.405 210.610 ;
        RECT 70.575 210.215 70.745 210.825 ;
        RECT 70.915 210.170 71.245 210.605 ;
        RECT 71.465 210.325 71.765 210.655 ;
        RECT 71.935 210.345 72.210 210.825 ;
        RECT 70.915 210.085 71.295 210.170 ;
        RECT 70.205 209.915 70.405 210.085 ;
        RECT 71.070 210.045 71.295 210.085 ;
        RECT 69.160 209.585 70.035 209.915 ;
        RECT 70.205 209.585 70.955 209.915 ;
        RECT 67.970 208.445 68.220 208.775 ;
        RECT 69.160 208.745 69.330 209.585 ;
        RECT 70.205 209.380 70.395 209.585 ;
        RECT 71.125 209.465 71.295 210.045 ;
        RECT 71.080 209.415 71.295 209.465 ;
        RECT 69.500 209.005 70.395 209.380 ;
        RECT 70.905 209.335 71.295 209.415 ;
        RECT 71.465 209.415 71.635 210.325 ;
        RECT 72.390 210.175 72.685 210.565 ;
        RECT 72.855 210.345 73.110 210.825 ;
        RECT 73.285 210.175 73.545 210.565 ;
        RECT 73.715 210.345 73.995 210.825 ;
        RECT 74.315 210.275 74.485 210.565 ;
        RECT 74.655 210.445 74.985 210.825 ;
        RECT 71.805 209.585 72.155 210.155 ;
        RECT 72.390 210.005 74.040 210.175 ;
        RECT 74.315 210.105 74.980 210.275 ;
        RECT 72.325 209.665 73.465 209.835 ;
        RECT 72.325 209.415 72.495 209.665 ;
        RECT 73.635 209.495 74.040 210.005 ;
        RECT 68.445 208.575 69.330 208.745 ;
        RECT 69.510 208.275 69.825 208.775 ;
        RECT 70.055 208.445 70.395 209.005 ;
        RECT 70.565 208.275 70.735 209.285 ;
        RECT 70.905 208.490 71.235 209.335 ;
        RECT 71.465 209.245 72.495 209.415 ;
        RECT 73.285 209.325 74.040 209.495 ;
        RECT 71.465 208.445 71.775 209.245 ;
        RECT 73.285 209.075 73.545 209.325 ;
        RECT 74.230 209.285 74.580 209.935 ;
        RECT 71.945 208.275 72.255 209.075 ;
        RECT 72.425 208.905 73.545 209.075 ;
        RECT 72.425 208.445 72.685 208.905 ;
        RECT 72.855 208.275 73.110 208.735 ;
        RECT 73.285 208.445 73.545 208.905 ;
        RECT 73.715 208.275 74.000 209.145 ;
        RECT 74.750 209.115 74.980 210.105 ;
        RECT 74.315 208.945 74.980 209.115 ;
        RECT 74.315 208.445 74.485 208.945 ;
        RECT 74.655 208.275 74.985 208.775 ;
        RECT 75.155 208.445 75.340 210.565 ;
        RECT 75.595 210.365 75.845 210.825 ;
        RECT 76.015 210.375 76.350 210.545 ;
        RECT 76.545 210.375 77.220 210.545 ;
        RECT 76.015 210.235 76.185 210.375 ;
        RECT 75.510 209.245 75.790 210.195 ;
        RECT 75.960 210.105 76.185 210.235 ;
        RECT 75.960 209.000 76.130 210.105 ;
        RECT 76.355 209.955 76.880 210.175 ;
        RECT 76.300 209.190 76.540 209.785 ;
        RECT 76.710 209.255 76.880 209.955 ;
        RECT 77.050 209.595 77.220 210.375 ;
        RECT 77.540 210.325 77.910 210.825 ;
        RECT 78.090 210.375 78.495 210.545 ;
        RECT 78.665 210.375 79.450 210.545 ;
        RECT 78.090 210.145 78.260 210.375 ;
        RECT 77.430 209.845 78.260 210.145 ;
        RECT 78.645 209.875 79.110 210.205 ;
        RECT 77.430 209.815 77.630 209.845 ;
        RECT 77.750 209.595 77.920 209.665 ;
        RECT 77.050 209.425 77.920 209.595 ;
        RECT 77.410 209.335 77.920 209.425 ;
        RECT 75.960 208.870 76.265 209.000 ;
        RECT 76.710 208.890 77.240 209.255 ;
        RECT 75.580 208.275 75.845 208.735 ;
        RECT 76.015 208.445 76.265 208.870 ;
        RECT 77.410 208.720 77.580 209.335 ;
        RECT 76.475 208.550 77.580 208.720 ;
        RECT 77.750 208.275 77.920 209.075 ;
        RECT 78.090 208.775 78.260 209.845 ;
        RECT 78.430 208.945 78.620 209.665 ;
        RECT 78.790 208.915 79.110 209.875 ;
        RECT 79.280 209.915 79.450 210.375 ;
        RECT 79.725 210.295 79.935 210.825 ;
        RECT 80.195 210.085 80.525 210.610 ;
        RECT 80.695 210.215 80.865 210.825 ;
        RECT 81.035 210.170 81.365 210.605 ;
        RECT 81.035 210.085 81.415 210.170 ;
        RECT 80.325 209.915 80.525 210.085 ;
        RECT 81.190 210.045 81.415 210.085 ;
        RECT 79.280 209.585 80.155 209.915 ;
        RECT 80.325 209.585 81.075 209.915 ;
        RECT 78.090 208.445 78.340 208.775 ;
        RECT 79.280 208.745 79.450 209.585 ;
        RECT 80.325 209.380 80.515 209.585 ;
        RECT 81.245 209.465 81.415 210.045 ;
        RECT 81.585 210.005 81.845 210.825 ;
        RECT 82.015 210.005 82.345 210.425 ;
        RECT 82.525 210.340 83.315 210.605 ;
        RECT 82.095 209.915 82.345 210.005 ;
        RECT 81.200 209.415 81.415 209.465 ;
        RECT 79.620 209.005 80.515 209.380 ;
        RECT 81.025 209.335 81.415 209.415 ;
        RECT 78.565 208.575 79.450 208.745 ;
        RECT 79.630 208.275 79.945 208.775 ;
        RECT 80.175 208.445 80.515 209.005 ;
        RECT 80.685 208.275 80.855 209.285 ;
        RECT 81.025 208.490 81.355 209.335 ;
        RECT 81.585 208.955 81.925 209.835 ;
        RECT 82.095 209.665 82.890 209.915 ;
        RECT 81.585 208.275 81.845 208.785 ;
        RECT 82.095 208.445 82.265 209.665 ;
        RECT 83.060 209.485 83.315 210.340 ;
        RECT 83.485 210.185 83.685 210.605 ;
        RECT 83.875 210.365 84.205 210.825 ;
        RECT 83.485 209.665 83.895 210.185 ;
        RECT 84.375 210.175 84.635 210.655 ;
        RECT 84.065 209.485 84.295 209.915 ;
        RECT 82.505 209.315 84.295 209.485 ;
        RECT 82.505 208.950 82.755 209.315 ;
        RECT 82.925 208.955 83.255 209.145 ;
        RECT 83.475 209.020 84.190 209.315 ;
        RECT 84.465 209.145 84.635 210.175 ;
        RECT 82.925 208.780 83.120 208.955 ;
        RECT 82.505 208.275 83.120 208.780 ;
        RECT 83.290 208.445 83.765 208.785 ;
        RECT 83.935 208.275 84.150 208.820 ;
        RECT 84.360 208.445 84.635 209.145 ;
        RECT 84.805 210.325 85.105 210.655 ;
        RECT 85.275 210.345 85.550 210.825 ;
        RECT 84.805 209.415 84.975 210.325 ;
        RECT 85.730 210.175 86.025 210.565 ;
        RECT 86.195 210.345 86.450 210.825 ;
        RECT 86.625 210.175 86.885 210.565 ;
        RECT 87.055 210.345 87.335 210.825 ;
        RECT 85.145 209.585 85.495 210.155 ;
        RECT 85.730 210.005 87.380 210.175 ;
        RECT 88.485 210.100 88.775 210.825 ;
        RECT 89.035 210.275 89.205 210.565 ;
        RECT 89.375 210.445 89.705 210.825 ;
        RECT 89.035 210.105 89.700 210.275 ;
        RECT 85.665 209.665 86.805 209.835 ;
        RECT 85.665 209.415 85.835 209.665 ;
        RECT 86.975 209.495 87.380 210.005 ;
        RECT 84.805 209.245 85.835 209.415 ;
        RECT 86.625 209.325 87.380 209.495 ;
        RECT 84.805 208.445 85.115 209.245 ;
        RECT 86.625 209.075 86.885 209.325 ;
        RECT 85.285 208.275 85.595 209.075 ;
        RECT 85.765 208.905 86.885 209.075 ;
        RECT 85.765 208.445 86.025 208.905 ;
        RECT 86.195 208.275 86.450 208.735 ;
        RECT 86.625 208.445 86.885 208.905 ;
        RECT 87.055 208.275 87.340 209.145 ;
        RECT 88.485 208.275 88.775 209.440 ;
        RECT 88.950 209.285 89.300 209.935 ;
        RECT 89.470 209.115 89.700 210.105 ;
        RECT 89.035 208.945 89.700 209.115 ;
        RECT 89.035 208.445 89.205 208.945 ;
        RECT 89.375 208.275 89.705 208.775 ;
        RECT 89.875 208.445 90.060 210.565 ;
        RECT 90.315 210.365 90.565 210.825 ;
        RECT 90.735 210.375 91.070 210.545 ;
        RECT 91.265 210.375 91.940 210.545 ;
        RECT 90.735 210.235 90.905 210.375 ;
        RECT 90.230 209.245 90.510 210.195 ;
        RECT 90.680 210.105 90.905 210.235 ;
        RECT 90.680 209.000 90.850 210.105 ;
        RECT 91.075 209.955 91.600 210.175 ;
        RECT 91.020 209.190 91.260 209.785 ;
        RECT 91.430 209.255 91.600 209.955 ;
        RECT 91.770 209.595 91.940 210.375 ;
        RECT 92.260 210.325 92.630 210.825 ;
        RECT 92.810 210.375 93.215 210.545 ;
        RECT 93.385 210.375 94.170 210.545 ;
        RECT 92.810 210.145 92.980 210.375 ;
        RECT 92.150 209.845 92.980 210.145 ;
        RECT 93.365 209.875 93.830 210.205 ;
        RECT 92.150 209.815 92.350 209.845 ;
        RECT 92.470 209.595 92.640 209.665 ;
        RECT 91.770 209.425 92.640 209.595 ;
        RECT 92.130 209.335 92.640 209.425 ;
        RECT 90.680 208.870 90.985 209.000 ;
        RECT 91.430 208.890 91.960 209.255 ;
        RECT 90.300 208.275 90.565 208.735 ;
        RECT 90.735 208.445 90.985 208.870 ;
        RECT 92.130 208.720 92.300 209.335 ;
        RECT 91.195 208.550 92.300 208.720 ;
        RECT 92.470 208.275 92.640 209.075 ;
        RECT 92.810 208.775 92.980 209.845 ;
        RECT 93.150 208.945 93.340 209.665 ;
        RECT 93.510 208.915 93.830 209.875 ;
        RECT 94.000 209.915 94.170 210.375 ;
        RECT 94.445 210.295 94.655 210.825 ;
        RECT 94.915 210.085 95.245 210.610 ;
        RECT 95.415 210.215 95.585 210.825 ;
        RECT 95.755 210.170 96.085 210.605 ;
        RECT 96.255 210.310 96.425 210.825 ;
        RECT 96.855 210.275 97.025 210.565 ;
        RECT 97.195 210.445 97.525 210.825 ;
        RECT 95.755 210.085 96.135 210.170 ;
        RECT 96.855 210.105 97.520 210.275 ;
        RECT 95.045 209.915 95.245 210.085 ;
        RECT 95.910 210.045 96.135 210.085 ;
        RECT 94.000 209.585 94.875 209.915 ;
        RECT 95.045 209.585 95.795 209.915 ;
        RECT 92.810 208.445 93.060 208.775 ;
        RECT 94.000 208.745 94.170 209.585 ;
        RECT 95.045 209.380 95.235 209.585 ;
        RECT 95.965 209.465 96.135 210.045 ;
        RECT 95.920 209.415 96.135 209.465 ;
        RECT 94.340 209.005 95.235 209.380 ;
        RECT 95.745 209.335 96.135 209.415 ;
        RECT 93.285 208.575 94.170 208.745 ;
        RECT 94.350 208.275 94.665 208.775 ;
        RECT 94.895 208.445 95.235 209.005 ;
        RECT 95.405 208.275 95.575 209.285 ;
        RECT 95.745 208.490 96.075 209.335 ;
        RECT 96.770 209.285 97.120 209.935 ;
        RECT 96.245 208.275 96.415 209.190 ;
        RECT 97.290 209.115 97.520 210.105 ;
        RECT 96.855 208.945 97.520 209.115 ;
        RECT 96.855 208.445 97.025 208.945 ;
        RECT 97.195 208.275 97.525 208.775 ;
        RECT 97.695 208.445 97.880 210.565 ;
        RECT 98.135 210.365 98.385 210.825 ;
        RECT 98.555 210.375 98.890 210.545 ;
        RECT 99.085 210.375 99.760 210.545 ;
        RECT 98.555 210.235 98.725 210.375 ;
        RECT 98.050 209.245 98.330 210.195 ;
        RECT 98.500 210.105 98.725 210.235 ;
        RECT 98.500 209.000 98.670 210.105 ;
        RECT 98.895 209.955 99.420 210.175 ;
        RECT 98.840 209.190 99.080 209.785 ;
        RECT 99.250 209.255 99.420 209.955 ;
        RECT 99.590 209.595 99.760 210.375 ;
        RECT 100.080 210.325 100.450 210.825 ;
        RECT 100.630 210.375 101.035 210.545 ;
        RECT 101.205 210.375 101.990 210.545 ;
        RECT 100.630 210.145 100.800 210.375 ;
        RECT 99.970 209.845 100.800 210.145 ;
        RECT 101.185 209.875 101.650 210.205 ;
        RECT 99.970 209.815 100.170 209.845 ;
        RECT 100.290 209.595 100.460 209.665 ;
        RECT 99.590 209.425 100.460 209.595 ;
        RECT 99.950 209.335 100.460 209.425 ;
        RECT 98.500 208.870 98.805 209.000 ;
        RECT 99.250 208.890 99.780 209.255 ;
        RECT 98.120 208.275 98.385 208.735 ;
        RECT 98.555 208.445 98.805 208.870 ;
        RECT 99.950 208.720 100.120 209.335 ;
        RECT 99.015 208.550 100.120 208.720 ;
        RECT 100.290 208.275 100.460 209.075 ;
        RECT 100.630 208.775 100.800 209.845 ;
        RECT 100.970 208.945 101.160 209.665 ;
        RECT 101.330 208.915 101.650 209.875 ;
        RECT 101.820 209.915 101.990 210.375 ;
        RECT 102.265 210.295 102.475 210.825 ;
        RECT 102.735 210.085 103.065 210.610 ;
        RECT 103.235 210.215 103.405 210.825 ;
        RECT 103.575 210.170 103.905 210.605 ;
        RECT 104.215 210.275 104.385 210.565 ;
        RECT 104.555 210.445 104.885 210.825 ;
        RECT 103.575 210.085 103.955 210.170 ;
        RECT 104.215 210.105 104.880 210.275 ;
        RECT 102.865 209.915 103.065 210.085 ;
        RECT 103.730 210.045 103.955 210.085 ;
        RECT 101.820 209.585 102.695 209.915 ;
        RECT 102.865 209.585 103.615 209.915 ;
        RECT 100.630 208.445 100.880 208.775 ;
        RECT 101.820 208.745 101.990 209.585 ;
        RECT 102.865 209.380 103.055 209.585 ;
        RECT 103.785 209.465 103.955 210.045 ;
        RECT 103.740 209.415 103.955 209.465 ;
        RECT 102.160 209.005 103.055 209.380 ;
        RECT 103.565 209.335 103.955 209.415 ;
        RECT 101.105 208.575 101.990 208.745 ;
        RECT 102.170 208.275 102.485 208.775 ;
        RECT 102.715 208.445 103.055 209.005 ;
        RECT 103.225 208.275 103.395 209.285 ;
        RECT 103.565 208.490 103.895 209.335 ;
        RECT 104.130 209.285 104.480 209.935 ;
        RECT 104.650 209.115 104.880 210.105 ;
        RECT 104.215 208.945 104.880 209.115 ;
        RECT 104.215 208.445 104.385 208.945 ;
        RECT 104.555 208.275 104.885 208.775 ;
        RECT 105.055 208.445 105.240 210.565 ;
        RECT 105.495 210.365 105.745 210.825 ;
        RECT 105.915 210.375 106.250 210.545 ;
        RECT 106.445 210.375 107.120 210.545 ;
        RECT 105.915 210.235 106.085 210.375 ;
        RECT 105.410 209.245 105.690 210.195 ;
        RECT 105.860 210.105 106.085 210.235 ;
        RECT 105.860 209.000 106.030 210.105 ;
        RECT 106.255 209.955 106.780 210.175 ;
        RECT 106.200 209.190 106.440 209.785 ;
        RECT 106.610 209.255 106.780 209.955 ;
        RECT 106.950 209.595 107.120 210.375 ;
        RECT 107.440 210.325 107.810 210.825 ;
        RECT 107.990 210.375 108.395 210.545 ;
        RECT 108.565 210.375 109.350 210.545 ;
        RECT 107.990 210.145 108.160 210.375 ;
        RECT 107.330 209.845 108.160 210.145 ;
        RECT 108.545 209.875 109.010 210.205 ;
        RECT 107.330 209.815 107.530 209.845 ;
        RECT 107.650 209.595 107.820 209.665 ;
        RECT 106.950 209.425 107.820 209.595 ;
        RECT 107.310 209.335 107.820 209.425 ;
        RECT 105.860 208.870 106.165 209.000 ;
        RECT 106.610 208.890 107.140 209.255 ;
        RECT 105.480 208.275 105.745 208.735 ;
        RECT 105.915 208.445 106.165 208.870 ;
        RECT 107.310 208.720 107.480 209.335 ;
        RECT 106.375 208.550 107.480 208.720 ;
        RECT 107.650 208.275 107.820 209.075 ;
        RECT 107.990 208.775 108.160 209.845 ;
        RECT 108.330 208.945 108.520 209.665 ;
        RECT 108.690 208.915 109.010 209.875 ;
        RECT 109.180 209.915 109.350 210.375 ;
        RECT 109.625 210.295 109.835 210.825 ;
        RECT 110.095 210.085 110.425 210.610 ;
        RECT 110.595 210.215 110.765 210.825 ;
        RECT 110.935 210.170 111.265 210.605 ;
        RECT 110.935 210.085 111.315 210.170 ;
        RECT 110.225 209.915 110.425 210.085 ;
        RECT 111.090 210.045 111.315 210.085 ;
        RECT 109.180 209.585 110.055 209.915 ;
        RECT 110.225 209.585 110.975 209.915 ;
        RECT 107.990 208.445 108.240 208.775 ;
        RECT 109.180 208.745 109.350 209.585 ;
        RECT 110.225 209.380 110.415 209.585 ;
        RECT 111.145 209.465 111.315 210.045 ;
        RECT 111.525 210.005 111.755 210.825 ;
        RECT 111.925 210.025 112.255 210.655 ;
        RECT 111.505 209.585 111.835 209.835 ;
        RECT 111.100 209.415 111.315 209.465 ;
        RECT 112.005 209.425 112.255 210.025 ;
        RECT 112.425 210.005 112.635 210.825 ;
        RECT 112.925 210.005 113.135 210.825 ;
        RECT 113.305 210.025 113.635 210.655 ;
        RECT 109.520 209.005 110.415 209.380 ;
        RECT 110.925 209.335 111.315 209.415 ;
        RECT 108.465 208.575 109.350 208.745 ;
        RECT 109.530 208.275 109.845 208.775 ;
        RECT 110.075 208.445 110.415 209.005 ;
        RECT 110.585 208.275 110.755 209.285 ;
        RECT 110.925 208.490 111.255 209.335 ;
        RECT 111.525 208.275 111.755 209.415 ;
        RECT 111.925 208.445 112.255 209.425 ;
        RECT 113.305 209.425 113.555 210.025 ;
        RECT 113.805 210.005 114.035 210.825 ;
        RECT 114.245 210.100 114.535 210.825 ;
        RECT 115.795 210.310 115.965 210.825 ;
        RECT 116.135 210.170 116.465 210.605 ;
        RECT 116.635 210.215 116.805 210.825 ;
        RECT 116.085 210.085 116.465 210.170 ;
        RECT 116.975 210.085 117.305 210.610 ;
        RECT 117.565 210.295 117.775 210.825 ;
        RECT 118.050 210.375 118.835 210.545 ;
        RECT 119.005 210.375 119.410 210.545 ;
        RECT 116.085 210.045 116.310 210.085 ;
        RECT 113.725 209.585 114.055 209.835 ;
        RECT 116.085 209.465 116.255 210.045 ;
        RECT 116.975 209.915 117.175 210.085 ;
        RECT 118.050 209.915 118.220 210.375 ;
        RECT 116.425 209.585 117.175 209.915 ;
        RECT 117.345 209.585 118.220 209.915 ;
        RECT 112.425 208.275 112.635 209.415 ;
        RECT 112.925 208.275 113.135 209.415 ;
        RECT 113.305 208.445 113.635 209.425 ;
        RECT 113.805 208.275 114.035 209.415 ;
        RECT 114.245 208.275 114.535 209.440 ;
        RECT 116.085 209.415 116.300 209.465 ;
        RECT 116.085 209.335 116.475 209.415 ;
        RECT 115.805 208.275 115.975 209.190 ;
        RECT 116.145 208.490 116.475 209.335 ;
        RECT 116.985 209.380 117.175 209.585 ;
        RECT 116.645 208.275 116.815 209.285 ;
        RECT 116.985 209.005 117.880 209.380 ;
        RECT 116.985 208.445 117.325 209.005 ;
        RECT 117.555 208.275 117.870 208.775 ;
        RECT 118.050 208.745 118.220 209.585 ;
        RECT 118.390 209.875 118.855 210.205 ;
        RECT 119.240 210.145 119.410 210.375 ;
        RECT 119.590 210.325 119.960 210.825 ;
        RECT 120.280 210.375 120.955 210.545 ;
        RECT 121.150 210.375 121.485 210.545 ;
        RECT 118.390 208.915 118.710 209.875 ;
        RECT 119.240 209.845 120.070 210.145 ;
        RECT 118.880 208.945 119.070 209.665 ;
        RECT 119.240 208.775 119.410 209.845 ;
        RECT 119.870 209.815 120.070 209.845 ;
        RECT 119.580 209.595 119.750 209.665 ;
        RECT 120.280 209.595 120.450 210.375 ;
        RECT 121.315 210.235 121.485 210.375 ;
        RECT 121.655 210.365 121.905 210.825 ;
        RECT 119.580 209.425 120.450 209.595 ;
        RECT 120.620 209.955 121.145 210.175 ;
        RECT 121.315 210.105 121.540 210.235 ;
        RECT 119.580 209.335 120.090 209.425 ;
        RECT 118.050 208.575 118.935 208.745 ;
        RECT 119.160 208.445 119.410 208.775 ;
        RECT 119.580 208.275 119.750 209.075 ;
        RECT 119.920 208.720 120.090 209.335 ;
        RECT 120.620 209.255 120.790 209.955 ;
        RECT 120.260 208.890 120.790 209.255 ;
        RECT 120.960 209.190 121.200 209.785 ;
        RECT 121.370 209.000 121.540 210.105 ;
        RECT 121.710 209.245 121.990 210.195 ;
        RECT 121.235 208.870 121.540 209.000 ;
        RECT 119.920 208.550 121.025 208.720 ;
        RECT 121.235 208.445 121.485 208.870 ;
        RECT 121.655 208.275 121.920 208.735 ;
        RECT 122.160 208.445 122.345 210.565 ;
        RECT 122.515 210.445 122.845 210.825 ;
        RECT 123.015 210.275 123.185 210.565 ;
        RECT 122.520 210.105 123.185 210.275 ;
        RECT 123.535 210.275 123.705 210.565 ;
        RECT 123.875 210.445 124.205 210.825 ;
        RECT 123.535 210.105 124.200 210.275 ;
        RECT 122.520 209.115 122.750 210.105 ;
        RECT 122.920 209.285 123.270 209.935 ;
        RECT 123.450 209.285 123.800 209.935 ;
        RECT 123.970 209.115 124.200 210.105 ;
        RECT 122.520 208.945 123.185 209.115 ;
        RECT 122.515 208.275 122.845 208.775 ;
        RECT 123.015 208.445 123.185 208.945 ;
        RECT 123.535 208.945 124.200 209.115 ;
        RECT 123.535 208.445 123.705 208.945 ;
        RECT 123.875 208.275 124.205 208.775 ;
        RECT 124.375 208.445 124.560 210.565 ;
        RECT 124.815 210.365 125.065 210.825 ;
        RECT 125.235 210.375 125.570 210.545 ;
        RECT 125.765 210.375 126.440 210.545 ;
        RECT 125.235 210.235 125.405 210.375 ;
        RECT 124.730 209.245 125.010 210.195 ;
        RECT 125.180 210.105 125.405 210.235 ;
        RECT 125.180 209.000 125.350 210.105 ;
        RECT 125.575 209.955 126.100 210.175 ;
        RECT 125.520 209.190 125.760 209.785 ;
        RECT 125.930 209.255 126.100 209.955 ;
        RECT 126.270 209.595 126.440 210.375 ;
        RECT 126.760 210.325 127.130 210.825 ;
        RECT 127.310 210.375 127.715 210.545 ;
        RECT 127.885 210.375 128.670 210.545 ;
        RECT 127.310 210.145 127.480 210.375 ;
        RECT 126.650 209.845 127.480 210.145 ;
        RECT 127.865 209.875 128.330 210.205 ;
        RECT 126.650 209.815 126.850 209.845 ;
        RECT 126.970 209.595 127.140 209.665 ;
        RECT 126.270 209.425 127.140 209.595 ;
        RECT 126.630 209.335 127.140 209.425 ;
        RECT 125.180 208.870 125.485 209.000 ;
        RECT 125.930 208.890 126.460 209.255 ;
        RECT 124.800 208.275 125.065 208.735 ;
        RECT 125.235 208.445 125.485 208.870 ;
        RECT 126.630 208.720 126.800 209.335 ;
        RECT 125.695 208.550 126.800 208.720 ;
        RECT 126.970 208.275 127.140 209.075 ;
        RECT 127.310 208.775 127.480 209.845 ;
        RECT 127.650 208.945 127.840 209.665 ;
        RECT 128.010 208.915 128.330 209.875 ;
        RECT 128.500 209.915 128.670 210.375 ;
        RECT 128.945 210.295 129.155 210.825 ;
        RECT 129.415 210.085 129.745 210.610 ;
        RECT 129.915 210.215 130.085 210.825 ;
        RECT 130.255 210.170 130.585 210.605 ;
        RECT 130.805 210.280 136.150 210.825 ;
        RECT 130.255 210.085 130.635 210.170 ;
        RECT 129.545 209.915 129.745 210.085 ;
        RECT 130.410 210.045 130.635 210.085 ;
        RECT 128.500 209.585 129.375 209.915 ;
        RECT 129.545 209.585 130.295 209.915 ;
        RECT 127.310 208.445 127.560 208.775 ;
        RECT 128.500 208.745 128.670 209.585 ;
        RECT 129.545 209.380 129.735 209.585 ;
        RECT 130.465 209.465 130.635 210.045 ;
        RECT 130.420 209.415 130.635 209.465 ;
        RECT 132.390 209.450 132.730 210.280 ;
        RECT 136.325 210.055 139.835 210.825 ;
        RECT 140.005 210.100 140.295 210.825 ;
        RECT 140.465 210.280 145.810 210.825 ;
        RECT 128.840 209.005 129.735 209.380 ;
        RECT 130.245 209.335 130.635 209.415 ;
        RECT 127.785 208.575 128.670 208.745 ;
        RECT 128.850 208.275 129.165 208.775 ;
        RECT 129.395 208.445 129.735 209.005 ;
        RECT 129.905 208.275 130.075 209.285 ;
        RECT 130.245 208.490 130.575 209.335 ;
        RECT 134.210 208.710 134.560 209.960 ;
        RECT 136.325 209.535 137.975 210.055 ;
        RECT 138.145 209.365 139.835 209.885 ;
        RECT 142.050 209.450 142.390 210.280 ;
        RECT 145.985 210.055 148.575 210.825 ;
        RECT 149.205 210.075 150.415 210.825 ;
        RECT 130.805 208.275 136.150 208.710 ;
        RECT 136.325 208.275 139.835 209.365 ;
        RECT 140.005 208.275 140.295 209.440 ;
        RECT 143.870 208.710 144.220 209.960 ;
        RECT 145.985 209.535 147.195 210.055 ;
        RECT 147.365 209.365 148.575 209.885 ;
        RECT 140.465 208.275 145.810 208.710 ;
        RECT 145.985 208.275 148.575 209.365 ;
        RECT 149.205 209.365 149.725 209.905 ;
        RECT 149.895 209.535 150.415 210.075 ;
        RECT 149.205 208.275 150.415 209.365 ;
        RECT 11.120 208.105 150.500 208.275 ;
        RECT 11.205 207.015 12.415 208.105 ;
        RECT 12.585 207.670 17.930 208.105 ;
        RECT 11.205 206.305 11.725 206.845 ;
        RECT 11.895 206.475 12.415 207.015 ;
        RECT 11.205 205.555 12.415 206.305 ;
        RECT 14.170 206.100 14.510 206.930 ;
        RECT 15.990 206.420 16.340 207.670 ;
        RECT 18.105 207.015 21.615 208.105 ;
        RECT 18.105 206.325 19.755 206.845 ;
        RECT 19.925 206.495 21.615 207.015 ;
        RECT 22.245 207.030 22.515 207.935 ;
        RECT 22.685 207.345 23.015 208.105 ;
        RECT 23.195 207.175 23.365 207.935 ;
        RECT 12.585 205.555 17.930 206.100 ;
        RECT 18.105 205.555 21.615 206.325 ;
        RECT 22.245 206.230 22.415 207.030 ;
        RECT 22.700 207.005 23.365 207.175 ;
        RECT 22.700 206.860 22.870 207.005 ;
        RECT 24.085 206.940 24.375 208.105 ;
        RECT 24.545 207.235 24.820 207.935 ;
        RECT 25.030 207.560 25.245 208.105 ;
        RECT 25.415 207.595 25.890 207.935 ;
        RECT 26.060 207.600 26.675 208.105 ;
        RECT 26.060 207.425 26.255 207.600 ;
        RECT 22.585 206.530 22.870 206.860 ;
        RECT 22.700 206.275 22.870 206.530 ;
        RECT 23.105 206.455 23.435 206.825 ;
        RECT 22.245 205.725 22.505 206.230 ;
        RECT 22.700 206.105 23.365 206.275 ;
        RECT 22.685 205.555 23.015 205.935 ;
        RECT 23.195 205.725 23.365 206.105 ;
        RECT 24.085 205.555 24.375 206.280 ;
        RECT 24.545 206.205 24.715 207.235 ;
        RECT 24.990 207.065 25.705 207.360 ;
        RECT 25.925 207.235 26.255 207.425 ;
        RECT 26.425 207.065 26.675 207.430 ;
        RECT 24.885 206.895 26.675 207.065 ;
        RECT 24.885 206.465 25.115 206.895 ;
        RECT 24.545 205.725 24.805 206.205 ;
        RECT 25.285 206.195 25.695 206.715 ;
        RECT 24.975 205.555 25.305 206.015 ;
        RECT 25.495 205.775 25.695 206.195 ;
        RECT 25.865 206.040 26.120 206.895 ;
        RECT 26.915 206.715 27.085 207.935 ;
        RECT 27.335 207.595 27.595 208.105 ;
        RECT 26.290 206.465 27.085 206.715 ;
        RECT 27.255 206.545 27.595 207.425 ;
        RECT 26.835 206.375 27.085 206.465 ;
        RECT 25.865 205.775 26.655 206.040 ;
        RECT 26.835 205.955 27.165 206.375 ;
        RECT 27.335 205.555 27.595 206.375 ;
        RECT 27.775 205.735 28.035 207.925 ;
        RECT 28.205 207.375 28.545 208.105 ;
        RECT 28.725 207.195 28.995 207.925 ;
        RECT 28.225 206.975 28.995 207.195 ;
        RECT 29.175 207.215 29.405 207.925 ;
        RECT 29.575 207.395 29.905 208.105 ;
        RECT 30.075 207.215 30.335 207.925 ;
        RECT 29.175 206.975 30.335 207.215 ;
        RECT 30.525 207.015 32.195 208.105 ;
        RECT 32.545 207.190 32.715 208.105 ;
        RECT 32.885 207.045 33.215 207.890 ;
        RECT 33.385 207.095 33.555 208.105 ;
        RECT 33.725 207.375 34.065 207.935 ;
        RECT 34.295 207.605 34.610 208.105 ;
        RECT 34.790 207.635 35.675 207.805 ;
        RECT 28.225 206.305 28.515 206.975 ;
        RECT 28.695 206.485 29.160 206.795 ;
        RECT 29.340 206.485 29.865 206.795 ;
        RECT 28.225 206.105 29.455 206.305 ;
        RECT 28.295 205.555 28.965 205.925 ;
        RECT 29.145 205.735 29.455 206.105 ;
        RECT 29.635 205.845 29.865 206.485 ;
        RECT 30.045 206.465 30.345 206.795 ;
        RECT 30.525 206.325 31.275 206.845 ;
        RECT 31.445 206.495 32.195 207.015 ;
        RECT 32.825 206.965 33.215 207.045 ;
        RECT 33.725 207.000 34.620 207.375 ;
        RECT 32.825 206.915 33.040 206.965 ;
        RECT 32.825 206.335 32.995 206.915 ;
        RECT 33.725 206.795 33.915 207.000 ;
        RECT 34.790 206.795 34.960 207.635 ;
        RECT 35.900 207.605 36.150 207.935 ;
        RECT 33.165 206.465 33.915 206.795 ;
        RECT 34.085 206.465 34.960 206.795 ;
        RECT 30.045 205.555 30.335 206.285 ;
        RECT 30.525 205.555 32.195 206.325 ;
        RECT 32.825 206.295 33.050 206.335 ;
        RECT 33.715 206.295 33.915 206.465 ;
        RECT 32.825 206.210 33.205 206.295 ;
        RECT 32.535 205.555 32.705 206.070 ;
        RECT 32.875 205.775 33.205 206.210 ;
        RECT 33.375 205.555 33.545 206.165 ;
        RECT 33.715 205.770 34.045 206.295 ;
        RECT 34.305 205.555 34.515 206.085 ;
        RECT 34.790 206.005 34.960 206.465 ;
        RECT 35.130 206.505 35.450 207.465 ;
        RECT 35.620 206.715 35.810 207.435 ;
        RECT 35.980 206.535 36.150 207.605 ;
        RECT 36.320 207.305 36.490 208.105 ;
        RECT 36.660 207.660 37.765 207.830 ;
        RECT 36.660 207.045 36.830 207.660 ;
        RECT 37.975 207.510 38.225 207.935 ;
        RECT 38.395 207.645 38.660 208.105 ;
        RECT 37.000 207.125 37.530 207.490 ;
        RECT 37.975 207.380 38.280 207.510 ;
        RECT 36.320 206.955 36.830 207.045 ;
        RECT 36.320 206.785 37.190 206.955 ;
        RECT 36.320 206.715 36.490 206.785 ;
        RECT 36.610 206.535 36.810 206.565 ;
        RECT 35.130 206.175 35.595 206.505 ;
        RECT 35.980 206.235 36.810 206.535 ;
        RECT 35.980 206.005 36.150 206.235 ;
        RECT 34.790 205.835 35.575 206.005 ;
        RECT 35.745 205.835 36.150 206.005 ;
        RECT 36.330 205.555 36.700 206.055 ;
        RECT 37.020 206.005 37.190 206.785 ;
        RECT 37.360 206.425 37.530 207.125 ;
        RECT 37.700 206.595 37.940 207.190 ;
        RECT 37.360 206.205 37.885 206.425 ;
        RECT 38.110 206.275 38.280 207.380 ;
        RECT 38.055 206.145 38.280 206.275 ;
        RECT 38.450 206.185 38.730 207.135 ;
        RECT 38.055 206.005 38.225 206.145 ;
        RECT 37.020 205.835 37.695 206.005 ;
        RECT 37.890 205.835 38.225 206.005 ;
        RECT 38.395 205.555 38.645 206.015 ;
        RECT 38.900 205.815 39.085 207.935 ;
        RECT 39.255 207.605 39.585 208.105 ;
        RECT 39.755 207.435 39.925 207.935 ;
        RECT 39.260 207.265 39.925 207.435 ;
        RECT 39.260 206.275 39.490 207.265 ;
        RECT 39.660 206.445 40.010 207.095 ;
        RECT 40.185 207.015 43.695 208.105 ;
        RECT 43.865 207.015 45.075 208.105 ;
        RECT 45.335 207.485 45.505 207.915 ;
        RECT 45.675 207.655 46.005 208.105 ;
        RECT 45.335 207.255 46.010 207.485 ;
        RECT 40.185 206.325 41.835 206.845 ;
        RECT 42.005 206.495 43.695 207.015 ;
        RECT 39.260 206.105 39.925 206.275 ;
        RECT 39.255 205.555 39.585 205.935 ;
        RECT 39.755 205.815 39.925 206.105 ;
        RECT 40.185 205.555 43.695 206.325 ;
        RECT 43.865 206.305 44.385 206.845 ;
        RECT 44.555 206.475 45.075 207.015 ;
        RECT 43.865 205.555 45.075 206.305 ;
        RECT 45.305 206.235 45.605 207.085 ;
        RECT 45.775 206.605 46.010 207.255 ;
        RECT 46.180 206.945 46.465 207.890 ;
        RECT 46.645 207.635 47.330 208.105 ;
        RECT 46.640 207.115 47.335 207.425 ;
        RECT 47.510 207.050 47.815 207.835 ;
        RECT 46.180 206.795 47.040 206.945 ;
        RECT 46.180 206.775 47.465 206.795 ;
        RECT 45.775 206.275 46.310 206.605 ;
        RECT 46.480 206.415 47.465 206.775 ;
        RECT 45.775 206.125 45.995 206.275 ;
        RECT 45.250 205.555 45.585 206.060 ;
        RECT 45.755 205.750 45.995 206.125 ;
        RECT 46.480 206.080 46.650 206.415 ;
        RECT 47.640 206.245 47.815 207.050 ;
        RECT 48.005 207.015 49.675 208.105 ;
        RECT 46.275 205.885 46.650 206.080 ;
        RECT 46.275 205.740 46.445 205.885 ;
        RECT 47.010 205.555 47.405 206.050 ;
        RECT 47.575 205.725 47.815 206.245 ;
        RECT 48.005 206.325 48.755 206.845 ;
        RECT 48.925 206.495 49.675 207.015 ;
        RECT 49.845 206.940 50.135 208.105 ;
        RECT 50.305 207.015 51.975 208.105 ;
        RECT 50.305 206.325 51.055 206.845 ;
        RECT 51.225 206.495 51.975 207.015 ;
        RECT 52.235 207.175 52.405 207.935 ;
        RECT 52.620 207.345 52.950 208.105 ;
        RECT 52.235 207.005 52.950 207.175 ;
        RECT 53.120 207.030 53.375 207.935 ;
        RECT 52.145 206.455 52.500 206.825 ;
        RECT 52.780 206.795 52.950 207.005 ;
        RECT 52.780 206.465 53.035 206.795 ;
        RECT 48.005 205.555 49.675 206.325 ;
        RECT 49.845 205.555 50.135 206.280 ;
        RECT 50.305 205.555 51.975 206.325 ;
        RECT 52.780 206.275 52.950 206.465 ;
        RECT 53.205 206.300 53.375 207.030 ;
        RECT 53.550 206.955 53.810 208.105 ;
        RECT 53.985 207.670 59.330 208.105 ;
        RECT 52.235 206.105 52.950 206.275 ;
        RECT 52.235 205.725 52.405 206.105 ;
        RECT 52.620 205.555 52.950 205.935 ;
        RECT 53.120 205.725 53.375 206.300 ;
        RECT 53.550 205.555 53.810 206.395 ;
        RECT 55.570 206.100 55.910 206.930 ;
        RECT 57.390 206.420 57.740 207.670 ;
        RECT 59.505 207.015 63.015 208.105 ;
        RECT 63.185 207.015 64.395 208.105 ;
        RECT 59.505 206.325 61.155 206.845 ;
        RECT 61.325 206.495 63.015 207.015 ;
        RECT 53.985 205.555 59.330 206.100 ;
        RECT 59.505 205.555 63.015 206.325 ;
        RECT 63.185 206.305 63.705 206.845 ;
        RECT 63.875 206.475 64.395 207.015 ;
        RECT 64.570 206.965 64.825 208.105 ;
        RECT 65.020 207.555 66.215 207.885 ;
        RECT 65.075 206.795 65.245 207.355 ;
        RECT 65.470 207.135 65.890 207.385 ;
        RECT 66.395 207.305 66.675 208.105 ;
        RECT 65.470 206.965 66.715 207.135 ;
        RECT 66.885 206.965 67.155 207.935 ;
        RECT 67.330 207.725 67.665 208.105 ;
        RECT 66.545 206.795 66.715 206.965 ;
        RECT 66.925 206.915 67.155 206.965 ;
        RECT 64.570 206.545 64.905 206.795 ;
        RECT 65.075 206.465 65.815 206.795 ;
        RECT 66.545 206.465 66.775 206.795 ;
        RECT 65.075 206.375 65.325 206.465 ;
        RECT 63.185 205.555 64.395 206.305 ;
        RECT 64.590 206.205 65.325 206.375 ;
        RECT 66.545 206.295 66.715 206.465 ;
        RECT 64.590 205.735 64.900 206.205 ;
        RECT 65.975 206.125 66.715 206.295 ;
        RECT 66.985 206.230 67.155 206.915 ;
        RECT 67.325 206.235 67.565 207.545 ;
        RECT 67.835 207.135 68.085 207.935 ;
        RECT 68.305 207.385 68.635 208.105 ;
        RECT 68.820 207.135 69.070 207.935 ;
        RECT 69.535 207.305 69.865 208.105 ;
        RECT 70.035 207.675 70.375 207.935 ;
        RECT 67.735 206.965 69.925 207.135 ;
        RECT 65.070 205.555 65.805 206.035 ;
        RECT 65.975 205.775 66.145 206.125 ;
        RECT 66.315 205.555 66.695 205.955 ;
        RECT 66.885 205.885 67.155 206.230 ;
        RECT 67.735 206.055 67.905 206.965 ;
        RECT 69.610 206.795 69.925 206.965 ;
        RECT 67.410 205.725 67.905 206.055 ;
        RECT 68.125 205.830 68.475 206.795 ;
        RECT 68.655 205.825 68.955 206.795 ;
        RECT 69.135 205.825 69.415 206.795 ;
        RECT 69.610 206.545 69.940 206.795 ;
        RECT 69.595 205.555 69.865 206.355 ;
        RECT 70.115 206.275 70.375 207.675 ;
        RECT 70.750 207.135 71.080 207.935 ;
        RECT 71.250 207.305 71.580 208.105 ;
        RECT 71.880 207.135 72.210 207.935 ;
        RECT 72.855 207.305 73.105 208.105 ;
        RECT 70.750 206.965 73.185 207.135 ;
        RECT 73.375 206.965 73.545 208.105 ;
        RECT 73.715 206.965 74.055 207.935 ;
        RECT 74.225 207.015 75.435 208.105 ;
        RECT 70.545 206.545 70.895 206.795 ;
        RECT 71.080 206.335 71.250 206.965 ;
        RECT 71.420 206.545 71.750 206.745 ;
        RECT 71.920 206.545 72.250 206.745 ;
        RECT 72.420 206.545 72.840 206.745 ;
        RECT 73.015 206.715 73.185 206.965 ;
        RECT 73.015 206.545 73.710 206.715 ;
        RECT 70.035 205.765 70.375 206.275 ;
        RECT 70.750 205.725 71.250 206.335 ;
        RECT 71.880 206.205 73.105 206.375 ;
        RECT 73.880 206.355 74.055 206.965 ;
        RECT 71.880 205.725 72.210 206.205 ;
        RECT 72.380 205.555 72.605 206.015 ;
        RECT 72.775 205.725 73.105 206.205 ;
        RECT 73.295 205.555 73.545 206.355 ;
        RECT 73.715 205.725 74.055 206.355 ;
        RECT 74.225 206.305 74.745 206.845 ;
        RECT 74.915 206.475 75.435 207.015 ;
        RECT 75.605 206.940 75.895 208.105 ;
        RECT 76.065 207.670 81.410 208.105 ;
        RECT 74.225 205.555 75.435 206.305 ;
        RECT 75.605 205.555 75.895 206.280 ;
        RECT 77.650 206.100 77.990 206.930 ;
        RECT 79.470 206.420 79.820 207.670 ;
        RECT 81.770 207.135 82.160 207.310 ;
        RECT 82.645 207.305 82.975 208.105 ;
        RECT 83.145 207.315 83.680 207.935 ;
        RECT 81.770 206.965 83.195 207.135 ;
        RECT 81.645 206.235 82.000 206.795 ;
        RECT 76.065 205.555 81.410 206.100 ;
        RECT 82.170 206.065 82.340 206.965 ;
        RECT 82.510 206.235 82.775 206.795 ;
        RECT 83.025 206.465 83.195 206.965 ;
        RECT 83.365 206.295 83.680 207.315 ;
        RECT 83.895 206.965 84.225 208.105 ;
        RECT 84.755 207.135 85.085 207.920 ;
        RECT 85.355 207.435 85.525 207.935 ;
        RECT 85.695 207.605 86.025 208.105 ;
        RECT 85.355 207.265 86.020 207.435 ;
        RECT 84.405 206.965 85.085 207.135 ;
        RECT 83.885 206.545 84.235 206.795 ;
        RECT 84.405 206.365 84.575 206.965 ;
        RECT 84.745 206.545 85.095 206.795 ;
        RECT 85.270 206.445 85.620 207.095 ;
        RECT 81.750 205.555 81.990 206.065 ;
        RECT 82.170 205.735 82.450 206.065 ;
        RECT 82.680 205.555 82.895 206.065 ;
        RECT 83.065 205.725 83.680 206.295 ;
        RECT 83.895 205.555 84.165 206.365 ;
        RECT 84.335 205.725 84.665 206.365 ;
        RECT 84.835 205.555 85.075 206.365 ;
        RECT 85.790 206.275 86.020 207.265 ;
        RECT 85.355 206.105 86.020 206.275 ;
        RECT 85.355 205.815 85.525 206.105 ;
        RECT 85.695 205.555 86.025 205.935 ;
        RECT 86.195 205.815 86.380 207.935 ;
        RECT 86.620 207.645 86.885 208.105 ;
        RECT 87.055 207.510 87.305 207.935 ;
        RECT 87.515 207.660 88.620 207.830 ;
        RECT 87.000 207.380 87.305 207.510 ;
        RECT 86.550 206.185 86.830 207.135 ;
        RECT 87.000 206.275 87.170 207.380 ;
        RECT 87.340 206.595 87.580 207.190 ;
        RECT 87.750 207.125 88.280 207.490 ;
        RECT 87.750 206.425 87.920 207.125 ;
        RECT 88.450 207.045 88.620 207.660 ;
        RECT 88.790 207.305 88.960 208.105 ;
        RECT 89.130 207.605 89.380 207.935 ;
        RECT 89.605 207.635 90.490 207.805 ;
        RECT 88.450 206.955 88.960 207.045 ;
        RECT 87.000 206.145 87.225 206.275 ;
        RECT 87.395 206.205 87.920 206.425 ;
        RECT 88.090 206.785 88.960 206.955 ;
        RECT 86.635 205.555 86.885 206.015 ;
        RECT 87.055 206.005 87.225 206.145 ;
        RECT 88.090 206.005 88.260 206.785 ;
        RECT 88.790 206.715 88.960 206.785 ;
        RECT 88.470 206.535 88.670 206.565 ;
        RECT 89.130 206.535 89.300 207.605 ;
        RECT 89.470 206.715 89.660 207.435 ;
        RECT 88.470 206.235 89.300 206.535 ;
        RECT 89.830 206.505 90.150 207.465 ;
        RECT 87.055 205.835 87.390 206.005 ;
        RECT 87.585 205.835 88.260 206.005 ;
        RECT 88.580 205.555 88.950 206.055 ;
        RECT 89.130 206.005 89.300 206.235 ;
        RECT 89.685 206.175 90.150 206.505 ;
        RECT 90.320 206.795 90.490 207.635 ;
        RECT 90.670 207.605 90.985 208.105 ;
        RECT 91.215 207.375 91.555 207.935 ;
        RECT 90.660 207.000 91.555 207.375 ;
        RECT 91.725 207.095 91.895 208.105 ;
        RECT 91.365 206.795 91.555 207.000 ;
        RECT 92.065 207.045 92.395 207.890 ;
        RECT 92.565 207.190 92.735 208.105 ;
        RECT 92.065 206.965 92.455 207.045 ;
        RECT 92.240 206.915 92.455 206.965 ;
        RECT 90.320 206.465 91.195 206.795 ;
        RECT 91.365 206.465 92.115 206.795 ;
        RECT 90.320 206.005 90.490 206.465 ;
        RECT 91.365 206.295 91.565 206.465 ;
        RECT 92.285 206.335 92.455 206.915 ;
        RECT 92.230 206.295 92.455 206.335 ;
        RECT 89.130 205.835 89.535 206.005 ;
        RECT 89.705 205.835 90.490 206.005 ;
        RECT 90.765 205.555 90.975 206.085 ;
        RECT 91.235 205.770 91.565 206.295 ;
        RECT 92.075 206.210 92.455 206.295 ;
        RECT 93.085 206.965 93.470 207.935 ;
        RECT 93.640 207.645 93.965 208.105 ;
        RECT 94.485 207.475 94.765 207.935 ;
        RECT 93.640 207.255 94.765 207.475 ;
        RECT 93.085 206.295 93.365 206.965 ;
        RECT 93.640 206.795 94.090 207.255 ;
        RECT 94.955 207.085 95.355 207.935 ;
        RECT 95.755 207.645 96.025 208.105 ;
        RECT 96.195 207.475 96.480 207.935 ;
        RECT 93.535 206.465 94.090 206.795 ;
        RECT 94.260 206.525 95.355 207.085 ;
        RECT 93.640 206.355 94.090 206.465 ;
        RECT 91.735 205.555 91.905 206.165 ;
        RECT 92.075 205.775 92.405 206.210 ;
        RECT 92.575 205.555 92.745 206.070 ;
        RECT 93.085 205.725 93.470 206.295 ;
        RECT 93.640 206.185 94.765 206.355 ;
        RECT 93.640 205.555 93.965 206.015 ;
        RECT 94.485 205.725 94.765 206.185 ;
        RECT 94.955 205.725 95.355 206.525 ;
        RECT 95.525 207.255 96.480 207.475 ;
        RECT 95.525 206.355 95.735 207.255 ;
        RECT 97.775 207.175 97.945 207.935 ;
        RECT 98.160 207.345 98.490 208.105 ;
        RECT 95.905 206.525 96.595 207.085 ;
        RECT 97.775 207.005 98.490 207.175 ;
        RECT 98.660 207.030 98.915 207.935 ;
        RECT 97.685 206.455 98.040 206.825 ;
        RECT 98.320 206.795 98.490 207.005 ;
        RECT 98.320 206.465 98.575 206.795 ;
        RECT 95.525 206.185 96.480 206.355 ;
        RECT 98.320 206.275 98.490 206.465 ;
        RECT 98.745 206.300 98.915 207.030 ;
        RECT 99.090 206.955 99.350 208.105 ;
        RECT 99.565 206.965 99.795 208.105 ;
        RECT 99.965 206.955 100.295 207.935 ;
        RECT 100.465 206.965 100.675 208.105 ;
        RECT 99.545 206.545 99.875 206.795 ;
        RECT 95.755 205.555 96.025 206.015 ;
        RECT 96.195 205.725 96.480 206.185 ;
        RECT 97.775 206.105 98.490 206.275 ;
        RECT 97.775 205.725 97.945 206.105 ;
        RECT 98.160 205.555 98.490 205.935 ;
        RECT 98.660 205.725 98.915 206.300 ;
        RECT 99.090 205.555 99.350 206.395 ;
        RECT 99.565 205.555 99.795 206.375 ;
        RECT 100.045 206.355 100.295 206.955 ;
        RECT 101.365 206.940 101.655 208.105 ;
        RECT 101.825 207.015 103.495 208.105 ;
        RECT 103.755 207.435 103.925 207.935 ;
        RECT 104.095 207.605 104.425 208.105 ;
        RECT 103.755 207.265 104.420 207.435 ;
        RECT 99.965 205.725 100.295 206.355 ;
        RECT 100.465 205.555 100.675 206.375 ;
        RECT 101.825 206.325 102.575 206.845 ;
        RECT 102.745 206.495 103.495 207.015 ;
        RECT 103.670 206.445 104.020 207.095 ;
        RECT 101.365 205.555 101.655 206.280 ;
        RECT 101.825 205.555 103.495 206.325 ;
        RECT 104.190 206.275 104.420 207.265 ;
        RECT 103.755 206.105 104.420 206.275 ;
        RECT 103.755 205.815 103.925 206.105 ;
        RECT 104.095 205.555 104.425 205.935 ;
        RECT 104.595 205.815 104.780 207.935 ;
        RECT 105.020 207.645 105.285 208.105 ;
        RECT 105.455 207.510 105.705 207.935 ;
        RECT 105.915 207.660 107.020 207.830 ;
        RECT 105.400 207.380 105.705 207.510 ;
        RECT 104.950 206.185 105.230 207.135 ;
        RECT 105.400 206.275 105.570 207.380 ;
        RECT 105.740 206.595 105.980 207.190 ;
        RECT 106.150 207.125 106.680 207.490 ;
        RECT 106.150 206.425 106.320 207.125 ;
        RECT 106.850 207.045 107.020 207.660 ;
        RECT 107.190 207.305 107.360 208.105 ;
        RECT 107.530 207.605 107.780 207.935 ;
        RECT 108.005 207.635 108.890 207.805 ;
        RECT 106.850 206.955 107.360 207.045 ;
        RECT 105.400 206.145 105.625 206.275 ;
        RECT 105.795 206.205 106.320 206.425 ;
        RECT 106.490 206.785 107.360 206.955 ;
        RECT 105.035 205.555 105.285 206.015 ;
        RECT 105.455 206.005 105.625 206.145 ;
        RECT 106.490 206.005 106.660 206.785 ;
        RECT 107.190 206.715 107.360 206.785 ;
        RECT 106.870 206.535 107.070 206.565 ;
        RECT 107.530 206.535 107.700 207.605 ;
        RECT 107.870 206.715 108.060 207.435 ;
        RECT 106.870 206.235 107.700 206.535 ;
        RECT 108.230 206.505 108.550 207.465 ;
        RECT 105.455 205.835 105.790 206.005 ;
        RECT 105.985 205.835 106.660 206.005 ;
        RECT 106.980 205.555 107.350 206.055 ;
        RECT 107.530 206.005 107.700 206.235 ;
        RECT 108.085 206.175 108.550 206.505 ;
        RECT 108.720 206.795 108.890 207.635 ;
        RECT 109.070 207.605 109.385 208.105 ;
        RECT 109.615 207.375 109.955 207.935 ;
        RECT 109.060 207.000 109.955 207.375 ;
        RECT 110.125 207.095 110.295 208.105 ;
        RECT 109.765 206.795 109.955 207.000 ;
        RECT 110.465 207.045 110.795 207.890 ;
        RECT 111.575 207.435 111.745 207.935 ;
        RECT 111.915 207.605 112.245 208.105 ;
        RECT 111.575 207.265 112.240 207.435 ;
        RECT 110.465 206.965 110.855 207.045 ;
        RECT 110.640 206.915 110.855 206.965 ;
        RECT 108.720 206.465 109.595 206.795 ;
        RECT 109.765 206.465 110.515 206.795 ;
        RECT 108.720 206.005 108.890 206.465 ;
        RECT 109.765 206.295 109.965 206.465 ;
        RECT 110.685 206.335 110.855 206.915 ;
        RECT 111.490 206.445 111.840 207.095 ;
        RECT 110.630 206.295 110.855 206.335 ;
        RECT 107.530 205.835 107.935 206.005 ;
        RECT 108.105 205.835 108.890 206.005 ;
        RECT 109.165 205.555 109.375 206.085 ;
        RECT 109.635 205.770 109.965 206.295 ;
        RECT 110.475 206.210 110.855 206.295 ;
        RECT 112.010 206.275 112.240 207.265 ;
        RECT 110.135 205.555 110.305 206.165 ;
        RECT 110.475 205.775 110.805 206.210 ;
        RECT 111.575 206.105 112.240 206.275 ;
        RECT 111.575 205.815 111.745 206.105 ;
        RECT 111.915 205.555 112.245 205.935 ;
        RECT 112.415 205.815 112.600 207.935 ;
        RECT 112.840 207.645 113.105 208.105 ;
        RECT 113.275 207.510 113.525 207.935 ;
        RECT 113.735 207.660 114.840 207.830 ;
        RECT 113.220 207.380 113.525 207.510 ;
        RECT 112.770 206.185 113.050 207.135 ;
        RECT 113.220 206.275 113.390 207.380 ;
        RECT 113.560 206.595 113.800 207.190 ;
        RECT 113.970 207.125 114.500 207.490 ;
        RECT 113.970 206.425 114.140 207.125 ;
        RECT 114.670 207.045 114.840 207.660 ;
        RECT 115.010 207.305 115.180 208.105 ;
        RECT 115.350 207.605 115.600 207.935 ;
        RECT 115.825 207.635 116.710 207.805 ;
        RECT 114.670 206.955 115.180 207.045 ;
        RECT 113.220 206.145 113.445 206.275 ;
        RECT 113.615 206.205 114.140 206.425 ;
        RECT 114.310 206.785 115.180 206.955 ;
        RECT 112.855 205.555 113.105 206.015 ;
        RECT 113.275 206.005 113.445 206.145 ;
        RECT 114.310 206.005 114.480 206.785 ;
        RECT 115.010 206.715 115.180 206.785 ;
        RECT 114.690 206.535 114.890 206.565 ;
        RECT 115.350 206.535 115.520 207.605 ;
        RECT 115.690 206.715 115.880 207.435 ;
        RECT 114.690 206.235 115.520 206.535 ;
        RECT 116.050 206.505 116.370 207.465 ;
        RECT 113.275 205.835 113.610 206.005 ;
        RECT 113.805 205.835 114.480 206.005 ;
        RECT 114.800 205.555 115.170 206.055 ;
        RECT 115.350 206.005 115.520 206.235 ;
        RECT 115.905 206.175 116.370 206.505 ;
        RECT 116.540 206.795 116.710 207.635 ;
        RECT 116.890 207.605 117.205 208.105 ;
        RECT 117.435 207.375 117.775 207.935 ;
        RECT 116.880 207.000 117.775 207.375 ;
        RECT 117.945 207.095 118.115 208.105 ;
        RECT 117.585 206.795 117.775 207.000 ;
        RECT 118.285 207.045 118.615 207.890 ;
        RECT 118.285 206.965 118.675 207.045 ;
        RECT 118.845 207.015 120.055 208.105 ;
        RECT 120.340 207.475 120.625 207.935 ;
        RECT 120.795 207.645 121.065 208.105 ;
        RECT 120.340 207.255 121.295 207.475 ;
        RECT 118.460 206.915 118.675 206.965 ;
        RECT 116.540 206.465 117.415 206.795 ;
        RECT 117.585 206.465 118.335 206.795 ;
        RECT 116.540 206.005 116.710 206.465 ;
        RECT 117.585 206.295 117.785 206.465 ;
        RECT 118.505 206.335 118.675 206.915 ;
        RECT 118.450 206.295 118.675 206.335 ;
        RECT 115.350 205.835 115.755 206.005 ;
        RECT 115.925 205.835 116.710 206.005 ;
        RECT 116.985 205.555 117.195 206.085 ;
        RECT 117.455 205.770 117.785 206.295 ;
        RECT 118.295 206.210 118.675 206.295 ;
        RECT 118.845 206.305 119.365 206.845 ;
        RECT 119.535 206.475 120.055 207.015 ;
        RECT 120.225 206.525 120.915 207.085 ;
        RECT 121.085 206.355 121.295 207.255 ;
        RECT 117.955 205.555 118.125 206.165 ;
        RECT 118.295 205.775 118.625 206.210 ;
        RECT 118.845 205.555 120.055 206.305 ;
        RECT 120.340 206.185 121.295 206.355 ;
        RECT 121.465 207.085 121.865 207.935 ;
        RECT 122.055 207.475 122.335 207.935 ;
        RECT 122.855 207.645 123.180 208.105 ;
        RECT 122.055 207.255 123.180 207.475 ;
        RECT 121.465 206.525 122.560 207.085 ;
        RECT 122.730 206.795 123.180 207.255 ;
        RECT 123.350 206.965 123.735 207.935 ;
        RECT 123.965 206.965 124.175 208.105 ;
        RECT 120.340 205.725 120.625 206.185 ;
        RECT 120.795 205.555 121.065 206.015 ;
        RECT 121.465 205.725 121.865 206.525 ;
        RECT 122.730 206.465 123.285 206.795 ;
        RECT 122.730 206.355 123.180 206.465 ;
        RECT 122.055 206.185 123.180 206.355 ;
        RECT 123.455 206.295 123.735 206.965 ;
        RECT 124.345 206.955 124.675 207.935 ;
        RECT 124.845 206.965 125.075 208.105 ;
        RECT 125.285 207.015 126.955 208.105 ;
        RECT 122.055 205.725 122.335 206.185 ;
        RECT 122.855 205.555 123.180 206.015 ;
        RECT 123.350 205.725 123.735 206.295 ;
        RECT 123.965 205.555 124.175 206.375 ;
        RECT 124.345 206.355 124.595 206.955 ;
        RECT 124.765 206.545 125.095 206.795 ;
        RECT 124.345 205.725 124.675 206.355 ;
        RECT 124.845 205.555 125.075 206.375 ;
        RECT 125.285 206.325 126.035 206.845 ;
        RECT 126.205 206.495 126.955 207.015 ;
        RECT 127.125 206.940 127.415 208.105 ;
        RECT 127.585 207.015 129.255 208.105 ;
        RECT 127.585 206.325 128.335 206.845 ;
        RECT 128.505 206.495 129.255 207.015 ;
        RECT 129.885 206.965 130.270 207.935 ;
        RECT 130.440 207.645 130.765 208.105 ;
        RECT 131.285 207.475 131.565 207.935 ;
        RECT 130.440 207.255 131.565 207.475 ;
        RECT 125.285 205.555 126.955 206.325 ;
        RECT 127.125 205.555 127.415 206.280 ;
        RECT 127.585 205.555 129.255 206.325 ;
        RECT 129.885 206.295 130.165 206.965 ;
        RECT 130.440 206.795 130.890 207.255 ;
        RECT 131.755 207.085 132.155 207.935 ;
        RECT 132.555 207.645 132.825 208.105 ;
        RECT 132.995 207.475 133.280 207.935 ;
        RECT 133.565 207.670 138.910 208.105 ;
        RECT 139.085 207.670 144.430 208.105 ;
        RECT 130.335 206.465 130.890 206.795 ;
        RECT 131.060 206.525 132.155 207.085 ;
        RECT 130.440 206.355 130.890 206.465 ;
        RECT 129.885 205.725 130.270 206.295 ;
        RECT 130.440 206.185 131.565 206.355 ;
        RECT 130.440 205.555 130.765 206.015 ;
        RECT 131.285 205.725 131.565 206.185 ;
        RECT 131.755 205.725 132.155 206.525 ;
        RECT 132.325 207.255 133.280 207.475 ;
        RECT 132.325 206.355 132.535 207.255 ;
        RECT 132.705 206.525 133.395 207.085 ;
        RECT 132.325 206.185 133.280 206.355 ;
        RECT 132.555 205.555 132.825 206.015 ;
        RECT 132.995 205.725 133.280 206.185 ;
        RECT 135.150 206.100 135.490 206.930 ;
        RECT 136.970 206.420 137.320 207.670 ;
        RECT 140.670 206.100 141.010 206.930 ;
        RECT 142.490 206.420 142.840 207.670 ;
        RECT 144.605 207.015 148.115 208.105 ;
        RECT 144.605 206.325 146.255 206.845 ;
        RECT 146.425 206.495 148.115 207.015 ;
        RECT 149.205 207.015 150.415 208.105 ;
        RECT 149.205 206.475 149.725 207.015 ;
        RECT 133.565 205.555 138.910 206.100 ;
        RECT 139.085 205.555 144.430 206.100 ;
        RECT 144.605 205.555 148.115 206.325 ;
        RECT 149.895 206.305 150.415 206.845 ;
        RECT 149.205 205.555 150.415 206.305 ;
        RECT 11.120 205.385 150.500 205.555 ;
        RECT 11.205 204.635 12.415 205.385 ;
        RECT 12.585 204.840 17.930 205.385 ;
        RECT 18.105 204.840 23.450 205.385 ;
        RECT 23.625 204.840 28.970 205.385 ;
        RECT 30.065 205.005 30.955 205.175 ;
        RECT 11.205 204.095 11.725 204.635 ;
        RECT 11.895 203.925 12.415 204.465 ;
        RECT 14.170 204.010 14.510 204.840 ;
        RECT 11.205 202.835 12.415 203.925 ;
        RECT 15.990 203.270 16.340 204.520 ;
        RECT 19.690 204.010 20.030 204.840 ;
        RECT 21.510 203.270 21.860 204.520 ;
        RECT 25.210 204.010 25.550 204.840 ;
        RECT 27.030 203.270 27.380 204.520 ;
        RECT 30.065 204.450 30.615 204.835 ;
        RECT 30.785 204.280 30.955 205.005 ;
        RECT 30.065 204.210 30.955 204.280 ;
        RECT 31.125 204.680 31.345 205.165 ;
        RECT 31.515 204.845 31.765 205.385 ;
        RECT 31.935 204.735 32.195 205.215 ;
        RECT 31.125 204.255 31.455 204.680 ;
        RECT 30.065 204.185 30.960 204.210 ;
        RECT 30.065 204.170 30.970 204.185 ;
        RECT 30.065 204.155 30.975 204.170 ;
        RECT 30.065 204.150 30.985 204.155 ;
        RECT 30.065 204.140 30.990 204.150 ;
        RECT 30.065 204.130 30.995 204.140 ;
        RECT 30.065 204.125 31.005 204.130 ;
        RECT 30.065 204.115 31.015 204.125 ;
        RECT 30.065 204.110 31.025 204.115 ;
        RECT 30.065 203.660 30.325 204.110 ;
        RECT 30.690 204.105 31.025 204.110 ;
        RECT 30.690 204.100 31.040 204.105 ;
        RECT 30.690 204.090 31.055 204.100 ;
        RECT 30.690 204.085 31.080 204.090 ;
        RECT 31.625 204.085 31.855 204.480 ;
        RECT 30.690 204.080 31.855 204.085 ;
        RECT 30.720 204.045 31.855 204.080 ;
        RECT 30.755 204.020 31.855 204.045 ;
        RECT 30.785 203.990 31.855 204.020 ;
        RECT 30.805 203.960 31.855 203.990 ;
        RECT 30.825 203.930 31.855 203.960 ;
        RECT 30.895 203.920 31.855 203.930 ;
        RECT 30.920 203.910 31.855 203.920 ;
        RECT 30.940 203.895 31.855 203.910 ;
        RECT 30.960 203.880 31.855 203.895 ;
        RECT 30.965 203.870 31.750 203.880 ;
        RECT 30.980 203.835 31.750 203.870 ;
        RECT 30.495 203.515 30.825 203.760 ;
        RECT 30.995 203.585 31.750 203.835 ;
        RECT 32.025 203.705 32.195 204.735 ;
        RECT 32.365 204.615 35.875 205.385 ;
        RECT 36.965 204.660 37.255 205.385 ;
        RECT 37.425 204.635 38.635 205.385 ;
        RECT 38.825 204.695 39.065 205.215 ;
        RECT 39.235 204.890 39.630 205.385 ;
        RECT 40.195 205.055 40.365 205.200 ;
        RECT 39.990 204.860 40.365 205.055 ;
        RECT 32.365 204.095 34.015 204.615 ;
        RECT 34.185 203.925 35.875 204.445 ;
        RECT 37.425 204.095 37.945 204.635 ;
        RECT 30.495 203.490 30.680 203.515 ;
        RECT 30.065 203.390 30.680 203.490 ;
        RECT 12.585 202.835 17.930 203.270 ;
        RECT 18.105 202.835 23.450 203.270 ;
        RECT 23.625 202.835 28.970 203.270 ;
        RECT 30.065 202.835 30.670 203.390 ;
        RECT 30.845 203.005 31.325 203.345 ;
        RECT 31.495 202.835 31.750 203.380 ;
        RECT 31.920 203.005 32.195 203.705 ;
        RECT 32.365 202.835 35.875 203.925 ;
        RECT 36.965 202.835 37.255 204.000 ;
        RECT 38.115 203.925 38.635 204.465 ;
        RECT 37.425 202.835 38.635 203.925 ;
        RECT 38.825 203.890 39.000 204.695 ;
        RECT 39.990 204.525 40.160 204.860 ;
        RECT 40.645 204.815 40.885 205.190 ;
        RECT 41.055 204.880 41.390 205.385 ;
        RECT 40.645 204.665 40.865 204.815 ;
        RECT 39.175 204.165 40.160 204.525 ;
        RECT 40.330 204.335 40.865 204.665 ;
        RECT 39.175 204.145 40.460 204.165 ;
        RECT 39.600 203.995 40.460 204.145 ;
        RECT 38.825 203.105 39.130 203.890 ;
        RECT 39.305 203.515 40.000 203.825 ;
        RECT 39.310 202.835 39.995 203.305 ;
        RECT 40.175 203.050 40.460 203.995 ;
        RECT 40.630 203.685 40.865 204.335 ;
        RECT 41.035 203.855 41.335 204.705 ;
        RECT 41.565 204.615 44.155 205.385 ;
        RECT 41.565 204.095 42.775 204.615 ;
        RECT 44.805 204.575 45.045 205.385 ;
        RECT 45.215 204.575 45.545 205.215 ;
        RECT 45.715 204.575 45.985 205.385 ;
        RECT 46.190 204.995 46.520 205.385 ;
        RECT 46.690 204.825 46.915 205.205 ;
        RECT 42.945 203.925 44.155 204.445 ;
        RECT 44.785 204.145 45.135 204.395 ;
        RECT 45.305 203.975 45.475 204.575 ;
        RECT 45.645 204.145 45.995 204.395 ;
        RECT 46.175 204.145 46.415 204.795 ;
        RECT 46.585 204.645 46.915 204.825 ;
        RECT 46.585 203.975 46.760 204.645 ;
        RECT 47.115 204.475 47.345 205.095 ;
        RECT 47.525 204.655 47.825 205.385 ;
        RECT 48.005 204.585 48.315 205.385 ;
        RECT 48.520 204.585 49.215 205.215 ;
        RECT 49.385 204.615 52.895 205.385 ;
        RECT 53.985 204.645 54.450 205.190 ;
        RECT 46.930 204.145 47.345 204.475 ;
        RECT 47.525 204.145 47.820 204.475 ;
        RECT 48.015 204.145 48.350 204.415 ;
        RECT 48.520 203.985 48.690 204.585 ;
        RECT 48.860 204.145 49.195 204.395 ;
        RECT 49.385 204.095 51.035 204.615 ;
        RECT 40.630 203.455 41.305 203.685 ;
        RECT 40.635 202.835 40.965 203.285 ;
        RECT 41.135 203.025 41.305 203.455 ;
        RECT 41.565 202.835 44.155 203.925 ;
        RECT 44.795 203.805 45.475 203.975 ;
        RECT 44.795 203.020 45.125 203.805 ;
        RECT 45.655 202.835 45.985 203.975 ;
        RECT 46.175 203.785 46.760 203.975 ;
        RECT 46.175 203.015 46.450 203.785 ;
        RECT 46.930 203.615 47.825 203.945 ;
        RECT 46.620 203.445 47.825 203.615 ;
        RECT 46.620 203.015 46.950 203.445 ;
        RECT 47.120 202.835 47.315 203.275 ;
        RECT 47.495 203.015 47.825 203.445 ;
        RECT 48.005 202.835 48.285 203.975 ;
        RECT 48.455 203.005 48.785 203.985 ;
        RECT 48.955 202.835 49.215 203.975 ;
        RECT 51.205 203.925 52.895 204.445 ;
        RECT 49.385 202.835 52.895 203.925 ;
        RECT 53.985 203.685 54.155 204.645 ;
        RECT 54.955 204.565 55.125 205.385 ;
        RECT 55.295 204.735 55.625 205.215 ;
        RECT 55.795 204.995 56.145 205.385 ;
        RECT 56.315 204.815 56.545 205.215 ;
        RECT 56.035 204.735 56.545 204.815 ;
        RECT 55.295 204.645 56.545 204.735 ;
        RECT 56.715 204.645 57.035 205.125 ;
        RECT 55.295 204.565 56.205 204.645 ;
        RECT 54.325 204.025 54.570 204.475 ;
        RECT 54.830 204.195 55.525 204.395 ;
        RECT 55.695 204.225 56.295 204.395 ;
        RECT 55.695 204.025 55.865 204.225 ;
        RECT 56.525 204.055 56.695 204.475 ;
        RECT 54.325 203.855 55.865 204.025 ;
        RECT 56.035 203.885 56.695 204.055 ;
        RECT 56.035 203.685 56.205 203.885 ;
        RECT 56.865 203.715 57.035 204.645 ;
        RECT 53.985 203.515 56.205 203.685 ;
        RECT 56.375 203.515 57.035 203.715 ;
        RECT 57.665 204.645 58.130 205.190 ;
        RECT 57.665 203.685 57.835 204.645 ;
        RECT 58.635 204.565 58.805 205.385 ;
        RECT 58.975 204.735 59.305 205.215 ;
        RECT 59.475 204.995 59.825 205.385 ;
        RECT 59.995 204.815 60.225 205.215 ;
        RECT 59.715 204.735 60.225 204.815 ;
        RECT 58.975 204.645 60.225 204.735 ;
        RECT 60.395 204.645 60.715 205.125 ;
        RECT 58.975 204.565 59.885 204.645 ;
        RECT 58.005 204.025 58.250 204.475 ;
        RECT 58.510 204.195 59.205 204.395 ;
        RECT 59.375 204.225 59.975 204.395 ;
        RECT 59.375 204.025 59.545 204.225 ;
        RECT 60.205 204.055 60.375 204.475 ;
        RECT 58.005 203.855 59.545 204.025 ;
        RECT 59.715 203.885 60.375 204.055 ;
        RECT 59.715 203.685 59.885 203.885 ;
        RECT 60.545 203.715 60.715 204.645 ;
        RECT 60.885 204.615 62.555 205.385 ;
        RECT 62.725 204.660 63.015 205.385 ;
        RECT 63.185 204.840 68.530 205.385 ;
        RECT 60.885 204.095 61.635 204.615 ;
        RECT 61.805 203.925 62.555 204.445 ;
        RECT 64.770 204.010 65.110 204.840 ;
        RECT 69.250 204.735 69.425 205.215 ;
        RECT 69.595 204.905 69.925 205.385 ;
        RECT 70.145 204.965 71.660 205.215 ;
        RECT 71.830 204.985 72.160 205.385 ;
        RECT 70.145 204.735 70.315 204.965 ;
        RECT 71.460 204.815 71.660 204.965 ;
        RECT 69.250 204.565 70.315 204.735 ;
        RECT 57.665 203.515 59.885 203.685 ;
        RECT 60.055 203.515 60.715 203.715 ;
        RECT 53.985 202.835 54.285 203.345 ;
        RECT 54.455 203.005 54.785 203.515 ;
        RECT 56.375 203.345 56.545 203.515 ;
        RECT 54.955 202.835 55.585 203.345 ;
        RECT 56.165 203.175 56.545 203.345 ;
        RECT 56.715 202.835 57.015 203.345 ;
        RECT 57.665 202.835 57.965 203.345 ;
        RECT 58.135 203.005 58.465 203.515 ;
        RECT 60.055 203.345 60.225 203.515 ;
        RECT 58.635 202.835 59.265 203.345 ;
        RECT 59.845 203.175 60.225 203.345 ;
        RECT 60.395 202.835 60.695 203.345 ;
        RECT 60.885 202.835 62.555 203.925 ;
        RECT 62.725 202.835 63.015 204.000 ;
        RECT 66.590 203.270 66.940 204.520 ;
        RECT 70.495 204.395 70.775 204.795 ;
        RECT 69.165 204.185 69.515 204.395 ;
        RECT 69.695 204.365 70.135 204.395 ;
        RECT 69.685 204.195 70.135 204.365 ;
        RECT 69.695 204.185 70.135 204.195 ;
        RECT 70.305 204.185 70.775 204.395 ;
        RECT 71.025 204.395 71.280 204.795 ;
        RECT 71.460 204.645 72.215 204.815 ;
        RECT 71.025 204.185 71.355 204.395 ;
        RECT 71.550 204.365 71.835 204.475 ;
        RECT 71.525 204.195 71.835 204.365 ;
        RECT 71.550 204.145 71.835 204.195 ;
        RECT 72.005 204.025 72.215 204.645 ;
        RECT 72.385 204.615 75.895 205.385 ;
        RECT 76.065 204.635 77.275 205.385 ;
        RECT 77.445 205.005 78.335 205.175 ;
        RECT 72.385 204.095 74.035 204.615 ;
        RECT 69.255 203.975 71.380 204.015 ;
        RECT 71.985 203.975 72.215 204.025 ;
        RECT 69.255 203.845 72.215 203.975 ;
        RECT 74.205 203.925 75.895 204.445 ;
        RECT 76.065 204.095 76.585 204.635 ;
        RECT 76.755 203.925 77.275 204.465 ;
        RECT 77.445 204.450 77.995 204.835 ;
        RECT 78.165 204.280 78.335 205.005 ;
        RECT 63.185 202.835 68.530 203.270 ;
        RECT 69.255 203.005 69.425 203.845 ;
        RECT 71.230 203.805 72.215 203.845 ;
        RECT 69.595 203.175 69.845 203.675 ;
        RECT 70.095 203.635 71.105 203.675 ;
        RECT 70.095 203.425 71.705 203.635 ;
        RECT 70.095 203.345 70.320 203.425 ;
        RECT 70.435 203.175 70.765 203.215 ;
        RECT 69.595 203.005 70.765 203.175 ;
        RECT 70.955 202.835 71.285 203.255 ;
        RECT 71.455 203.005 71.705 203.425 ;
        RECT 71.875 202.835 72.205 203.595 ;
        RECT 72.385 202.835 75.895 203.925 ;
        RECT 76.065 202.835 77.275 203.925 ;
        RECT 77.445 204.210 78.335 204.280 ;
        RECT 78.505 204.680 78.725 205.165 ;
        RECT 78.895 204.845 79.145 205.385 ;
        RECT 79.315 204.735 79.575 205.215 ;
        RECT 78.505 204.255 78.835 204.680 ;
        RECT 77.445 204.185 78.340 204.210 ;
        RECT 77.445 204.170 78.350 204.185 ;
        RECT 77.445 204.155 78.355 204.170 ;
        RECT 77.445 204.150 78.365 204.155 ;
        RECT 77.445 204.140 78.370 204.150 ;
        RECT 77.445 204.130 78.375 204.140 ;
        RECT 77.445 204.125 78.385 204.130 ;
        RECT 77.445 204.115 78.395 204.125 ;
        RECT 77.445 204.110 78.405 204.115 ;
        RECT 77.445 203.660 77.705 204.110 ;
        RECT 78.070 204.105 78.405 204.110 ;
        RECT 78.070 204.100 78.420 204.105 ;
        RECT 78.070 204.090 78.435 204.100 ;
        RECT 78.070 204.085 78.460 204.090 ;
        RECT 79.005 204.085 79.235 204.480 ;
        RECT 78.070 204.080 79.235 204.085 ;
        RECT 78.100 204.045 79.235 204.080 ;
        RECT 78.135 204.020 79.235 204.045 ;
        RECT 78.165 203.990 79.235 204.020 ;
        RECT 78.185 203.960 79.235 203.990 ;
        RECT 78.205 203.930 79.235 203.960 ;
        RECT 78.275 203.920 79.235 203.930 ;
        RECT 78.300 203.910 79.235 203.920 ;
        RECT 78.320 203.895 79.235 203.910 ;
        RECT 78.340 203.880 79.235 203.895 ;
        RECT 78.345 203.870 79.130 203.880 ;
        RECT 78.360 203.835 79.130 203.870 ;
        RECT 77.875 203.515 78.205 203.760 ;
        RECT 78.375 203.585 79.130 203.835 ;
        RECT 79.405 203.705 79.575 204.735 ;
        RECT 80.405 204.755 80.735 205.115 ;
        RECT 81.355 204.925 81.605 205.385 ;
        RECT 81.775 204.925 82.335 205.215 ;
        RECT 82.595 205.045 82.765 205.080 ;
        RECT 80.405 204.565 81.795 204.755 ;
        RECT 81.625 204.475 81.795 204.565 ;
        RECT 80.220 204.145 80.895 204.395 ;
        RECT 81.115 204.145 81.455 204.395 ;
        RECT 81.625 204.145 81.915 204.475 ;
        RECT 80.220 203.785 80.485 204.145 ;
        RECT 81.625 203.895 81.795 204.145 ;
        RECT 77.875 203.490 78.060 203.515 ;
        RECT 77.445 203.390 78.060 203.490 ;
        RECT 77.445 202.835 78.050 203.390 ;
        RECT 78.225 203.005 78.705 203.345 ;
        RECT 78.875 202.835 79.130 203.380 ;
        RECT 79.300 203.005 79.575 203.705 ;
        RECT 80.855 203.725 81.795 203.895 ;
        RECT 80.405 202.835 80.685 203.505 ;
        RECT 80.855 203.175 81.155 203.725 ;
        RECT 82.085 203.555 82.335 204.925 ;
        RECT 82.565 204.875 82.765 205.045 ;
        RECT 82.595 204.515 82.765 204.875 ;
        RECT 82.955 204.855 83.185 205.160 ;
        RECT 83.355 205.025 83.685 205.385 ;
        RECT 83.880 204.855 84.170 205.205 ;
        RECT 82.955 204.685 84.170 204.855 ;
        RECT 84.345 204.615 87.855 205.385 ;
        RECT 88.485 204.660 88.775 205.385 ;
        RECT 88.945 204.615 90.615 205.385 ;
        RECT 90.875 204.835 91.045 205.125 ;
        RECT 91.215 205.005 91.545 205.385 ;
        RECT 90.875 204.665 91.540 204.835 ;
        RECT 82.595 204.345 83.115 204.515 ;
        RECT 82.510 203.815 82.755 204.175 ;
        RECT 82.945 203.965 83.115 204.345 ;
        RECT 83.285 204.145 83.670 204.475 ;
        RECT 83.850 204.365 84.110 204.475 ;
        RECT 83.850 204.195 84.115 204.365 ;
        RECT 83.850 204.145 84.110 204.195 ;
        RECT 82.945 203.685 83.295 203.965 ;
        RECT 81.355 202.835 81.685 203.555 ;
        RECT 81.875 203.005 82.335 203.555 ;
        RECT 82.510 202.835 82.765 203.635 ;
        RECT 82.965 203.005 83.295 203.685 ;
        RECT 83.475 203.095 83.670 204.145 ;
        RECT 84.345 204.095 85.995 204.615 ;
        RECT 83.850 202.835 84.170 203.975 ;
        RECT 86.165 203.925 87.855 204.445 ;
        RECT 88.945 204.095 89.695 204.615 ;
        RECT 84.345 202.835 87.855 203.925 ;
        RECT 88.485 202.835 88.775 204.000 ;
        RECT 89.865 203.925 90.615 204.445 ;
        RECT 88.945 202.835 90.615 203.925 ;
        RECT 90.790 203.845 91.140 204.495 ;
        RECT 91.310 203.675 91.540 204.665 ;
        RECT 90.875 203.505 91.540 203.675 ;
        RECT 90.875 203.005 91.045 203.505 ;
        RECT 91.215 202.835 91.545 203.335 ;
        RECT 91.715 203.005 91.900 205.125 ;
        RECT 92.155 204.925 92.405 205.385 ;
        RECT 92.575 204.935 92.910 205.105 ;
        RECT 93.105 204.935 93.780 205.105 ;
        RECT 92.575 204.795 92.745 204.935 ;
        RECT 92.070 203.805 92.350 204.755 ;
        RECT 92.520 204.665 92.745 204.795 ;
        RECT 92.520 203.560 92.690 204.665 ;
        RECT 92.915 204.515 93.440 204.735 ;
        RECT 92.860 203.750 93.100 204.345 ;
        RECT 93.270 203.815 93.440 204.515 ;
        RECT 93.610 204.155 93.780 204.935 ;
        RECT 94.100 204.885 94.470 205.385 ;
        RECT 94.650 204.935 95.055 205.105 ;
        RECT 95.225 204.935 96.010 205.105 ;
        RECT 94.650 204.705 94.820 204.935 ;
        RECT 93.990 204.405 94.820 204.705 ;
        RECT 95.205 204.435 95.670 204.765 ;
        RECT 93.990 204.375 94.190 204.405 ;
        RECT 94.310 204.155 94.480 204.225 ;
        RECT 93.610 203.985 94.480 204.155 ;
        RECT 93.970 203.895 94.480 203.985 ;
        RECT 92.520 203.430 92.825 203.560 ;
        RECT 93.270 203.450 93.800 203.815 ;
        RECT 92.140 202.835 92.405 203.295 ;
        RECT 92.575 203.005 92.825 203.430 ;
        RECT 93.970 203.280 94.140 203.895 ;
        RECT 93.035 203.110 94.140 203.280 ;
        RECT 94.310 202.835 94.480 203.635 ;
        RECT 94.650 203.335 94.820 204.405 ;
        RECT 94.990 203.505 95.180 204.225 ;
        RECT 95.350 203.475 95.670 204.435 ;
        RECT 95.840 204.475 96.010 204.935 ;
        RECT 96.285 204.855 96.495 205.385 ;
        RECT 96.755 204.645 97.085 205.170 ;
        RECT 97.255 204.775 97.425 205.385 ;
        RECT 97.595 204.730 97.925 205.165 ;
        RECT 98.095 204.870 98.265 205.385 ;
        RECT 98.605 204.840 103.950 205.385 ;
        RECT 97.595 204.645 97.975 204.730 ;
        RECT 96.885 204.475 97.085 204.645 ;
        RECT 97.750 204.605 97.975 204.645 ;
        RECT 95.840 204.145 96.715 204.475 ;
        RECT 96.885 204.145 97.635 204.475 ;
        RECT 94.650 203.005 94.900 203.335 ;
        RECT 95.840 203.305 96.010 204.145 ;
        RECT 96.885 203.940 97.075 204.145 ;
        RECT 97.805 204.025 97.975 204.605 ;
        RECT 97.760 203.975 97.975 204.025 ;
        RECT 100.190 204.010 100.530 204.840 ;
        RECT 104.125 204.615 106.715 205.385 ;
        RECT 106.935 204.730 107.265 205.165 ;
        RECT 107.435 204.775 107.605 205.385 ;
        RECT 106.885 204.645 107.265 204.730 ;
        RECT 107.775 204.645 108.105 205.170 ;
        RECT 108.365 204.855 108.575 205.385 ;
        RECT 108.850 204.935 109.635 205.105 ;
        RECT 109.805 204.935 110.210 205.105 ;
        RECT 96.180 203.565 97.075 203.940 ;
        RECT 97.585 203.895 97.975 203.975 ;
        RECT 95.125 203.135 96.010 203.305 ;
        RECT 96.190 202.835 96.505 203.335 ;
        RECT 96.735 203.005 97.075 203.565 ;
        RECT 97.245 202.835 97.415 203.845 ;
        RECT 97.585 203.050 97.915 203.895 ;
        RECT 98.085 202.835 98.255 203.750 ;
        RECT 102.010 203.270 102.360 204.520 ;
        RECT 104.125 204.095 105.335 204.615 ;
        RECT 106.885 204.605 107.110 204.645 ;
        RECT 105.505 203.925 106.715 204.445 ;
        RECT 98.605 202.835 103.950 203.270 ;
        RECT 104.125 202.835 106.715 203.925 ;
        RECT 106.885 204.025 107.055 204.605 ;
        RECT 107.775 204.475 107.975 204.645 ;
        RECT 108.850 204.475 109.020 204.935 ;
        RECT 107.225 204.145 107.975 204.475 ;
        RECT 108.145 204.145 109.020 204.475 ;
        RECT 106.885 203.975 107.100 204.025 ;
        RECT 106.885 203.895 107.275 203.975 ;
        RECT 106.945 203.050 107.275 203.895 ;
        RECT 107.785 203.940 107.975 204.145 ;
        RECT 107.445 202.835 107.615 203.845 ;
        RECT 107.785 203.565 108.680 203.940 ;
        RECT 107.785 203.005 108.125 203.565 ;
        RECT 108.355 202.835 108.670 203.335 ;
        RECT 108.850 203.305 109.020 204.145 ;
        RECT 109.190 204.435 109.655 204.765 ;
        RECT 110.040 204.705 110.210 204.935 ;
        RECT 110.390 204.885 110.760 205.385 ;
        RECT 111.080 204.935 111.755 205.105 ;
        RECT 111.950 204.935 112.285 205.105 ;
        RECT 109.190 203.475 109.510 204.435 ;
        RECT 110.040 204.405 110.870 204.705 ;
        RECT 109.680 203.505 109.870 204.225 ;
        RECT 110.040 203.335 110.210 204.405 ;
        RECT 110.670 204.375 110.870 204.405 ;
        RECT 110.380 204.155 110.550 204.225 ;
        RECT 111.080 204.155 111.250 204.935 ;
        RECT 112.115 204.795 112.285 204.935 ;
        RECT 112.455 204.925 112.705 205.385 ;
        RECT 110.380 203.985 111.250 204.155 ;
        RECT 111.420 204.515 111.945 204.735 ;
        RECT 112.115 204.665 112.340 204.795 ;
        RECT 110.380 203.895 110.890 203.985 ;
        RECT 108.850 203.135 109.735 203.305 ;
        RECT 109.960 203.005 110.210 203.335 ;
        RECT 110.380 202.835 110.550 203.635 ;
        RECT 110.720 203.280 110.890 203.895 ;
        RECT 111.420 203.815 111.590 204.515 ;
        RECT 111.060 203.450 111.590 203.815 ;
        RECT 111.760 203.750 112.000 204.345 ;
        RECT 112.170 203.560 112.340 204.665 ;
        RECT 112.510 203.805 112.790 204.755 ;
        RECT 112.035 203.430 112.340 203.560 ;
        RECT 110.720 203.110 111.825 203.280 ;
        RECT 112.035 203.005 112.285 203.430 ;
        RECT 112.455 202.835 112.720 203.295 ;
        RECT 112.960 203.005 113.145 205.125 ;
        RECT 113.315 205.005 113.645 205.385 ;
        RECT 113.815 204.835 113.985 205.125 ;
        RECT 113.320 204.665 113.985 204.835 ;
        RECT 113.320 203.675 113.550 204.665 ;
        RECT 114.245 204.660 114.535 205.385 ;
        RECT 114.705 204.840 120.050 205.385 ;
        RECT 120.225 204.840 125.570 205.385 ;
        RECT 125.745 204.840 131.090 205.385 ;
        RECT 131.265 204.840 136.610 205.385 ;
        RECT 113.720 203.845 114.070 204.495 ;
        RECT 116.290 204.010 116.630 204.840 ;
        RECT 113.320 203.505 113.985 203.675 ;
        RECT 113.315 202.835 113.645 203.335 ;
        RECT 113.815 203.005 113.985 203.505 ;
        RECT 114.245 202.835 114.535 204.000 ;
        RECT 118.110 203.270 118.460 204.520 ;
        RECT 121.810 204.010 122.150 204.840 ;
        RECT 123.630 203.270 123.980 204.520 ;
        RECT 127.330 204.010 127.670 204.840 ;
        RECT 129.150 203.270 129.500 204.520 ;
        RECT 132.850 204.010 133.190 204.840 ;
        RECT 136.785 204.615 139.375 205.385 ;
        RECT 140.005 204.660 140.295 205.385 ;
        RECT 140.465 204.840 145.810 205.385 ;
        RECT 134.670 203.270 135.020 204.520 ;
        RECT 136.785 204.095 137.995 204.615 ;
        RECT 138.165 203.925 139.375 204.445 ;
        RECT 142.050 204.010 142.390 204.840 ;
        RECT 145.985 204.615 148.575 205.385 ;
        RECT 149.205 204.635 150.415 205.385 ;
        RECT 114.705 202.835 120.050 203.270 ;
        RECT 120.225 202.835 125.570 203.270 ;
        RECT 125.745 202.835 131.090 203.270 ;
        RECT 131.265 202.835 136.610 203.270 ;
        RECT 136.785 202.835 139.375 203.925 ;
        RECT 140.005 202.835 140.295 204.000 ;
        RECT 143.870 203.270 144.220 204.520 ;
        RECT 145.985 204.095 147.195 204.615 ;
        RECT 147.365 203.925 148.575 204.445 ;
        RECT 140.465 202.835 145.810 203.270 ;
        RECT 145.985 202.835 148.575 203.925 ;
        RECT 149.205 203.925 149.725 204.465 ;
        RECT 149.895 204.095 150.415 204.635 ;
        RECT 149.205 202.835 150.415 203.925 ;
        RECT 11.120 202.665 150.500 202.835 ;
        RECT 11.205 201.575 12.415 202.665 ;
        RECT 12.585 201.575 16.095 202.665 ;
        RECT 16.815 201.995 16.985 202.495 ;
        RECT 17.155 202.165 17.485 202.665 ;
        RECT 16.815 201.825 17.480 201.995 ;
        RECT 11.205 200.865 11.725 201.405 ;
        RECT 11.895 201.035 12.415 201.575 ;
        RECT 12.585 200.885 14.235 201.405 ;
        RECT 14.405 201.055 16.095 201.575 ;
        RECT 16.730 201.005 17.080 201.655 ;
        RECT 11.205 200.115 12.415 200.865 ;
        RECT 12.585 200.115 16.095 200.885 ;
        RECT 17.250 200.835 17.480 201.825 ;
        RECT 16.815 200.665 17.480 200.835 ;
        RECT 16.815 200.375 16.985 200.665 ;
        RECT 17.155 200.115 17.485 200.495 ;
        RECT 17.655 200.375 17.840 202.495 ;
        RECT 18.080 202.205 18.345 202.665 ;
        RECT 18.515 202.070 18.765 202.495 ;
        RECT 18.975 202.220 20.080 202.390 ;
        RECT 18.460 201.940 18.765 202.070 ;
        RECT 18.010 200.745 18.290 201.695 ;
        RECT 18.460 200.835 18.630 201.940 ;
        RECT 18.800 201.155 19.040 201.750 ;
        RECT 19.210 201.685 19.740 202.050 ;
        RECT 19.210 200.985 19.380 201.685 ;
        RECT 19.910 201.605 20.080 202.220 ;
        RECT 20.250 201.865 20.420 202.665 ;
        RECT 20.590 202.165 20.840 202.495 ;
        RECT 21.065 202.195 21.950 202.365 ;
        RECT 19.910 201.515 20.420 201.605 ;
        RECT 18.460 200.705 18.685 200.835 ;
        RECT 18.855 200.765 19.380 200.985 ;
        RECT 19.550 201.345 20.420 201.515 ;
        RECT 18.095 200.115 18.345 200.575 ;
        RECT 18.515 200.565 18.685 200.705 ;
        RECT 19.550 200.565 19.720 201.345 ;
        RECT 20.250 201.275 20.420 201.345 ;
        RECT 19.930 201.095 20.130 201.125 ;
        RECT 20.590 201.095 20.760 202.165 ;
        RECT 20.930 201.275 21.120 201.995 ;
        RECT 19.930 200.795 20.760 201.095 ;
        RECT 21.290 201.065 21.610 202.025 ;
        RECT 18.515 200.395 18.850 200.565 ;
        RECT 19.045 200.395 19.720 200.565 ;
        RECT 20.040 200.115 20.410 200.615 ;
        RECT 20.590 200.565 20.760 200.795 ;
        RECT 21.145 200.735 21.610 201.065 ;
        RECT 21.780 201.355 21.950 202.195 ;
        RECT 22.130 202.165 22.445 202.665 ;
        RECT 22.675 201.935 23.015 202.495 ;
        RECT 22.120 201.560 23.015 201.935 ;
        RECT 23.185 201.655 23.355 202.665 ;
        RECT 22.825 201.355 23.015 201.560 ;
        RECT 23.525 201.605 23.855 202.450 ;
        RECT 23.525 201.525 23.915 201.605 ;
        RECT 23.700 201.475 23.915 201.525 ;
        RECT 24.085 201.500 24.375 202.665 ;
        RECT 24.545 201.525 24.930 202.495 ;
        RECT 25.100 202.205 25.425 202.665 ;
        RECT 25.945 202.035 26.225 202.495 ;
        RECT 25.100 201.815 26.225 202.035 ;
        RECT 21.780 201.025 22.655 201.355 ;
        RECT 22.825 201.025 23.575 201.355 ;
        RECT 21.780 200.565 21.950 201.025 ;
        RECT 22.825 200.855 23.025 201.025 ;
        RECT 23.745 200.895 23.915 201.475 ;
        RECT 23.690 200.855 23.915 200.895 ;
        RECT 20.590 200.395 20.995 200.565 ;
        RECT 21.165 200.395 21.950 200.565 ;
        RECT 22.225 200.115 22.435 200.645 ;
        RECT 22.695 200.330 23.025 200.855 ;
        RECT 23.535 200.770 23.915 200.855 ;
        RECT 24.545 200.855 24.825 201.525 ;
        RECT 25.100 201.355 25.550 201.815 ;
        RECT 26.415 201.645 26.815 202.495 ;
        RECT 27.215 202.205 27.485 202.665 ;
        RECT 27.655 202.035 27.940 202.495 ;
        RECT 24.995 201.025 25.550 201.355 ;
        RECT 25.720 201.085 26.815 201.645 ;
        RECT 25.100 200.915 25.550 201.025 ;
        RECT 23.195 200.115 23.365 200.725 ;
        RECT 23.535 200.335 23.865 200.770 ;
        RECT 24.085 200.115 24.375 200.840 ;
        RECT 24.545 200.285 24.930 200.855 ;
        RECT 25.100 200.745 26.225 200.915 ;
        RECT 25.100 200.115 25.425 200.575 ;
        RECT 25.945 200.285 26.225 200.745 ;
        RECT 26.415 200.285 26.815 201.085 ;
        RECT 26.985 201.815 27.940 202.035 ;
        RECT 29.235 201.995 29.405 202.495 ;
        RECT 29.575 202.165 29.905 202.665 ;
        RECT 29.235 201.825 29.900 201.995 ;
        RECT 26.985 200.915 27.195 201.815 ;
        RECT 27.365 201.085 28.055 201.645 ;
        RECT 29.150 201.005 29.500 201.655 ;
        RECT 26.985 200.745 27.940 200.915 ;
        RECT 29.670 200.835 29.900 201.825 ;
        RECT 27.215 200.115 27.485 200.575 ;
        RECT 27.655 200.285 27.940 200.745 ;
        RECT 29.235 200.665 29.900 200.835 ;
        RECT 29.235 200.375 29.405 200.665 ;
        RECT 29.575 200.115 29.905 200.495 ;
        RECT 30.075 200.375 30.260 202.495 ;
        RECT 30.500 202.205 30.765 202.665 ;
        RECT 30.935 202.070 31.185 202.495 ;
        RECT 31.395 202.220 32.500 202.390 ;
        RECT 30.880 201.940 31.185 202.070 ;
        RECT 30.430 200.745 30.710 201.695 ;
        RECT 30.880 200.835 31.050 201.940 ;
        RECT 31.220 201.155 31.460 201.750 ;
        RECT 31.630 201.685 32.160 202.050 ;
        RECT 31.630 200.985 31.800 201.685 ;
        RECT 32.330 201.605 32.500 202.220 ;
        RECT 32.670 201.865 32.840 202.665 ;
        RECT 33.010 202.165 33.260 202.495 ;
        RECT 33.485 202.195 34.370 202.365 ;
        RECT 32.330 201.515 32.840 201.605 ;
        RECT 30.880 200.705 31.105 200.835 ;
        RECT 31.275 200.765 31.800 200.985 ;
        RECT 31.970 201.345 32.840 201.515 ;
        RECT 30.515 200.115 30.765 200.575 ;
        RECT 30.935 200.565 31.105 200.705 ;
        RECT 31.970 200.565 32.140 201.345 ;
        RECT 32.670 201.275 32.840 201.345 ;
        RECT 32.350 201.095 32.550 201.125 ;
        RECT 33.010 201.095 33.180 202.165 ;
        RECT 33.350 201.275 33.540 201.995 ;
        RECT 32.350 200.795 33.180 201.095 ;
        RECT 33.710 201.065 34.030 202.025 ;
        RECT 30.935 200.395 31.270 200.565 ;
        RECT 31.465 200.395 32.140 200.565 ;
        RECT 32.460 200.115 32.830 200.615 ;
        RECT 33.010 200.565 33.180 200.795 ;
        RECT 33.565 200.735 34.030 201.065 ;
        RECT 34.200 201.355 34.370 202.195 ;
        RECT 34.550 202.165 34.865 202.665 ;
        RECT 35.095 201.935 35.435 202.495 ;
        RECT 34.540 201.560 35.435 201.935 ;
        RECT 35.605 201.655 35.775 202.665 ;
        RECT 35.245 201.355 35.435 201.560 ;
        RECT 35.945 201.605 36.275 202.450 ;
        RECT 36.445 201.750 36.615 202.665 ;
        RECT 35.945 201.525 36.335 201.605 ;
        RECT 37.430 201.525 37.685 202.665 ;
        RECT 37.880 202.115 39.075 202.445 ;
        RECT 36.120 201.475 36.335 201.525 ;
        RECT 34.200 201.025 35.075 201.355 ;
        RECT 35.245 201.025 35.995 201.355 ;
        RECT 34.200 200.565 34.370 201.025 ;
        RECT 35.245 200.855 35.445 201.025 ;
        RECT 36.165 200.895 36.335 201.475 ;
        RECT 37.935 201.355 38.105 201.915 ;
        RECT 38.330 201.695 38.750 201.945 ;
        RECT 39.255 201.865 39.535 202.665 ;
        RECT 38.330 201.525 39.575 201.695 ;
        RECT 39.745 201.525 40.015 202.495 ;
        RECT 39.405 201.355 39.575 201.525 ;
        RECT 37.430 201.105 37.765 201.355 ;
        RECT 37.935 201.025 38.675 201.355 ;
        RECT 39.405 201.025 39.635 201.355 ;
        RECT 37.935 200.935 38.185 201.025 ;
        RECT 36.110 200.855 36.335 200.895 ;
        RECT 33.010 200.395 33.415 200.565 ;
        RECT 33.585 200.395 34.370 200.565 ;
        RECT 34.645 200.115 34.855 200.645 ;
        RECT 35.115 200.330 35.445 200.855 ;
        RECT 35.955 200.770 36.335 200.855 ;
        RECT 35.615 200.115 35.785 200.725 ;
        RECT 35.955 200.335 36.285 200.770 ;
        RECT 37.450 200.765 38.185 200.935 ;
        RECT 39.405 200.855 39.575 201.025 ;
        RECT 36.455 200.115 36.625 200.630 ;
        RECT 37.450 200.295 37.760 200.765 ;
        RECT 38.835 200.685 39.575 200.855 ;
        RECT 39.845 200.790 40.015 201.525 ;
        RECT 37.930 200.115 38.665 200.595 ;
        RECT 38.835 200.335 39.005 200.685 ;
        RECT 39.175 200.115 39.555 200.515 ;
        RECT 39.745 200.445 40.015 200.790 ;
        RECT 40.205 201.610 40.510 202.395 ;
        RECT 40.690 202.195 41.375 202.665 ;
        RECT 40.685 201.675 41.380 201.985 ;
        RECT 40.205 200.805 40.380 201.610 ;
        RECT 41.555 201.505 41.840 202.450 ;
        RECT 42.015 202.215 42.345 202.665 ;
        RECT 42.515 202.045 42.685 202.475 ;
        RECT 40.980 201.355 41.840 201.505 ;
        RECT 40.555 201.335 41.840 201.355 ;
        RECT 42.010 201.815 42.685 202.045 ;
        RECT 40.555 200.975 41.540 201.335 ;
        RECT 42.010 201.165 42.245 201.815 ;
        RECT 42.955 201.715 43.230 202.485 ;
        RECT 43.400 202.055 43.730 202.485 ;
        RECT 43.900 202.225 44.095 202.665 ;
        RECT 44.275 202.055 44.605 202.485 ;
        RECT 43.400 201.885 44.605 202.055 ;
        RECT 40.205 200.285 40.445 200.805 ;
        RECT 41.370 200.640 41.540 200.975 ;
        RECT 41.710 200.835 42.245 201.165 ;
        RECT 42.025 200.685 42.245 200.835 ;
        RECT 42.415 200.795 42.715 201.645 ;
        RECT 42.955 201.525 43.540 201.715 ;
        RECT 43.710 201.555 44.605 201.885 ;
        RECT 44.785 201.575 48.295 202.665 ;
        RECT 48.465 201.575 49.675 202.665 ;
        RECT 42.955 200.705 43.195 201.355 ;
        RECT 43.365 200.855 43.540 201.525 ;
        RECT 43.710 201.025 44.125 201.355 ;
        RECT 44.305 201.025 44.600 201.355 ;
        RECT 40.615 200.115 41.010 200.610 ;
        RECT 41.370 200.445 41.745 200.640 ;
        RECT 41.575 200.300 41.745 200.445 ;
        RECT 42.025 200.310 42.265 200.685 ;
        RECT 43.365 200.675 43.695 200.855 ;
        RECT 42.435 200.115 42.770 200.620 ;
        RECT 42.970 200.115 43.300 200.505 ;
        RECT 43.470 200.295 43.695 200.675 ;
        RECT 43.895 200.405 44.125 201.025 ;
        RECT 44.785 200.885 46.435 201.405 ;
        RECT 46.605 201.055 48.295 201.575 ;
        RECT 44.305 200.115 44.605 200.845 ;
        RECT 44.785 200.115 48.295 200.885 ;
        RECT 48.465 200.865 48.985 201.405 ;
        RECT 49.155 201.035 49.675 201.575 ;
        RECT 49.845 201.500 50.135 202.665 ;
        RECT 48.465 200.115 49.675 200.865 ;
        RECT 49.845 200.115 50.135 200.840 ;
        RECT 50.315 200.295 50.575 202.485 ;
        RECT 50.745 201.935 51.085 202.665 ;
        RECT 51.265 201.755 51.535 202.485 ;
        RECT 50.765 201.535 51.535 201.755 ;
        RECT 51.715 201.775 51.945 202.485 ;
        RECT 52.115 201.955 52.445 202.665 ;
        RECT 52.615 201.775 52.875 202.485 ;
        RECT 53.065 202.230 58.410 202.665 ;
        RECT 51.715 201.535 52.875 201.775 ;
        RECT 50.765 200.865 51.055 201.535 ;
        RECT 51.235 201.045 51.700 201.355 ;
        RECT 51.880 201.045 52.405 201.355 ;
        RECT 50.765 200.665 51.995 200.865 ;
        RECT 50.835 200.115 51.505 200.485 ;
        RECT 51.685 200.295 51.995 200.665 ;
        RECT 52.175 200.405 52.405 201.045 ;
        RECT 52.585 201.025 52.885 201.355 ;
        RECT 52.585 200.115 52.875 200.845 ;
        RECT 54.650 200.660 54.990 201.490 ;
        RECT 56.470 200.980 56.820 202.230 ;
        RECT 58.585 201.575 61.175 202.665 ;
        RECT 61.435 202.045 61.605 202.475 ;
        RECT 61.775 202.215 62.105 202.665 ;
        RECT 61.435 201.815 62.110 202.045 ;
        RECT 58.585 200.885 59.795 201.405 ;
        RECT 59.965 201.055 61.175 201.575 ;
        RECT 53.065 200.115 58.410 200.660 ;
        RECT 58.585 200.115 61.175 200.885 ;
        RECT 61.405 200.795 61.705 201.645 ;
        RECT 61.875 201.165 62.110 201.815 ;
        RECT 62.280 201.505 62.565 202.450 ;
        RECT 62.745 202.195 63.430 202.665 ;
        RECT 62.740 201.675 63.435 201.985 ;
        RECT 63.610 201.610 63.915 202.395 ;
        RECT 62.280 201.355 63.140 201.505 ;
        RECT 63.705 201.475 63.915 201.610 ;
        RECT 62.280 201.335 63.565 201.355 ;
        RECT 61.875 200.835 62.410 201.165 ;
        RECT 62.580 200.975 63.565 201.335 ;
        RECT 61.875 200.685 62.095 200.835 ;
        RECT 61.350 200.115 61.685 200.620 ;
        RECT 61.855 200.310 62.095 200.685 ;
        RECT 62.580 200.640 62.750 200.975 ;
        RECT 63.740 200.805 63.915 201.475 ;
        RECT 62.375 200.445 62.750 200.640 ;
        RECT 62.375 200.300 62.545 200.445 ;
        RECT 63.110 200.115 63.505 200.610 ;
        RECT 63.675 200.285 63.915 200.805 ;
        RECT 64.115 200.295 64.375 202.485 ;
        RECT 64.545 201.935 64.885 202.665 ;
        RECT 65.065 201.755 65.335 202.485 ;
        RECT 64.565 201.535 65.335 201.755 ;
        RECT 65.515 201.775 65.745 202.485 ;
        RECT 65.915 201.955 66.245 202.665 ;
        RECT 66.415 201.775 66.675 202.485 ;
        RECT 65.515 201.535 66.675 201.775 ;
        RECT 64.565 200.865 64.855 201.535 ;
        RECT 66.865 201.525 67.135 202.495 ;
        RECT 67.345 201.865 67.625 202.665 ;
        RECT 67.805 202.115 69.000 202.445 ;
        RECT 68.130 201.695 68.550 201.945 ;
        RECT 67.305 201.525 68.550 201.695 ;
        RECT 65.035 201.045 65.500 201.355 ;
        RECT 65.680 201.045 66.205 201.355 ;
        RECT 64.565 200.665 65.795 200.865 ;
        RECT 64.635 200.115 65.305 200.485 ;
        RECT 65.485 200.295 65.795 200.665 ;
        RECT 65.975 200.405 66.205 201.045 ;
        RECT 66.385 201.025 66.685 201.355 ;
        RECT 66.385 200.115 66.675 200.845 ;
        RECT 66.865 200.790 67.035 201.525 ;
        RECT 67.305 201.355 67.475 201.525 ;
        RECT 68.775 201.355 68.945 201.915 ;
        RECT 69.195 201.525 69.450 202.665 ;
        RECT 69.625 201.575 70.835 202.665 ;
        RECT 67.245 201.025 67.475 201.355 ;
        RECT 68.205 201.025 68.945 201.355 ;
        RECT 69.115 201.105 69.450 201.355 ;
        RECT 67.305 200.855 67.475 201.025 ;
        RECT 68.695 200.935 68.945 201.025 ;
        RECT 66.865 200.445 67.135 200.790 ;
        RECT 67.305 200.685 68.045 200.855 ;
        RECT 68.695 200.765 69.430 200.935 ;
        RECT 67.325 200.115 67.705 200.515 ;
        RECT 67.875 200.335 68.045 200.685 ;
        RECT 68.215 200.115 68.950 200.595 ;
        RECT 69.120 200.295 69.430 200.765 ;
        RECT 69.625 200.865 70.145 201.405 ;
        RECT 70.315 201.035 70.835 201.575 ;
        RECT 71.040 201.875 71.575 202.495 ;
        RECT 69.625 200.115 70.835 200.865 ;
        RECT 71.040 200.855 71.355 201.875 ;
        RECT 71.745 201.865 72.075 202.665 ;
        RECT 72.560 201.695 72.950 201.870 ;
        RECT 71.525 201.525 72.950 201.695 ;
        RECT 73.305 201.525 73.585 202.665 ;
        RECT 71.525 201.025 71.695 201.525 ;
        RECT 71.040 200.285 71.655 200.855 ;
        RECT 71.945 200.795 72.210 201.355 ;
        RECT 72.380 200.625 72.550 201.525 ;
        RECT 73.755 201.515 74.085 202.495 ;
        RECT 74.255 201.525 74.515 202.665 ;
        RECT 72.720 200.795 73.075 201.355 ;
        RECT 73.315 201.085 73.650 201.355 ;
        RECT 73.820 200.915 73.990 201.515 ;
        RECT 75.605 201.500 75.895 202.665 ;
        RECT 76.065 202.230 81.410 202.665 ;
        RECT 74.160 201.105 74.495 201.355 ;
        RECT 71.825 200.115 72.040 200.625 ;
        RECT 72.270 200.295 72.550 200.625 ;
        RECT 72.730 200.115 72.970 200.625 ;
        RECT 73.305 200.115 73.615 200.915 ;
        RECT 73.820 200.285 74.515 200.915 ;
        RECT 75.605 200.115 75.895 200.840 ;
        RECT 77.650 200.660 77.990 201.490 ;
        RECT 79.470 200.980 79.820 202.230 ;
        RECT 81.585 201.575 82.795 202.665 ;
        RECT 82.965 202.155 83.225 202.665 ;
        RECT 81.585 200.865 82.105 201.405 ;
        RECT 82.275 201.035 82.795 201.575 ;
        RECT 82.965 201.105 83.305 201.985 ;
        RECT 83.475 201.275 83.645 202.495 ;
        RECT 83.885 202.160 84.500 202.665 ;
        RECT 83.885 201.625 84.135 201.990 ;
        RECT 84.305 201.985 84.500 202.160 ;
        RECT 84.670 202.155 85.145 202.495 ;
        RECT 85.315 202.120 85.530 202.665 ;
        RECT 84.305 201.795 84.635 201.985 ;
        RECT 84.855 201.625 85.570 201.920 ;
        RECT 85.740 201.795 86.015 202.495 ;
        RECT 83.885 201.455 85.675 201.625 ;
        RECT 83.475 201.025 84.270 201.275 ;
        RECT 83.475 200.935 83.725 201.025 ;
        RECT 76.065 200.115 81.410 200.660 ;
        RECT 81.585 200.115 82.795 200.865 ;
        RECT 82.965 200.115 83.225 200.935 ;
        RECT 83.395 200.515 83.725 200.935 ;
        RECT 84.440 200.600 84.695 201.455 ;
        RECT 83.905 200.335 84.695 200.600 ;
        RECT 84.865 200.755 85.275 201.275 ;
        RECT 85.445 201.025 85.675 201.455 ;
        RECT 85.845 200.765 86.015 201.795 ;
        RECT 86.185 201.575 88.775 202.665 ;
        RECT 84.865 200.335 85.065 200.755 ;
        RECT 85.255 200.115 85.585 200.575 ;
        RECT 85.755 200.285 86.015 200.765 ;
        RECT 86.185 200.885 87.395 201.405 ;
        RECT 87.565 201.055 88.775 201.575 ;
        RECT 89.035 201.735 89.205 202.495 ;
        RECT 89.385 201.905 89.715 202.665 ;
        RECT 89.035 201.565 89.700 201.735 ;
        RECT 89.885 201.590 90.155 202.495 ;
        RECT 90.325 202.230 95.670 202.665 ;
        RECT 89.530 201.420 89.700 201.565 ;
        RECT 88.965 201.015 89.295 201.385 ;
        RECT 89.530 201.090 89.815 201.420 ;
        RECT 86.185 200.115 88.775 200.885 ;
        RECT 89.530 200.835 89.700 201.090 ;
        RECT 89.035 200.665 89.700 200.835 ;
        RECT 89.985 200.790 90.155 201.590 ;
        RECT 89.035 200.285 89.205 200.665 ;
        RECT 89.385 200.115 89.715 200.495 ;
        RECT 89.895 200.285 90.155 200.790 ;
        RECT 91.910 200.660 92.250 201.490 ;
        RECT 93.730 200.980 94.080 202.230 ;
        RECT 95.845 201.575 99.355 202.665 ;
        RECT 95.845 200.885 97.495 201.405 ;
        RECT 97.665 201.055 99.355 201.575 ;
        RECT 100.075 201.735 100.245 202.495 ;
        RECT 100.425 201.905 100.755 202.665 ;
        RECT 100.075 201.565 100.740 201.735 ;
        RECT 100.925 201.590 101.195 202.495 ;
        RECT 100.570 201.420 100.740 201.565 ;
        RECT 100.005 201.015 100.335 201.385 ;
        RECT 100.570 201.090 100.855 201.420 ;
        RECT 90.325 200.115 95.670 200.660 ;
        RECT 95.845 200.115 99.355 200.885 ;
        RECT 100.570 200.835 100.740 201.090 ;
        RECT 100.075 200.665 100.740 200.835 ;
        RECT 101.025 200.790 101.195 201.590 ;
        RECT 101.365 201.500 101.655 202.665 ;
        RECT 101.885 201.605 102.215 202.450 ;
        RECT 102.385 201.655 102.555 202.665 ;
        RECT 102.725 201.935 103.065 202.495 ;
        RECT 103.295 202.165 103.610 202.665 ;
        RECT 103.790 202.195 104.675 202.365 ;
        RECT 101.825 201.525 102.215 201.605 ;
        RECT 102.725 201.560 103.620 201.935 ;
        RECT 101.825 201.475 102.040 201.525 ;
        RECT 101.825 200.895 101.995 201.475 ;
        RECT 102.725 201.355 102.915 201.560 ;
        RECT 103.790 201.355 103.960 202.195 ;
        RECT 104.900 202.165 105.150 202.495 ;
        RECT 102.165 201.025 102.915 201.355 ;
        RECT 103.085 201.025 103.960 201.355 ;
        RECT 101.825 200.855 102.050 200.895 ;
        RECT 102.715 200.855 102.915 201.025 ;
        RECT 100.075 200.285 100.245 200.665 ;
        RECT 100.425 200.115 100.755 200.495 ;
        RECT 100.935 200.285 101.195 200.790 ;
        RECT 101.365 200.115 101.655 200.840 ;
        RECT 101.825 200.770 102.205 200.855 ;
        RECT 101.875 200.335 102.205 200.770 ;
        RECT 102.375 200.115 102.545 200.725 ;
        RECT 102.715 200.330 103.045 200.855 ;
        RECT 103.305 200.115 103.515 200.645 ;
        RECT 103.790 200.565 103.960 201.025 ;
        RECT 104.130 201.065 104.450 202.025 ;
        RECT 104.620 201.275 104.810 201.995 ;
        RECT 104.980 201.095 105.150 202.165 ;
        RECT 105.320 201.865 105.490 202.665 ;
        RECT 105.660 202.220 106.765 202.390 ;
        RECT 105.660 201.605 105.830 202.220 ;
        RECT 106.975 202.070 107.225 202.495 ;
        RECT 107.395 202.205 107.660 202.665 ;
        RECT 106.000 201.685 106.530 202.050 ;
        RECT 106.975 201.940 107.280 202.070 ;
        RECT 105.320 201.515 105.830 201.605 ;
        RECT 105.320 201.345 106.190 201.515 ;
        RECT 105.320 201.275 105.490 201.345 ;
        RECT 105.610 201.095 105.810 201.125 ;
        RECT 104.130 200.735 104.595 201.065 ;
        RECT 104.980 200.795 105.810 201.095 ;
        RECT 104.980 200.565 105.150 200.795 ;
        RECT 103.790 200.395 104.575 200.565 ;
        RECT 104.745 200.395 105.150 200.565 ;
        RECT 105.330 200.115 105.700 200.615 ;
        RECT 106.020 200.565 106.190 201.345 ;
        RECT 106.360 200.985 106.530 201.685 ;
        RECT 106.700 201.155 106.940 201.750 ;
        RECT 106.360 200.765 106.885 200.985 ;
        RECT 107.110 200.835 107.280 201.940 ;
        RECT 107.055 200.705 107.280 200.835 ;
        RECT 107.450 200.745 107.730 201.695 ;
        RECT 107.055 200.565 107.225 200.705 ;
        RECT 106.020 200.395 106.695 200.565 ;
        RECT 106.890 200.395 107.225 200.565 ;
        RECT 107.395 200.115 107.645 200.575 ;
        RECT 107.900 200.375 108.085 202.495 ;
        RECT 108.255 202.165 108.585 202.665 ;
        RECT 108.755 201.995 108.925 202.495 ;
        RECT 108.260 201.825 108.925 201.995 ;
        RECT 109.760 202.035 110.045 202.495 ;
        RECT 110.215 202.205 110.485 202.665 ;
        RECT 108.260 200.835 108.490 201.825 ;
        RECT 109.760 201.815 110.715 202.035 ;
        RECT 108.660 201.005 109.010 201.655 ;
        RECT 109.645 201.085 110.335 201.645 ;
        RECT 110.505 200.915 110.715 201.815 ;
        RECT 108.260 200.665 108.925 200.835 ;
        RECT 108.255 200.115 108.585 200.495 ;
        RECT 108.755 200.375 108.925 200.665 ;
        RECT 109.760 200.745 110.715 200.915 ;
        RECT 110.885 201.645 111.285 202.495 ;
        RECT 111.475 202.035 111.755 202.495 ;
        RECT 112.275 202.205 112.600 202.665 ;
        RECT 111.475 201.815 112.600 202.035 ;
        RECT 110.885 201.085 111.980 201.645 ;
        RECT 112.150 201.355 112.600 201.815 ;
        RECT 112.770 201.525 113.155 202.495 ;
        RECT 113.325 201.575 114.535 202.665 ;
        RECT 114.795 201.995 114.965 202.495 ;
        RECT 115.135 202.165 115.465 202.665 ;
        RECT 114.795 201.825 115.460 201.995 ;
        RECT 109.760 200.285 110.045 200.745 ;
        RECT 110.215 200.115 110.485 200.575 ;
        RECT 110.885 200.285 111.285 201.085 ;
        RECT 112.150 201.025 112.705 201.355 ;
        RECT 112.150 200.915 112.600 201.025 ;
        RECT 111.475 200.745 112.600 200.915 ;
        RECT 112.875 200.855 113.155 201.525 ;
        RECT 111.475 200.285 111.755 200.745 ;
        RECT 112.275 200.115 112.600 200.575 ;
        RECT 112.770 200.285 113.155 200.855 ;
        RECT 113.325 200.865 113.845 201.405 ;
        RECT 114.015 201.035 114.535 201.575 ;
        RECT 114.710 201.005 115.060 201.655 ;
        RECT 113.325 200.115 114.535 200.865 ;
        RECT 115.230 200.835 115.460 201.825 ;
        RECT 114.795 200.665 115.460 200.835 ;
        RECT 114.795 200.375 114.965 200.665 ;
        RECT 115.135 200.115 115.465 200.495 ;
        RECT 115.635 200.375 115.820 202.495 ;
        RECT 116.060 202.205 116.325 202.665 ;
        RECT 116.495 202.070 116.745 202.495 ;
        RECT 116.955 202.220 118.060 202.390 ;
        RECT 116.440 201.940 116.745 202.070 ;
        RECT 115.990 200.745 116.270 201.695 ;
        RECT 116.440 200.835 116.610 201.940 ;
        RECT 116.780 201.155 117.020 201.750 ;
        RECT 117.190 201.685 117.720 202.050 ;
        RECT 117.190 200.985 117.360 201.685 ;
        RECT 117.890 201.605 118.060 202.220 ;
        RECT 118.230 201.865 118.400 202.665 ;
        RECT 118.570 202.165 118.820 202.495 ;
        RECT 119.045 202.195 119.930 202.365 ;
        RECT 117.890 201.515 118.400 201.605 ;
        RECT 116.440 200.705 116.665 200.835 ;
        RECT 116.835 200.765 117.360 200.985 ;
        RECT 117.530 201.345 118.400 201.515 ;
        RECT 116.075 200.115 116.325 200.575 ;
        RECT 116.495 200.565 116.665 200.705 ;
        RECT 117.530 200.565 117.700 201.345 ;
        RECT 118.230 201.275 118.400 201.345 ;
        RECT 117.910 201.095 118.110 201.125 ;
        RECT 118.570 201.095 118.740 202.165 ;
        RECT 118.910 201.275 119.100 201.995 ;
        RECT 117.910 200.795 118.740 201.095 ;
        RECT 119.270 201.065 119.590 202.025 ;
        RECT 116.495 200.395 116.830 200.565 ;
        RECT 117.025 200.395 117.700 200.565 ;
        RECT 118.020 200.115 118.390 200.615 ;
        RECT 118.570 200.565 118.740 200.795 ;
        RECT 119.125 200.735 119.590 201.065 ;
        RECT 119.760 201.355 119.930 202.195 ;
        RECT 120.110 202.165 120.425 202.665 ;
        RECT 120.655 201.935 120.995 202.495 ;
        RECT 120.100 201.560 120.995 201.935 ;
        RECT 121.165 201.655 121.335 202.665 ;
        RECT 120.805 201.355 120.995 201.560 ;
        RECT 121.505 201.605 121.835 202.450 ;
        RECT 122.005 201.750 122.175 202.665 ;
        RECT 121.505 201.525 121.895 201.605 ;
        RECT 122.525 201.575 126.035 202.665 ;
        RECT 121.680 201.475 121.895 201.525 ;
        RECT 119.760 201.025 120.635 201.355 ;
        RECT 120.805 201.025 121.555 201.355 ;
        RECT 119.760 200.565 119.930 201.025 ;
        RECT 120.805 200.855 121.005 201.025 ;
        RECT 121.725 200.895 121.895 201.475 ;
        RECT 121.670 200.855 121.895 200.895 ;
        RECT 118.570 200.395 118.975 200.565 ;
        RECT 119.145 200.395 119.930 200.565 ;
        RECT 120.205 200.115 120.415 200.645 ;
        RECT 120.675 200.330 121.005 200.855 ;
        RECT 121.515 200.770 121.895 200.855 ;
        RECT 122.525 200.885 124.175 201.405 ;
        RECT 124.345 201.055 126.035 201.575 ;
        RECT 127.125 201.500 127.415 202.665 ;
        RECT 127.585 202.230 132.930 202.665 ;
        RECT 133.105 202.230 138.450 202.665 ;
        RECT 138.625 202.230 143.970 202.665 ;
        RECT 121.175 200.115 121.345 200.725 ;
        RECT 121.515 200.335 121.845 200.770 ;
        RECT 122.015 200.115 122.185 200.630 ;
        RECT 122.525 200.115 126.035 200.885 ;
        RECT 127.125 200.115 127.415 200.840 ;
        RECT 129.170 200.660 129.510 201.490 ;
        RECT 130.990 200.980 131.340 202.230 ;
        RECT 134.690 200.660 135.030 201.490 ;
        RECT 136.510 200.980 136.860 202.230 ;
        RECT 140.210 200.660 140.550 201.490 ;
        RECT 142.030 200.980 142.380 202.230 ;
        RECT 144.145 201.575 147.655 202.665 ;
        RECT 147.825 201.575 149.035 202.665 ;
        RECT 144.145 200.885 145.795 201.405 ;
        RECT 145.965 201.055 147.655 201.575 ;
        RECT 127.585 200.115 132.930 200.660 ;
        RECT 133.105 200.115 138.450 200.660 ;
        RECT 138.625 200.115 143.970 200.660 ;
        RECT 144.145 200.115 147.655 200.885 ;
        RECT 147.825 200.865 148.345 201.405 ;
        RECT 148.515 201.035 149.035 201.575 ;
        RECT 149.205 201.575 150.415 202.665 ;
        RECT 149.205 201.035 149.725 201.575 ;
        RECT 149.895 200.865 150.415 201.405 ;
        RECT 147.825 200.115 149.035 200.865 ;
        RECT 149.205 200.115 150.415 200.865 ;
        RECT 11.120 199.945 150.500 200.115 ;
        RECT 11.205 199.195 12.415 199.945 ;
        RECT 12.585 199.400 17.930 199.945 ;
        RECT 11.205 198.655 11.725 199.195 ;
        RECT 11.895 198.485 12.415 199.025 ;
        RECT 14.170 198.570 14.510 199.400 ;
        RECT 18.105 199.175 21.615 199.945 ;
        RECT 21.785 199.195 22.995 199.945 ;
        RECT 23.190 199.555 23.520 199.945 ;
        RECT 23.690 199.385 23.915 199.765 ;
        RECT 11.205 197.395 12.415 198.485 ;
        RECT 15.990 197.830 16.340 199.080 ;
        RECT 18.105 198.655 19.755 199.175 ;
        RECT 19.925 198.485 21.615 199.005 ;
        RECT 21.785 198.655 22.305 199.195 ;
        RECT 22.475 198.485 22.995 199.025 ;
        RECT 23.175 198.705 23.415 199.355 ;
        RECT 23.585 199.205 23.915 199.385 ;
        RECT 23.585 198.535 23.760 199.205 ;
        RECT 24.115 199.035 24.345 199.655 ;
        RECT 24.525 199.215 24.825 199.945 ;
        RECT 25.010 199.415 25.300 199.765 ;
        RECT 25.495 199.585 25.825 199.945 ;
        RECT 25.995 199.415 26.225 199.720 ;
        RECT 25.010 199.245 26.225 199.415 ;
        RECT 26.415 199.075 26.585 199.640 ;
        RECT 23.930 198.705 24.345 199.035 ;
        RECT 24.525 198.705 24.820 199.035 ;
        RECT 25.070 198.925 25.330 199.035 ;
        RECT 25.065 198.755 25.330 198.925 ;
        RECT 25.070 198.705 25.330 198.755 ;
        RECT 25.510 198.705 25.895 199.035 ;
        RECT 26.065 198.905 26.585 199.075 ;
        RECT 26.845 199.295 27.105 199.775 ;
        RECT 27.275 199.405 27.525 199.945 ;
        RECT 12.585 197.395 17.930 197.830 ;
        RECT 18.105 197.395 21.615 198.485 ;
        RECT 21.785 197.395 22.995 198.485 ;
        RECT 23.175 198.345 23.760 198.535 ;
        RECT 23.175 197.575 23.450 198.345 ;
        RECT 23.930 198.175 24.825 198.505 ;
        RECT 23.620 198.005 24.825 198.175 ;
        RECT 23.620 197.575 23.950 198.005 ;
        RECT 24.120 197.395 24.315 197.835 ;
        RECT 24.495 197.575 24.825 198.005 ;
        RECT 25.010 197.395 25.330 198.535 ;
        RECT 25.510 197.655 25.705 198.705 ;
        RECT 26.065 198.525 26.235 198.905 ;
        RECT 25.885 198.245 26.235 198.525 ;
        RECT 26.425 198.375 26.670 198.735 ;
        RECT 26.845 198.265 27.015 199.295 ;
        RECT 27.695 199.240 27.915 199.725 ;
        RECT 27.185 198.645 27.415 199.040 ;
        RECT 27.585 198.815 27.915 199.240 ;
        RECT 28.085 199.565 28.975 199.735 ;
        RECT 28.085 198.840 28.255 199.565 ;
        RECT 28.425 199.010 28.975 199.395 ;
        RECT 29.145 199.175 31.735 199.945 ;
        RECT 31.905 199.270 32.165 199.775 ;
        RECT 32.345 199.565 32.675 199.945 ;
        RECT 32.855 199.395 33.025 199.775 ;
        RECT 28.085 198.770 28.975 198.840 ;
        RECT 28.080 198.745 28.975 198.770 ;
        RECT 28.070 198.730 28.975 198.745 ;
        RECT 28.065 198.715 28.975 198.730 ;
        RECT 28.055 198.710 28.975 198.715 ;
        RECT 28.050 198.700 28.975 198.710 ;
        RECT 28.045 198.690 28.975 198.700 ;
        RECT 28.035 198.685 28.975 198.690 ;
        RECT 28.025 198.675 28.975 198.685 ;
        RECT 28.015 198.670 28.975 198.675 ;
        RECT 28.015 198.665 28.350 198.670 ;
        RECT 28.000 198.660 28.350 198.665 ;
        RECT 27.985 198.650 28.350 198.660 ;
        RECT 27.960 198.645 28.350 198.650 ;
        RECT 27.185 198.640 28.350 198.645 ;
        RECT 27.185 198.605 28.320 198.640 ;
        RECT 27.185 198.580 28.285 198.605 ;
        RECT 27.185 198.550 28.255 198.580 ;
        RECT 27.185 198.520 28.235 198.550 ;
        RECT 27.185 198.490 28.215 198.520 ;
        RECT 27.185 198.480 28.145 198.490 ;
        RECT 27.185 198.470 28.120 198.480 ;
        RECT 27.185 198.455 28.100 198.470 ;
        RECT 27.185 198.440 28.080 198.455 ;
        RECT 27.290 198.430 28.075 198.440 ;
        RECT 27.290 198.395 28.060 198.430 ;
        RECT 25.885 197.565 26.215 198.245 ;
        RECT 26.415 197.395 26.670 198.195 ;
        RECT 26.845 197.565 27.120 198.265 ;
        RECT 27.290 198.145 28.045 198.395 ;
        RECT 28.215 198.075 28.545 198.320 ;
        RECT 28.715 198.220 28.975 198.670 ;
        RECT 29.145 198.655 30.355 199.175 ;
        RECT 30.525 198.485 31.735 199.005 ;
        RECT 28.360 198.050 28.545 198.075 ;
        RECT 28.360 197.950 28.975 198.050 ;
        RECT 27.290 197.395 27.545 197.940 ;
        RECT 27.715 197.565 28.195 197.905 ;
        RECT 28.370 197.395 28.975 197.950 ;
        RECT 29.145 197.395 31.735 198.485 ;
        RECT 31.905 198.470 32.075 199.270 ;
        RECT 32.360 199.225 33.025 199.395 ;
        RECT 32.360 198.970 32.530 199.225 ;
        RECT 33.285 199.175 36.795 199.945 ;
        RECT 36.965 199.220 37.255 199.945 ;
        RECT 37.425 199.400 42.770 199.945 ;
        RECT 32.245 198.640 32.530 198.970 ;
        RECT 32.765 198.675 33.095 199.045 ;
        RECT 33.285 198.655 34.935 199.175 ;
        RECT 32.360 198.495 32.530 198.640 ;
        RECT 31.905 197.565 32.175 198.470 ;
        RECT 32.360 198.325 33.025 198.495 ;
        RECT 35.105 198.485 36.795 199.005 ;
        RECT 39.010 198.570 39.350 199.400 ;
        RECT 42.945 199.175 46.455 199.945 ;
        RECT 32.345 197.395 32.675 198.155 ;
        RECT 32.855 197.565 33.025 198.325 ;
        RECT 33.285 197.395 36.795 198.485 ;
        RECT 36.965 197.395 37.255 198.560 ;
        RECT 40.830 197.830 41.180 199.080 ;
        RECT 42.945 198.655 44.595 199.175 ;
        RECT 47.565 199.135 47.805 199.945 ;
        RECT 47.975 199.135 48.305 199.775 ;
        RECT 48.475 199.135 48.745 199.945 ;
        RECT 48.925 199.145 49.235 199.945 ;
        RECT 49.440 199.145 50.135 199.775 ;
        RECT 51.225 199.205 51.690 199.750 ;
        RECT 44.765 198.485 46.455 199.005 ;
        RECT 47.545 198.705 47.895 198.955 ;
        RECT 48.065 198.535 48.235 199.135 ;
        RECT 48.405 198.705 48.755 198.955 ;
        RECT 48.935 198.705 49.270 198.975 ;
        RECT 49.440 198.545 49.610 199.145 ;
        RECT 49.780 198.705 50.115 198.955 ;
        RECT 37.425 197.395 42.770 197.830 ;
        RECT 42.945 197.395 46.455 198.485 ;
        RECT 47.555 198.365 48.235 198.535 ;
        RECT 47.555 197.580 47.885 198.365 ;
        RECT 48.415 197.395 48.745 198.535 ;
        RECT 48.925 197.395 49.205 198.535 ;
        RECT 49.375 197.565 49.705 198.545 ;
        RECT 49.875 197.395 50.135 198.535 ;
        RECT 51.225 198.245 51.395 199.205 ;
        RECT 52.195 199.125 52.365 199.945 ;
        RECT 52.535 199.295 52.865 199.775 ;
        RECT 53.035 199.555 53.385 199.945 ;
        RECT 53.555 199.375 53.785 199.775 ;
        RECT 53.275 199.295 53.785 199.375 ;
        RECT 52.535 199.205 53.785 199.295 ;
        RECT 53.955 199.205 54.275 199.685 ;
        RECT 54.445 199.400 59.790 199.945 ;
        RECT 52.535 199.125 53.445 199.205 ;
        RECT 51.565 198.585 51.810 199.035 ;
        RECT 52.070 198.755 52.765 198.955 ;
        RECT 52.935 198.785 53.535 198.955 ;
        RECT 52.935 198.585 53.105 198.785 ;
        RECT 53.765 198.615 53.935 199.035 ;
        RECT 51.565 198.415 53.105 198.585 ;
        RECT 53.275 198.445 53.935 198.615 ;
        RECT 53.275 198.245 53.445 198.445 ;
        RECT 54.105 198.275 54.275 199.205 ;
        RECT 56.030 198.570 56.370 199.400 ;
        RECT 59.965 199.175 62.555 199.945 ;
        RECT 62.725 199.220 63.015 199.945 ;
        RECT 63.185 199.400 68.530 199.945 ;
        RECT 51.225 198.075 53.445 198.245 ;
        RECT 53.615 198.075 54.275 198.275 ;
        RECT 51.225 197.395 51.525 197.905 ;
        RECT 51.695 197.565 52.025 198.075 ;
        RECT 53.615 197.905 53.785 198.075 ;
        RECT 52.195 197.395 52.825 197.905 ;
        RECT 53.405 197.735 53.785 197.905 ;
        RECT 53.955 197.395 54.255 197.905 ;
        RECT 57.850 197.830 58.200 199.080 ;
        RECT 59.965 198.655 61.175 199.175 ;
        RECT 61.345 198.485 62.555 199.005 ;
        RECT 64.770 198.570 65.110 199.400 ;
        RECT 69.625 199.270 69.895 199.615 ;
        RECT 70.085 199.545 70.465 199.945 ;
        RECT 70.635 199.375 70.805 199.725 ;
        RECT 70.975 199.465 71.710 199.945 ;
        RECT 54.445 197.395 59.790 197.830 ;
        RECT 59.965 197.395 62.555 198.485 ;
        RECT 62.725 197.395 63.015 198.560 ;
        RECT 66.590 197.830 66.940 199.080 ;
        RECT 69.625 198.535 69.795 199.270 ;
        RECT 70.065 199.205 70.805 199.375 ;
        RECT 71.880 199.295 72.190 199.765 ;
        RECT 70.065 199.035 70.235 199.205 ;
        RECT 71.455 199.125 72.190 199.295 ;
        RECT 72.385 199.175 75.895 199.945 ;
        RECT 76.525 199.565 77.415 199.735 ;
        RECT 71.455 199.035 71.705 199.125 ;
        RECT 70.005 198.705 70.235 199.035 ;
        RECT 70.965 198.705 71.705 199.035 ;
        RECT 71.875 198.705 72.210 198.955 ;
        RECT 70.065 198.535 70.235 198.705 ;
        RECT 63.185 197.395 68.530 197.830 ;
        RECT 69.625 197.565 69.895 198.535 ;
        RECT 70.065 198.365 71.310 198.535 ;
        RECT 70.105 197.395 70.385 198.195 ;
        RECT 70.890 198.115 71.310 198.365 ;
        RECT 71.535 198.145 71.705 198.705 ;
        RECT 72.385 198.655 74.035 199.175 ;
        RECT 76.525 199.010 77.075 199.395 ;
        RECT 70.565 197.615 71.760 197.945 ;
        RECT 71.955 197.395 72.210 198.535 ;
        RECT 74.205 198.485 75.895 199.005 ;
        RECT 77.245 198.840 77.415 199.565 ;
        RECT 72.385 197.395 75.895 198.485 ;
        RECT 76.525 198.770 77.415 198.840 ;
        RECT 77.585 199.265 77.805 199.725 ;
        RECT 77.975 199.405 78.225 199.945 ;
        RECT 78.395 199.295 78.655 199.775 ;
        RECT 79.285 199.565 80.175 199.735 ;
        RECT 77.585 199.240 77.835 199.265 ;
        RECT 77.585 198.815 77.915 199.240 ;
        RECT 76.525 198.745 77.420 198.770 ;
        RECT 76.525 198.730 77.430 198.745 ;
        RECT 76.525 198.715 77.435 198.730 ;
        RECT 76.525 198.710 77.445 198.715 ;
        RECT 76.525 198.700 77.450 198.710 ;
        RECT 76.525 198.690 77.455 198.700 ;
        RECT 76.525 198.685 77.465 198.690 ;
        RECT 76.525 198.675 77.475 198.685 ;
        RECT 76.525 198.670 77.485 198.675 ;
        RECT 76.525 198.220 76.785 198.670 ;
        RECT 77.150 198.665 77.485 198.670 ;
        RECT 77.150 198.660 77.500 198.665 ;
        RECT 77.150 198.650 77.515 198.660 ;
        RECT 77.150 198.645 77.540 198.650 ;
        RECT 78.085 198.645 78.315 199.040 ;
        RECT 77.150 198.640 78.315 198.645 ;
        RECT 77.180 198.605 78.315 198.640 ;
        RECT 77.215 198.580 78.315 198.605 ;
        RECT 77.245 198.550 78.315 198.580 ;
        RECT 77.265 198.520 78.315 198.550 ;
        RECT 77.285 198.490 78.315 198.520 ;
        RECT 77.355 198.480 78.315 198.490 ;
        RECT 77.380 198.470 78.315 198.480 ;
        RECT 77.400 198.455 78.315 198.470 ;
        RECT 77.420 198.440 78.315 198.455 ;
        RECT 77.425 198.430 78.210 198.440 ;
        RECT 77.440 198.395 78.210 198.430 ;
        RECT 76.955 198.075 77.285 198.320 ;
        RECT 77.455 198.145 78.210 198.395 ;
        RECT 78.485 198.265 78.655 199.295 ;
        RECT 79.285 199.010 79.835 199.395 ;
        RECT 80.005 198.840 80.175 199.565 ;
        RECT 76.955 198.050 77.140 198.075 ;
        RECT 76.525 197.950 77.140 198.050 ;
        RECT 76.525 197.395 77.130 197.950 ;
        RECT 77.305 197.565 77.785 197.905 ;
        RECT 77.955 197.395 78.210 197.940 ;
        RECT 78.380 197.565 78.655 198.265 ;
        RECT 79.285 198.770 80.175 198.840 ;
        RECT 80.345 199.240 80.565 199.725 ;
        RECT 80.735 199.405 80.985 199.945 ;
        RECT 81.155 199.295 81.415 199.775 ;
        RECT 80.345 198.815 80.675 199.240 ;
        RECT 79.285 198.745 80.180 198.770 ;
        RECT 79.285 198.730 80.190 198.745 ;
        RECT 79.285 198.715 80.195 198.730 ;
        RECT 79.285 198.710 80.205 198.715 ;
        RECT 79.285 198.700 80.210 198.710 ;
        RECT 79.285 198.690 80.215 198.700 ;
        RECT 79.285 198.685 80.225 198.690 ;
        RECT 79.285 198.675 80.235 198.685 ;
        RECT 79.285 198.670 80.245 198.675 ;
        RECT 79.285 198.220 79.545 198.670 ;
        RECT 79.910 198.665 80.245 198.670 ;
        RECT 79.910 198.660 80.260 198.665 ;
        RECT 79.910 198.650 80.275 198.660 ;
        RECT 79.910 198.645 80.300 198.650 ;
        RECT 80.845 198.645 81.075 199.040 ;
        RECT 79.910 198.640 81.075 198.645 ;
        RECT 79.940 198.605 81.075 198.640 ;
        RECT 79.975 198.580 81.075 198.605 ;
        RECT 80.005 198.550 81.075 198.580 ;
        RECT 80.025 198.520 81.075 198.550 ;
        RECT 80.045 198.490 81.075 198.520 ;
        RECT 80.115 198.480 81.075 198.490 ;
        RECT 80.140 198.470 81.075 198.480 ;
        RECT 80.160 198.455 81.075 198.470 ;
        RECT 80.180 198.440 81.075 198.455 ;
        RECT 80.185 198.430 80.970 198.440 ;
        RECT 80.200 198.395 80.970 198.430 ;
        RECT 79.715 198.075 80.045 198.320 ;
        RECT 80.215 198.145 80.970 198.395 ;
        RECT 81.245 198.265 81.415 199.295 ;
        RECT 81.585 199.195 82.795 199.945 ;
        RECT 83.130 199.435 83.370 199.945 ;
        RECT 83.550 199.435 83.830 199.765 ;
        RECT 84.060 199.435 84.275 199.945 ;
        RECT 81.585 198.655 82.105 199.195 ;
        RECT 82.275 198.485 82.795 199.025 ;
        RECT 83.025 198.705 83.380 199.265 ;
        RECT 83.550 198.535 83.720 199.435 ;
        RECT 83.890 198.705 84.155 199.265 ;
        RECT 84.445 199.205 85.060 199.775 ;
        RECT 84.405 198.535 84.575 199.035 ;
        RECT 79.715 198.050 79.900 198.075 ;
        RECT 79.285 197.950 79.900 198.050 ;
        RECT 79.285 197.395 79.890 197.950 ;
        RECT 80.065 197.565 80.545 197.905 ;
        RECT 80.715 197.395 80.970 197.940 ;
        RECT 81.140 197.565 81.415 198.265 ;
        RECT 81.585 197.395 82.795 198.485 ;
        RECT 83.150 198.365 84.575 198.535 ;
        RECT 83.150 198.190 83.540 198.365 ;
        RECT 84.025 197.395 84.355 198.195 ;
        RECT 84.745 198.185 85.060 199.205 ;
        RECT 85.265 199.175 87.855 199.945 ;
        RECT 88.485 199.220 88.775 199.945 ;
        RECT 88.945 199.175 90.615 199.945 ;
        RECT 91.295 199.555 91.625 199.945 ;
        RECT 91.795 199.375 91.965 199.695 ;
        RECT 92.135 199.555 92.465 199.945 ;
        RECT 92.880 199.545 93.835 199.715 ;
        RECT 91.245 199.205 93.495 199.375 ;
        RECT 85.265 198.655 86.475 199.175 ;
        RECT 86.645 198.485 87.855 199.005 ;
        RECT 88.945 198.655 89.695 199.175 ;
        RECT 84.525 197.565 85.060 198.185 ;
        RECT 85.265 197.395 87.855 198.485 ;
        RECT 88.485 197.395 88.775 198.560 ;
        RECT 89.865 198.485 90.615 199.005 ;
        RECT 88.945 197.395 90.615 198.485 ;
        RECT 91.245 198.245 91.415 199.205 ;
        RECT 91.585 198.585 91.830 199.035 ;
        RECT 92.000 198.755 92.550 198.955 ;
        RECT 92.720 198.785 93.095 198.955 ;
        RECT 92.720 198.585 92.890 198.785 ;
        RECT 93.265 198.705 93.495 199.205 ;
        RECT 91.585 198.415 92.890 198.585 ;
        RECT 93.665 198.665 93.835 199.545 ;
        RECT 94.005 199.110 94.295 199.945 ;
        RECT 94.465 199.175 97.975 199.945 ;
        RECT 98.605 199.565 99.495 199.735 ;
        RECT 93.665 198.495 94.295 198.665 ;
        RECT 94.465 198.655 96.115 199.175 ;
        RECT 98.605 199.010 99.155 199.395 ;
        RECT 91.245 197.565 91.625 198.245 ;
        RECT 92.215 197.395 92.385 198.245 ;
        RECT 92.555 198.075 93.795 198.245 ;
        RECT 92.555 197.565 92.885 198.075 ;
        RECT 93.055 197.395 93.225 197.905 ;
        RECT 93.395 197.565 93.795 198.075 ;
        RECT 93.975 197.565 94.295 198.495 ;
        RECT 96.285 198.485 97.975 199.005 ;
        RECT 99.325 198.840 99.495 199.565 ;
        RECT 94.465 197.395 97.975 198.485 ;
        RECT 98.605 198.770 99.495 198.840 ;
        RECT 99.665 199.265 99.885 199.725 ;
        RECT 100.055 199.405 100.305 199.945 ;
        RECT 100.475 199.295 100.735 199.775 ;
        RECT 99.665 199.240 99.915 199.265 ;
        RECT 99.665 198.815 99.995 199.240 ;
        RECT 98.605 198.745 99.500 198.770 ;
        RECT 98.605 198.730 99.510 198.745 ;
        RECT 98.605 198.715 99.515 198.730 ;
        RECT 98.605 198.710 99.525 198.715 ;
        RECT 98.605 198.700 99.530 198.710 ;
        RECT 98.605 198.690 99.535 198.700 ;
        RECT 98.605 198.685 99.545 198.690 ;
        RECT 98.605 198.675 99.555 198.685 ;
        RECT 98.605 198.670 99.565 198.675 ;
        RECT 98.605 198.220 98.865 198.670 ;
        RECT 99.230 198.665 99.565 198.670 ;
        RECT 99.230 198.660 99.580 198.665 ;
        RECT 99.230 198.650 99.595 198.660 ;
        RECT 99.230 198.645 99.620 198.650 ;
        RECT 100.165 198.645 100.395 199.040 ;
        RECT 99.230 198.640 100.395 198.645 ;
        RECT 99.260 198.605 100.395 198.640 ;
        RECT 99.295 198.580 100.395 198.605 ;
        RECT 99.325 198.550 100.395 198.580 ;
        RECT 99.345 198.520 100.395 198.550 ;
        RECT 99.365 198.490 100.395 198.520 ;
        RECT 99.435 198.480 100.395 198.490 ;
        RECT 99.460 198.470 100.395 198.480 ;
        RECT 99.480 198.455 100.395 198.470 ;
        RECT 99.500 198.440 100.395 198.455 ;
        RECT 99.505 198.430 100.290 198.440 ;
        RECT 99.520 198.395 100.290 198.430 ;
        RECT 99.035 198.075 99.365 198.320 ;
        RECT 99.535 198.145 100.290 198.395 ;
        RECT 100.565 198.265 100.735 199.295 ;
        RECT 99.035 198.050 99.220 198.075 ;
        RECT 98.605 197.950 99.220 198.050 ;
        RECT 98.605 197.395 99.210 197.950 ;
        RECT 99.385 197.565 99.865 197.905 ;
        RECT 100.035 197.395 100.290 197.940 ;
        RECT 100.460 197.565 100.735 198.265 ;
        RECT 100.905 199.205 101.290 199.775 ;
        RECT 101.460 199.485 101.785 199.945 ;
        RECT 102.305 199.315 102.585 199.775 ;
        RECT 100.905 198.535 101.185 199.205 ;
        RECT 101.460 199.145 102.585 199.315 ;
        RECT 101.460 199.035 101.910 199.145 ;
        RECT 101.355 198.705 101.910 199.035 ;
        RECT 102.775 198.975 103.175 199.775 ;
        RECT 103.575 199.485 103.845 199.945 ;
        RECT 104.015 199.315 104.300 199.775 ;
        RECT 100.905 197.565 101.290 198.535 ;
        RECT 101.460 198.245 101.910 198.705 ;
        RECT 102.080 198.415 103.175 198.975 ;
        RECT 101.460 198.025 102.585 198.245 ;
        RECT 101.460 197.395 101.785 197.855 ;
        RECT 102.305 197.565 102.585 198.025 ;
        RECT 102.775 197.565 103.175 198.415 ;
        RECT 103.345 199.145 104.300 199.315 ;
        RECT 105.135 199.395 105.305 199.685 ;
        RECT 105.475 199.565 105.805 199.945 ;
        RECT 105.135 199.225 105.800 199.395 ;
        RECT 103.345 198.245 103.555 199.145 ;
        RECT 103.725 198.415 104.415 198.975 ;
        RECT 105.050 198.405 105.400 199.055 ;
        RECT 103.345 198.025 104.300 198.245 ;
        RECT 105.570 198.235 105.800 199.225 ;
        RECT 103.575 197.395 103.845 197.855 ;
        RECT 104.015 197.565 104.300 198.025 ;
        RECT 105.135 198.065 105.800 198.235 ;
        RECT 105.135 197.565 105.305 198.065 ;
        RECT 105.475 197.395 105.805 197.895 ;
        RECT 105.975 197.565 106.160 199.685 ;
        RECT 106.415 199.485 106.665 199.945 ;
        RECT 106.835 199.495 107.170 199.665 ;
        RECT 107.365 199.495 108.040 199.665 ;
        RECT 106.835 199.355 107.005 199.495 ;
        RECT 106.330 198.365 106.610 199.315 ;
        RECT 106.780 199.225 107.005 199.355 ;
        RECT 106.780 198.120 106.950 199.225 ;
        RECT 107.175 199.075 107.700 199.295 ;
        RECT 107.120 198.310 107.360 198.905 ;
        RECT 107.530 198.375 107.700 199.075 ;
        RECT 107.870 198.715 108.040 199.495 ;
        RECT 108.360 199.445 108.730 199.945 ;
        RECT 108.910 199.495 109.315 199.665 ;
        RECT 109.485 199.495 110.270 199.665 ;
        RECT 108.910 199.265 109.080 199.495 ;
        RECT 108.250 198.965 109.080 199.265 ;
        RECT 109.465 198.995 109.930 199.325 ;
        RECT 108.250 198.935 108.450 198.965 ;
        RECT 108.570 198.715 108.740 198.785 ;
        RECT 107.870 198.545 108.740 198.715 ;
        RECT 108.230 198.455 108.740 198.545 ;
        RECT 106.780 197.990 107.085 198.120 ;
        RECT 107.530 198.010 108.060 198.375 ;
        RECT 106.400 197.395 106.665 197.855 ;
        RECT 106.835 197.565 107.085 197.990 ;
        RECT 108.230 197.840 108.400 198.455 ;
        RECT 107.295 197.670 108.400 197.840 ;
        RECT 108.570 197.395 108.740 198.195 ;
        RECT 108.910 197.895 109.080 198.965 ;
        RECT 109.250 198.065 109.440 198.785 ;
        RECT 109.610 198.035 109.930 198.995 ;
        RECT 110.100 199.035 110.270 199.495 ;
        RECT 110.545 199.415 110.755 199.945 ;
        RECT 111.015 199.205 111.345 199.730 ;
        RECT 111.515 199.335 111.685 199.945 ;
        RECT 111.855 199.290 112.185 199.725 ;
        RECT 112.355 199.430 112.525 199.945 ;
        RECT 111.855 199.205 112.235 199.290 ;
        RECT 111.145 199.035 111.345 199.205 ;
        RECT 112.010 199.165 112.235 199.205 ;
        RECT 110.100 198.705 110.975 199.035 ;
        RECT 111.145 198.705 111.895 199.035 ;
        RECT 108.910 197.565 109.160 197.895 ;
        RECT 110.100 197.865 110.270 198.705 ;
        RECT 111.145 198.500 111.335 198.705 ;
        RECT 112.065 198.585 112.235 199.165 ;
        RECT 112.865 199.195 114.075 199.945 ;
        RECT 114.245 199.220 114.535 199.945 ;
        RECT 114.905 199.315 115.235 199.675 ;
        RECT 115.855 199.485 116.105 199.945 ;
        RECT 116.275 199.485 116.835 199.775 ;
        RECT 112.865 198.655 113.385 199.195 ;
        RECT 114.905 199.125 116.295 199.315 ;
        RECT 116.125 199.035 116.295 199.125 ;
        RECT 112.020 198.535 112.235 198.585 ;
        RECT 110.440 198.125 111.335 198.500 ;
        RECT 111.845 198.455 112.235 198.535 ;
        RECT 113.555 198.485 114.075 199.025 ;
        RECT 114.720 198.705 115.395 198.955 ;
        RECT 115.615 198.705 115.955 198.955 ;
        RECT 116.125 198.705 116.415 199.035 ;
        RECT 109.385 197.695 110.270 197.865 ;
        RECT 110.450 197.395 110.765 197.895 ;
        RECT 110.995 197.565 111.335 198.125 ;
        RECT 111.505 197.395 111.675 198.405 ;
        RECT 111.845 197.610 112.175 198.455 ;
        RECT 112.345 197.395 112.515 198.310 ;
        RECT 112.865 197.395 114.075 198.485 ;
        RECT 114.245 197.395 114.535 198.560 ;
        RECT 114.720 198.345 114.985 198.705 ;
        RECT 116.125 198.455 116.295 198.705 ;
        RECT 115.355 198.285 116.295 198.455 ;
        RECT 114.905 197.395 115.185 198.065 ;
        RECT 115.355 197.735 115.655 198.285 ;
        RECT 116.585 198.115 116.835 199.485 ;
        RECT 115.855 197.395 116.185 198.115 ;
        RECT 116.375 197.565 116.835 198.115 ;
        RECT 117.005 199.270 117.265 199.775 ;
        RECT 117.445 199.565 117.775 199.945 ;
        RECT 117.955 199.395 118.125 199.775 ;
        RECT 117.005 198.470 117.175 199.270 ;
        RECT 117.460 199.225 118.125 199.395 ;
        RECT 117.460 198.970 117.630 199.225 ;
        RECT 118.385 199.175 121.895 199.945 ;
        RECT 123.035 199.290 123.365 199.725 ;
        RECT 123.535 199.335 123.705 199.945 ;
        RECT 122.985 199.205 123.365 199.290 ;
        RECT 123.875 199.205 124.205 199.730 ;
        RECT 124.465 199.415 124.675 199.945 ;
        RECT 124.950 199.495 125.735 199.665 ;
        RECT 125.905 199.495 126.310 199.665 ;
        RECT 117.345 198.640 117.630 198.970 ;
        RECT 117.865 198.675 118.195 199.045 ;
        RECT 118.385 198.655 120.035 199.175 ;
        RECT 122.985 199.165 123.210 199.205 ;
        RECT 117.460 198.495 117.630 198.640 ;
        RECT 117.005 197.565 117.275 198.470 ;
        RECT 117.460 198.325 118.125 198.495 ;
        RECT 120.205 198.485 121.895 199.005 ;
        RECT 117.445 197.395 117.775 198.155 ;
        RECT 117.955 197.565 118.125 198.325 ;
        RECT 118.385 197.395 121.895 198.485 ;
        RECT 122.985 198.585 123.155 199.165 ;
        RECT 123.875 199.035 124.075 199.205 ;
        RECT 124.950 199.035 125.120 199.495 ;
        RECT 123.325 198.705 124.075 199.035 ;
        RECT 124.245 198.705 125.120 199.035 ;
        RECT 122.985 198.535 123.200 198.585 ;
        RECT 122.985 198.455 123.375 198.535 ;
        RECT 123.045 197.610 123.375 198.455 ;
        RECT 123.885 198.500 124.075 198.705 ;
        RECT 123.545 197.395 123.715 198.405 ;
        RECT 123.885 198.125 124.780 198.500 ;
        RECT 123.885 197.565 124.225 198.125 ;
        RECT 124.455 197.395 124.770 197.895 ;
        RECT 124.950 197.865 125.120 198.705 ;
        RECT 125.290 198.995 125.755 199.325 ;
        RECT 126.140 199.265 126.310 199.495 ;
        RECT 126.490 199.445 126.860 199.945 ;
        RECT 127.180 199.495 127.855 199.665 ;
        RECT 128.050 199.495 128.385 199.665 ;
        RECT 125.290 198.035 125.610 198.995 ;
        RECT 126.140 198.965 126.970 199.265 ;
        RECT 125.780 198.065 125.970 198.785 ;
        RECT 126.140 197.895 126.310 198.965 ;
        RECT 126.770 198.935 126.970 198.965 ;
        RECT 126.480 198.715 126.650 198.785 ;
        RECT 127.180 198.715 127.350 199.495 ;
        RECT 128.215 199.355 128.385 199.495 ;
        RECT 128.555 199.485 128.805 199.945 ;
        RECT 126.480 198.545 127.350 198.715 ;
        RECT 127.520 199.075 128.045 199.295 ;
        RECT 128.215 199.225 128.440 199.355 ;
        RECT 126.480 198.455 126.990 198.545 ;
        RECT 124.950 197.695 125.835 197.865 ;
        RECT 126.060 197.565 126.310 197.895 ;
        RECT 126.480 197.395 126.650 198.195 ;
        RECT 126.820 197.840 126.990 198.455 ;
        RECT 127.520 198.375 127.690 199.075 ;
        RECT 127.160 198.010 127.690 198.375 ;
        RECT 127.860 198.310 128.100 198.905 ;
        RECT 128.270 198.120 128.440 199.225 ;
        RECT 128.610 198.365 128.890 199.315 ;
        RECT 128.135 197.990 128.440 198.120 ;
        RECT 126.820 197.670 127.925 197.840 ;
        RECT 128.135 197.565 128.385 197.990 ;
        RECT 128.555 197.395 128.820 197.855 ;
        RECT 129.060 197.565 129.245 199.685 ;
        RECT 129.415 199.565 129.745 199.945 ;
        RECT 129.915 199.395 130.085 199.685 ;
        RECT 130.345 199.400 135.690 199.945 ;
        RECT 129.420 199.225 130.085 199.395 ;
        RECT 129.420 198.235 129.650 199.225 ;
        RECT 129.820 198.405 130.170 199.055 ;
        RECT 131.930 198.570 132.270 199.400 ;
        RECT 135.865 199.175 139.375 199.945 ;
        RECT 140.005 199.220 140.295 199.945 ;
        RECT 140.465 199.400 145.810 199.945 ;
        RECT 129.420 198.065 130.085 198.235 ;
        RECT 129.415 197.395 129.745 197.895 ;
        RECT 129.915 197.565 130.085 198.065 ;
        RECT 133.750 197.830 134.100 199.080 ;
        RECT 135.865 198.655 137.515 199.175 ;
        RECT 137.685 198.485 139.375 199.005 ;
        RECT 142.050 198.570 142.390 199.400 ;
        RECT 145.985 199.175 148.575 199.945 ;
        RECT 149.205 199.195 150.415 199.945 ;
        RECT 130.345 197.395 135.690 197.830 ;
        RECT 135.865 197.395 139.375 198.485 ;
        RECT 140.005 197.395 140.295 198.560 ;
        RECT 143.870 197.830 144.220 199.080 ;
        RECT 145.985 198.655 147.195 199.175 ;
        RECT 147.365 198.485 148.575 199.005 ;
        RECT 140.465 197.395 145.810 197.830 ;
        RECT 145.985 197.395 148.575 198.485 ;
        RECT 149.205 198.485 149.725 199.025 ;
        RECT 149.895 198.655 150.415 199.195 ;
        RECT 149.205 197.395 150.415 198.485 ;
        RECT 11.120 197.225 150.500 197.395 ;
        RECT 11.205 196.135 12.415 197.225 ;
        RECT 12.585 196.790 17.930 197.225 ;
        RECT 18.105 196.790 23.450 197.225 ;
        RECT 11.205 195.425 11.725 195.965 ;
        RECT 11.895 195.595 12.415 196.135 ;
        RECT 11.205 194.675 12.415 195.425 ;
        RECT 14.170 195.220 14.510 196.050 ;
        RECT 15.990 195.540 16.340 196.790 ;
        RECT 19.690 195.220 20.030 196.050 ;
        RECT 21.510 195.540 21.860 196.790 ;
        RECT 24.085 196.060 24.375 197.225 ;
        RECT 24.545 196.790 29.890 197.225 ;
        RECT 30.065 196.790 35.410 197.225 ;
        RECT 12.585 194.675 17.930 195.220 ;
        RECT 18.105 194.675 23.450 195.220 ;
        RECT 24.085 194.675 24.375 195.400 ;
        RECT 26.130 195.220 26.470 196.050 ;
        RECT 27.950 195.540 28.300 196.790 ;
        RECT 31.650 195.220 31.990 196.050 ;
        RECT 33.470 195.540 33.820 196.790 ;
        RECT 35.585 196.135 38.175 197.225 ;
        RECT 38.435 196.605 38.605 197.035 ;
        RECT 38.775 196.775 39.105 197.225 ;
        RECT 38.435 196.375 39.110 196.605 ;
        RECT 35.585 195.445 36.795 195.965 ;
        RECT 36.965 195.615 38.175 196.135 ;
        RECT 24.545 194.675 29.890 195.220 ;
        RECT 30.065 194.675 35.410 195.220 ;
        RECT 35.585 194.675 38.175 195.445 ;
        RECT 38.405 195.355 38.705 196.205 ;
        RECT 38.875 195.725 39.110 196.375 ;
        RECT 39.280 196.065 39.565 197.010 ;
        RECT 39.745 196.755 40.430 197.225 ;
        RECT 39.740 196.235 40.435 196.545 ;
        RECT 40.610 196.170 40.915 196.955 ;
        RECT 39.280 195.915 40.140 196.065 ;
        RECT 40.705 196.035 40.915 196.170 ;
        RECT 41.110 196.085 41.365 197.225 ;
        RECT 41.560 196.675 42.755 197.005 ;
        RECT 39.280 195.895 40.565 195.915 ;
        RECT 38.875 195.395 39.410 195.725 ;
        RECT 39.580 195.535 40.565 195.895 ;
        RECT 38.875 195.245 39.095 195.395 ;
        RECT 38.350 194.675 38.685 195.180 ;
        RECT 38.855 194.870 39.095 195.245 ;
        RECT 39.580 195.200 39.750 195.535 ;
        RECT 40.740 195.365 40.915 196.035 ;
        RECT 41.615 195.915 41.785 196.475 ;
        RECT 42.010 196.255 42.430 196.505 ;
        RECT 42.935 196.425 43.215 197.225 ;
        RECT 42.010 196.085 43.255 196.255 ;
        RECT 43.425 196.085 43.695 197.055 ;
        RECT 43.870 196.425 44.125 197.225 ;
        RECT 44.325 196.375 44.655 197.055 ;
        RECT 43.085 195.915 43.255 196.085 ;
        RECT 43.465 196.035 43.695 196.085 ;
        RECT 41.110 195.665 41.445 195.915 ;
        RECT 41.615 195.585 42.355 195.915 ;
        RECT 43.085 195.585 43.315 195.915 ;
        RECT 41.615 195.495 41.865 195.585 ;
        RECT 39.375 195.005 39.750 195.200 ;
        RECT 39.375 194.860 39.545 195.005 ;
        RECT 40.110 194.675 40.505 195.170 ;
        RECT 40.675 194.845 40.915 195.365 ;
        RECT 41.130 195.325 41.865 195.495 ;
        RECT 43.085 195.415 43.255 195.585 ;
        RECT 41.130 194.855 41.440 195.325 ;
        RECT 42.515 195.245 43.255 195.415 ;
        RECT 43.525 195.350 43.695 196.035 ;
        RECT 43.870 195.885 44.115 196.245 ;
        RECT 44.305 196.095 44.655 196.375 ;
        RECT 44.305 195.715 44.475 196.095 ;
        RECT 44.835 195.915 45.030 196.965 ;
        RECT 45.210 196.085 45.530 197.225 ;
        RECT 45.705 196.135 49.215 197.225 ;
        RECT 41.610 194.675 42.345 195.155 ;
        RECT 42.515 194.895 42.685 195.245 ;
        RECT 42.855 194.675 43.235 195.075 ;
        RECT 43.425 195.005 43.695 195.350 ;
        RECT 43.955 195.545 44.475 195.715 ;
        RECT 44.645 195.585 45.030 195.915 ;
        RECT 45.210 195.865 45.470 195.915 ;
        RECT 45.210 195.695 45.475 195.865 ;
        RECT 45.210 195.585 45.470 195.695 ;
        RECT 43.955 194.980 44.125 195.545 ;
        RECT 45.705 195.445 47.355 195.965 ;
        RECT 47.525 195.615 49.215 196.135 ;
        RECT 49.845 196.060 50.135 197.225 ;
        RECT 50.305 196.790 55.650 197.225 ;
        RECT 44.315 195.205 45.530 195.375 ;
        RECT 44.315 194.900 44.545 195.205 ;
        RECT 44.715 194.675 45.045 195.035 ;
        RECT 45.240 194.855 45.530 195.205 ;
        RECT 45.705 194.675 49.215 195.445 ;
        RECT 49.845 194.675 50.135 195.400 ;
        RECT 51.890 195.220 52.230 196.050 ;
        RECT 53.710 195.540 54.060 196.790 ;
        RECT 55.825 196.135 57.495 197.225 ;
        RECT 57.665 196.715 57.925 197.225 ;
        RECT 55.825 195.445 56.575 195.965 ;
        RECT 56.745 195.615 57.495 196.135 ;
        RECT 57.665 195.665 58.005 196.545 ;
        RECT 58.175 195.835 58.345 197.055 ;
        RECT 58.585 196.720 59.200 197.225 ;
        RECT 58.585 196.185 58.835 196.550 ;
        RECT 59.005 196.545 59.200 196.720 ;
        RECT 59.370 196.715 59.845 197.055 ;
        RECT 60.015 196.680 60.230 197.225 ;
        RECT 59.005 196.355 59.335 196.545 ;
        RECT 59.555 196.185 60.270 196.480 ;
        RECT 60.440 196.355 60.715 197.055 ;
        RECT 60.975 196.555 61.145 197.055 ;
        RECT 61.315 196.725 61.645 197.225 ;
        RECT 60.975 196.385 61.640 196.555 ;
        RECT 58.585 196.015 60.375 196.185 ;
        RECT 58.175 195.585 58.970 195.835 ;
        RECT 58.175 195.495 58.425 195.585 ;
        RECT 50.305 194.675 55.650 195.220 ;
        RECT 55.825 194.675 57.495 195.445 ;
        RECT 57.665 194.675 57.925 195.495 ;
        RECT 58.095 195.075 58.425 195.495 ;
        RECT 59.140 195.160 59.395 196.015 ;
        RECT 58.605 194.895 59.395 195.160 ;
        RECT 59.565 195.315 59.975 195.835 ;
        RECT 60.145 195.585 60.375 196.015 ;
        RECT 60.545 195.325 60.715 196.355 ;
        RECT 60.890 195.565 61.240 196.215 ;
        RECT 61.410 195.395 61.640 196.385 ;
        RECT 59.565 194.895 59.765 195.315 ;
        RECT 59.955 194.675 60.285 195.135 ;
        RECT 60.455 194.845 60.715 195.325 ;
        RECT 60.975 195.225 61.640 195.395 ;
        RECT 60.975 194.935 61.145 195.225 ;
        RECT 61.315 194.675 61.645 195.055 ;
        RECT 61.815 194.935 62.000 197.055 ;
        RECT 62.240 196.765 62.505 197.225 ;
        RECT 62.675 196.630 62.925 197.055 ;
        RECT 63.135 196.780 64.240 196.950 ;
        RECT 62.620 196.500 62.925 196.630 ;
        RECT 62.170 195.305 62.450 196.255 ;
        RECT 62.620 195.395 62.790 196.500 ;
        RECT 62.960 195.715 63.200 196.310 ;
        RECT 63.370 196.245 63.900 196.610 ;
        RECT 63.370 195.545 63.540 196.245 ;
        RECT 64.070 196.165 64.240 196.780 ;
        RECT 64.410 196.425 64.580 197.225 ;
        RECT 64.750 196.725 65.000 197.055 ;
        RECT 65.225 196.755 66.110 196.925 ;
        RECT 64.070 196.075 64.580 196.165 ;
        RECT 62.620 195.265 62.845 195.395 ;
        RECT 63.015 195.325 63.540 195.545 ;
        RECT 63.710 195.905 64.580 196.075 ;
        RECT 62.255 194.675 62.505 195.135 ;
        RECT 62.675 195.125 62.845 195.265 ;
        RECT 63.710 195.125 63.880 195.905 ;
        RECT 64.410 195.835 64.580 195.905 ;
        RECT 64.090 195.655 64.290 195.685 ;
        RECT 64.750 195.655 64.920 196.725 ;
        RECT 65.090 195.835 65.280 196.555 ;
        RECT 64.090 195.355 64.920 195.655 ;
        RECT 65.450 195.625 65.770 196.585 ;
        RECT 62.675 194.955 63.010 195.125 ;
        RECT 63.205 194.955 63.880 195.125 ;
        RECT 64.200 194.675 64.570 195.175 ;
        RECT 64.750 195.125 64.920 195.355 ;
        RECT 65.305 195.295 65.770 195.625 ;
        RECT 65.940 195.915 66.110 196.755 ;
        RECT 66.290 196.725 66.605 197.225 ;
        RECT 66.835 196.495 67.175 197.055 ;
        RECT 66.280 196.120 67.175 196.495 ;
        RECT 67.345 196.215 67.515 197.225 ;
        RECT 66.985 195.915 67.175 196.120 ;
        RECT 67.685 196.165 68.015 197.010 ;
        RECT 67.685 196.085 68.075 196.165 ;
        RECT 68.245 196.135 69.915 197.225 ;
        RECT 67.860 196.035 68.075 196.085 ;
        RECT 65.940 195.585 66.815 195.915 ;
        RECT 66.985 195.585 67.735 195.915 ;
        RECT 65.940 195.125 66.110 195.585 ;
        RECT 66.985 195.415 67.185 195.585 ;
        RECT 67.905 195.455 68.075 196.035 ;
        RECT 67.850 195.415 68.075 195.455 ;
        RECT 64.750 194.955 65.155 195.125 ;
        RECT 65.325 194.955 66.110 195.125 ;
        RECT 66.385 194.675 66.595 195.205 ;
        RECT 66.855 194.890 67.185 195.415 ;
        RECT 67.695 195.330 68.075 195.415 ;
        RECT 68.245 195.445 68.995 195.965 ;
        RECT 69.165 195.615 69.915 196.135 ;
        RECT 70.085 196.085 70.355 197.055 ;
        RECT 70.565 196.425 70.845 197.225 ;
        RECT 71.025 196.675 72.220 197.005 ;
        RECT 71.350 196.255 71.770 196.505 ;
        RECT 70.525 196.085 71.770 196.255 ;
        RECT 70.085 196.035 70.315 196.085 ;
        RECT 67.355 194.675 67.525 195.285 ;
        RECT 67.695 194.895 68.025 195.330 ;
        RECT 68.245 194.675 69.915 195.445 ;
        RECT 70.085 195.350 70.255 196.035 ;
        RECT 70.525 195.915 70.695 196.085 ;
        RECT 71.995 195.915 72.165 196.475 ;
        RECT 72.415 196.085 72.670 197.225 ;
        RECT 72.845 196.135 75.435 197.225 ;
        RECT 70.465 195.585 70.695 195.915 ;
        RECT 71.425 195.585 72.165 195.915 ;
        RECT 72.335 195.665 72.670 195.915 ;
        RECT 70.525 195.415 70.695 195.585 ;
        RECT 71.915 195.495 72.165 195.585 ;
        RECT 70.085 195.005 70.355 195.350 ;
        RECT 70.525 195.245 71.265 195.415 ;
        RECT 71.915 195.325 72.650 195.495 ;
        RECT 70.545 194.675 70.925 195.075 ;
        RECT 71.095 194.895 71.265 195.245 ;
        RECT 71.435 194.675 72.170 195.155 ;
        RECT 72.340 194.855 72.650 195.325 ;
        RECT 72.845 195.445 74.055 195.965 ;
        RECT 74.225 195.615 75.435 196.135 ;
        RECT 75.605 196.060 75.895 197.225 ;
        RECT 76.065 196.135 77.735 197.225 ;
        RECT 76.065 195.445 76.815 195.965 ;
        RECT 76.985 195.615 77.735 196.135 ;
        RECT 78.090 196.255 78.480 196.430 ;
        RECT 78.965 196.425 79.295 197.225 ;
        RECT 79.465 196.435 80.000 197.055 ;
        RECT 78.090 196.085 79.515 196.255 ;
        RECT 72.845 194.675 75.435 195.445 ;
        RECT 75.605 194.675 75.895 195.400 ;
        RECT 76.065 194.675 77.735 195.445 ;
        RECT 77.965 195.355 78.320 195.915 ;
        RECT 78.490 195.185 78.660 196.085 ;
        RECT 78.830 195.355 79.095 195.915 ;
        RECT 79.345 195.585 79.515 196.085 ;
        RECT 79.685 195.415 80.000 196.435 ;
        RECT 80.390 196.255 80.780 196.430 ;
        RECT 81.265 196.425 81.595 197.225 ;
        RECT 81.765 196.435 82.300 197.055 ;
        RECT 82.505 196.715 82.765 197.225 ;
        RECT 80.390 196.085 81.815 196.255 ;
        RECT 78.070 194.675 78.310 195.185 ;
        RECT 78.490 194.855 78.770 195.185 ;
        RECT 79.000 194.675 79.215 195.185 ;
        RECT 79.385 194.845 80.000 195.415 ;
        RECT 80.265 195.355 80.620 195.915 ;
        RECT 80.790 195.185 80.960 196.085 ;
        RECT 81.130 195.355 81.395 195.915 ;
        RECT 81.645 195.585 81.815 196.085 ;
        RECT 81.985 195.415 82.300 196.435 ;
        RECT 82.505 195.665 82.845 196.545 ;
        RECT 83.015 195.835 83.185 197.055 ;
        RECT 83.425 196.720 84.040 197.225 ;
        RECT 83.425 196.185 83.675 196.550 ;
        RECT 83.845 196.545 84.040 196.720 ;
        RECT 84.210 196.715 84.685 197.055 ;
        RECT 84.855 196.680 85.070 197.225 ;
        RECT 83.845 196.355 84.175 196.545 ;
        RECT 84.395 196.185 85.110 196.480 ;
        RECT 85.280 196.355 85.555 197.055 ;
        RECT 83.425 196.015 85.215 196.185 ;
        RECT 83.015 195.585 83.810 195.835 ;
        RECT 83.015 195.495 83.265 195.585 ;
        RECT 80.370 194.675 80.610 195.185 ;
        RECT 80.790 194.855 81.070 195.185 ;
        RECT 81.300 194.675 81.515 195.185 ;
        RECT 81.685 194.845 82.300 195.415 ;
        RECT 82.505 194.675 82.765 195.495 ;
        RECT 82.935 195.075 83.265 195.495 ;
        RECT 83.980 195.160 84.235 196.015 ;
        RECT 83.445 194.895 84.235 195.160 ;
        RECT 84.405 195.315 84.815 195.835 ;
        RECT 84.985 195.585 85.215 196.015 ;
        RECT 85.385 195.325 85.555 196.355 ;
        RECT 85.725 196.135 87.395 197.225 ;
        RECT 84.405 194.895 84.605 195.315 ;
        RECT 84.795 194.675 85.125 195.135 ;
        RECT 85.295 194.845 85.555 195.325 ;
        RECT 85.725 195.445 86.475 195.965 ;
        RECT 86.645 195.615 87.395 196.135 ;
        RECT 88.115 196.295 88.285 197.055 ;
        RECT 88.465 196.465 88.795 197.225 ;
        RECT 88.115 196.125 88.780 196.295 ;
        RECT 88.965 196.150 89.235 197.055 ;
        RECT 89.495 196.555 89.665 197.055 ;
        RECT 89.835 196.725 90.165 197.225 ;
        RECT 89.495 196.385 90.160 196.555 ;
        RECT 88.610 195.980 88.780 196.125 ;
        RECT 88.045 195.575 88.375 195.945 ;
        RECT 88.610 195.650 88.895 195.980 ;
        RECT 85.725 194.675 87.395 195.445 ;
        RECT 88.610 195.395 88.780 195.650 ;
        RECT 88.115 195.225 88.780 195.395 ;
        RECT 89.065 195.350 89.235 196.150 ;
        RECT 89.410 195.565 89.760 196.215 ;
        RECT 89.930 195.395 90.160 196.385 ;
        RECT 88.115 194.845 88.285 195.225 ;
        RECT 88.465 194.675 88.795 195.055 ;
        RECT 88.975 194.845 89.235 195.350 ;
        RECT 89.495 195.225 90.160 195.395 ;
        RECT 89.495 194.935 89.665 195.225 ;
        RECT 89.835 194.675 90.165 195.055 ;
        RECT 90.335 194.935 90.520 197.055 ;
        RECT 90.760 196.765 91.025 197.225 ;
        RECT 91.195 196.630 91.445 197.055 ;
        RECT 91.655 196.780 92.760 196.950 ;
        RECT 91.140 196.500 91.445 196.630 ;
        RECT 90.690 195.305 90.970 196.255 ;
        RECT 91.140 195.395 91.310 196.500 ;
        RECT 91.480 195.715 91.720 196.310 ;
        RECT 91.890 196.245 92.420 196.610 ;
        RECT 91.890 195.545 92.060 196.245 ;
        RECT 92.590 196.165 92.760 196.780 ;
        RECT 92.930 196.425 93.100 197.225 ;
        RECT 93.270 196.725 93.520 197.055 ;
        RECT 93.745 196.755 94.630 196.925 ;
        RECT 92.590 196.075 93.100 196.165 ;
        RECT 91.140 195.265 91.365 195.395 ;
        RECT 91.535 195.325 92.060 195.545 ;
        RECT 92.230 195.905 93.100 196.075 ;
        RECT 90.775 194.675 91.025 195.135 ;
        RECT 91.195 195.125 91.365 195.265 ;
        RECT 92.230 195.125 92.400 195.905 ;
        RECT 92.930 195.835 93.100 195.905 ;
        RECT 92.610 195.655 92.810 195.685 ;
        RECT 93.270 195.655 93.440 196.725 ;
        RECT 93.610 195.835 93.800 196.555 ;
        RECT 92.610 195.355 93.440 195.655 ;
        RECT 93.970 195.625 94.290 196.585 ;
        RECT 91.195 194.955 91.530 195.125 ;
        RECT 91.725 194.955 92.400 195.125 ;
        RECT 92.720 194.675 93.090 195.175 ;
        RECT 93.270 195.125 93.440 195.355 ;
        RECT 93.825 195.295 94.290 195.625 ;
        RECT 94.460 195.915 94.630 196.755 ;
        RECT 94.810 196.725 95.125 197.225 ;
        RECT 95.355 196.495 95.695 197.055 ;
        RECT 94.800 196.120 95.695 196.495 ;
        RECT 95.865 196.215 96.035 197.225 ;
        RECT 95.505 195.915 95.695 196.120 ;
        RECT 96.205 196.165 96.535 197.010 ;
        RECT 96.705 196.310 96.875 197.225 ;
        RECT 96.205 196.085 96.595 196.165 ;
        RECT 97.225 196.135 100.735 197.225 ;
        RECT 96.380 196.035 96.595 196.085 ;
        RECT 94.460 195.585 95.335 195.915 ;
        RECT 95.505 195.585 96.255 195.915 ;
        RECT 94.460 195.125 94.630 195.585 ;
        RECT 95.505 195.415 95.705 195.585 ;
        RECT 96.425 195.455 96.595 196.035 ;
        RECT 96.370 195.415 96.595 195.455 ;
        RECT 93.270 194.955 93.675 195.125 ;
        RECT 93.845 194.955 94.630 195.125 ;
        RECT 94.905 194.675 95.115 195.205 ;
        RECT 95.375 194.890 95.705 195.415 ;
        RECT 96.215 195.330 96.595 195.415 ;
        RECT 97.225 195.445 98.875 195.965 ;
        RECT 99.045 195.615 100.735 196.135 ;
        RECT 101.365 196.060 101.655 197.225 ;
        RECT 101.825 196.670 102.430 197.225 ;
        RECT 102.605 196.715 103.085 197.055 ;
        RECT 103.255 196.680 103.510 197.225 ;
        RECT 101.825 196.570 102.440 196.670 ;
        RECT 102.255 196.545 102.440 196.570 ;
        RECT 101.825 195.950 102.085 196.400 ;
        RECT 102.255 196.300 102.585 196.545 ;
        RECT 102.755 196.225 103.510 196.475 ;
        RECT 103.680 196.355 103.955 197.055 ;
        RECT 102.740 196.190 103.510 196.225 ;
        RECT 102.725 196.180 103.510 196.190 ;
        RECT 102.720 196.165 103.615 196.180 ;
        RECT 102.700 196.150 103.615 196.165 ;
        RECT 102.680 196.140 103.615 196.150 ;
        RECT 102.655 196.130 103.615 196.140 ;
        RECT 102.585 196.100 103.615 196.130 ;
        RECT 102.565 196.070 103.615 196.100 ;
        RECT 102.545 196.040 103.615 196.070 ;
        RECT 102.515 196.015 103.615 196.040 ;
        RECT 102.480 195.980 103.615 196.015 ;
        RECT 102.450 195.975 103.615 195.980 ;
        RECT 102.450 195.970 102.840 195.975 ;
        RECT 102.450 195.960 102.815 195.970 ;
        RECT 102.450 195.955 102.800 195.960 ;
        RECT 102.450 195.950 102.785 195.955 ;
        RECT 101.825 195.945 102.785 195.950 ;
        RECT 101.825 195.935 102.775 195.945 ;
        RECT 101.825 195.930 102.765 195.935 ;
        RECT 101.825 195.920 102.755 195.930 ;
        RECT 101.825 195.910 102.750 195.920 ;
        RECT 101.825 195.905 102.745 195.910 ;
        RECT 101.825 195.890 102.735 195.905 ;
        RECT 101.825 195.875 102.730 195.890 ;
        RECT 101.825 195.850 102.720 195.875 ;
        RECT 101.825 195.780 102.715 195.850 ;
        RECT 95.875 194.675 96.045 195.285 ;
        RECT 96.215 194.895 96.545 195.330 ;
        RECT 96.715 194.675 96.885 195.190 ;
        RECT 97.225 194.675 100.735 195.445 ;
        RECT 101.365 194.675 101.655 195.400 ;
        RECT 101.825 195.225 102.375 195.610 ;
        RECT 102.545 195.055 102.715 195.780 ;
        RECT 101.825 194.885 102.715 195.055 ;
        RECT 102.885 195.380 103.215 195.805 ;
        RECT 103.385 195.580 103.615 195.975 ;
        RECT 102.885 194.895 103.105 195.380 ;
        RECT 103.785 195.325 103.955 196.355 ;
        RECT 103.275 194.675 103.525 195.215 ;
        RECT 103.695 194.845 103.955 195.325 ;
        RECT 104.160 196.435 104.695 197.055 ;
        RECT 104.160 195.415 104.475 196.435 ;
        RECT 104.865 196.425 105.195 197.225 ;
        RECT 105.680 196.255 106.070 196.430 ;
        RECT 104.645 196.085 106.070 196.255 ;
        RECT 106.425 196.150 106.695 197.055 ;
        RECT 106.865 196.465 107.195 197.225 ;
        RECT 107.375 196.295 107.545 197.055 ;
        RECT 104.645 195.585 104.815 196.085 ;
        RECT 104.160 194.845 104.775 195.415 ;
        RECT 105.065 195.355 105.330 195.915 ;
        RECT 105.500 195.185 105.670 196.085 ;
        RECT 105.840 195.355 106.195 195.915 ;
        RECT 106.425 195.350 106.595 196.150 ;
        RECT 106.880 196.125 107.545 196.295 ;
        RECT 107.805 196.135 111.315 197.225 ;
        RECT 106.880 195.980 107.050 196.125 ;
        RECT 106.765 195.650 107.050 195.980 ;
        RECT 106.880 195.395 107.050 195.650 ;
        RECT 107.285 195.575 107.615 195.945 ;
        RECT 107.805 195.445 109.455 195.965 ;
        RECT 109.625 195.615 111.315 196.135 ;
        RECT 112.405 196.465 112.920 196.875 ;
        RECT 113.155 196.465 113.325 197.225 ;
        RECT 113.495 196.885 115.525 197.055 ;
        RECT 112.405 195.655 112.745 196.465 ;
        RECT 113.495 196.220 113.665 196.885 ;
        RECT 114.060 196.545 115.185 196.715 ;
        RECT 112.915 196.030 113.665 196.220 ;
        RECT 113.835 196.205 114.845 196.375 ;
        RECT 112.405 195.485 113.635 195.655 ;
        RECT 104.945 194.675 105.160 195.185 ;
        RECT 105.390 194.855 105.670 195.185 ;
        RECT 105.850 194.675 106.090 195.185 ;
        RECT 106.425 194.845 106.685 195.350 ;
        RECT 106.880 195.225 107.545 195.395 ;
        RECT 106.865 194.675 107.195 195.055 ;
        RECT 107.375 194.845 107.545 195.225 ;
        RECT 107.805 194.675 111.315 195.445 ;
        RECT 112.680 194.880 112.925 195.485 ;
        RECT 113.145 194.675 113.655 195.210 ;
        RECT 113.835 194.845 114.025 196.205 ;
        RECT 114.195 195.525 114.470 196.005 ;
        RECT 114.195 195.355 114.475 195.525 ;
        RECT 114.675 195.405 114.845 196.205 ;
        RECT 115.015 195.415 115.185 196.545 ;
        RECT 115.355 195.915 115.525 196.885 ;
        RECT 115.695 196.085 115.865 197.225 ;
        RECT 116.035 196.085 116.370 197.055 ;
        RECT 116.545 196.135 120.055 197.225 ;
        RECT 115.355 195.585 115.550 195.915 ;
        RECT 115.775 195.585 116.030 195.915 ;
        RECT 115.775 195.415 115.945 195.585 ;
        RECT 116.200 195.415 116.370 196.085 ;
        RECT 114.195 194.845 114.470 195.355 ;
        RECT 115.015 195.245 115.945 195.415 ;
        RECT 115.015 195.210 115.190 195.245 ;
        RECT 114.660 194.845 115.190 195.210 ;
        RECT 115.615 194.675 115.945 195.075 ;
        RECT 116.115 194.845 116.370 195.415 ;
        RECT 116.545 195.445 118.195 195.965 ;
        RECT 118.365 195.615 120.055 196.135 ;
        RECT 120.230 196.085 120.550 197.225 ;
        RECT 120.730 195.915 120.925 196.965 ;
        RECT 121.105 196.375 121.435 197.055 ;
        RECT 121.635 196.425 121.890 197.225 ;
        RECT 121.105 196.095 121.455 196.375 ;
        RECT 120.290 195.865 120.550 195.915 ;
        RECT 120.285 195.695 120.550 195.865 ;
        RECT 120.290 195.585 120.550 195.695 ;
        RECT 120.730 195.585 121.115 195.915 ;
        RECT 121.285 195.715 121.455 196.095 ;
        RECT 121.645 195.885 121.890 196.245 ;
        RECT 122.065 196.135 125.575 197.225 ;
        RECT 125.745 196.135 126.955 197.225 ;
        RECT 121.285 195.545 121.805 195.715 ;
        RECT 116.545 194.675 120.055 195.445 ;
        RECT 120.230 195.205 121.445 195.375 ;
        RECT 120.230 194.855 120.520 195.205 ;
        RECT 120.715 194.675 121.045 195.035 ;
        RECT 121.215 194.900 121.445 195.205 ;
        RECT 121.635 195.185 121.805 195.545 ;
        RECT 122.065 195.445 123.715 195.965 ;
        RECT 123.885 195.615 125.575 196.135 ;
        RECT 121.635 195.015 121.835 195.185 ;
        RECT 121.635 194.980 121.805 195.015 ;
        RECT 122.065 194.675 125.575 195.445 ;
        RECT 125.745 195.425 126.265 195.965 ;
        RECT 126.435 195.595 126.955 196.135 ;
        RECT 127.125 196.060 127.415 197.225 ;
        RECT 127.585 196.790 132.930 197.225 ;
        RECT 133.105 196.790 138.450 197.225 ;
        RECT 138.625 196.790 143.970 197.225 ;
        RECT 125.745 194.675 126.955 195.425 ;
        RECT 127.125 194.675 127.415 195.400 ;
        RECT 129.170 195.220 129.510 196.050 ;
        RECT 130.990 195.540 131.340 196.790 ;
        RECT 134.690 195.220 135.030 196.050 ;
        RECT 136.510 195.540 136.860 196.790 ;
        RECT 140.210 195.220 140.550 196.050 ;
        RECT 142.030 195.540 142.380 196.790 ;
        RECT 144.145 196.135 147.655 197.225 ;
        RECT 147.825 196.135 149.035 197.225 ;
        RECT 144.145 195.445 145.795 195.965 ;
        RECT 145.965 195.615 147.655 196.135 ;
        RECT 127.585 194.675 132.930 195.220 ;
        RECT 133.105 194.675 138.450 195.220 ;
        RECT 138.625 194.675 143.970 195.220 ;
        RECT 144.145 194.675 147.655 195.445 ;
        RECT 147.825 195.425 148.345 195.965 ;
        RECT 148.515 195.595 149.035 196.135 ;
        RECT 149.205 196.135 150.415 197.225 ;
        RECT 149.205 195.595 149.725 196.135 ;
        RECT 149.895 195.425 150.415 195.965 ;
        RECT 147.825 194.675 149.035 195.425 ;
        RECT 149.205 194.675 150.415 195.425 ;
        RECT 11.120 194.505 150.500 194.675 ;
        RECT 11.205 193.755 12.415 194.505 ;
        RECT 12.585 193.755 13.795 194.505 ;
        RECT 13.965 193.830 14.225 194.335 ;
        RECT 14.405 194.125 14.735 194.505 ;
        RECT 14.915 193.955 15.085 194.335 ;
        RECT 11.205 193.215 11.725 193.755 ;
        RECT 11.895 193.045 12.415 193.585 ;
        RECT 12.585 193.215 13.105 193.755 ;
        RECT 13.275 193.045 13.795 193.585 ;
        RECT 11.205 191.955 12.415 193.045 ;
        RECT 12.585 191.955 13.795 193.045 ;
        RECT 13.965 193.030 14.135 193.830 ;
        RECT 14.420 193.785 15.085 193.955 ;
        RECT 15.895 193.955 16.065 194.245 ;
        RECT 16.235 194.125 16.565 194.505 ;
        RECT 15.895 193.785 16.560 193.955 ;
        RECT 14.420 193.530 14.590 193.785 ;
        RECT 14.305 193.200 14.590 193.530 ;
        RECT 14.825 193.235 15.155 193.605 ;
        RECT 14.420 193.055 14.590 193.200 ;
        RECT 13.965 192.125 14.235 193.030 ;
        RECT 14.420 192.885 15.085 193.055 ;
        RECT 15.810 192.965 16.160 193.615 ;
        RECT 14.405 191.955 14.735 192.715 ;
        RECT 14.915 192.125 15.085 192.885 ;
        RECT 16.330 192.795 16.560 193.785 ;
        RECT 15.895 192.625 16.560 192.795 ;
        RECT 15.895 192.125 16.065 192.625 ;
        RECT 16.235 191.955 16.565 192.455 ;
        RECT 16.735 192.125 16.920 194.245 ;
        RECT 17.175 194.045 17.425 194.505 ;
        RECT 17.595 194.055 17.930 194.225 ;
        RECT 18.125 194.055 18.800 194.225 ;
        RECT 17.595 193.915 17.765 194.055 ;
        RECT 17.090 192.925 17.370 193.875 ;
        RECT 17.540 193.785 17.765 193.915 ;
        RECT 17.540 192.680 17.710 193.785 ;
        RECT 17.935 193.635 18.460 193.855 ;
        RECT 17.880 192.870 18.120 193.465 ;
        RECT 18.290 192.935 18.460 193.635 ;
        RECT 18.630 193.275 18.800 194.055 ;
        RECT 19.120 194.005 19.490 194.505 ;
        RECT 19.670 194.055 20.075 194.225 ;
        RECT 20.245 194.055 21.030 194.225 ;
        RECT 19.670 193.825 19.840 194.055 ;
        RECT 19.010 193.525 19.840 193.825 ;
        RECT 20.225 193.555 20.690 193.885 ;
        RECT 19.010 193.495 19.210 193.525 ;
        RECT 19.330 193.275 19.500 193.345 ;
        RECT 18.630 193.105 19.500 193.275 ;
        RECT 18.990 193.015 19.500 193.105 ;
        RECT 17.540 192.550 17.845 192.680 ;
        RECT 18.290 192.570 18.820 192.935 ;
        RECT 17.160 191.955 17.425 192.415 ;
        RECT 17.595 192.125 17.845 192.550 ;
        RECT 18.990 192.400 19.160 193.015 ;
        RECT 18.055 192.230 19.160 192.400 ;
        RECT 19.330 191.955 19.500 192.755 ;
        RECT 19.670 192.455 19.840 193.525 ;
        RECT 20.010 192.625 20.200 193.345 ;
        RECT 20.370 192.595 20.690 193.555 ;
        RECT 20.860 193.595 21.030 194.055 ;
        RECT 21.305 193.975 21.515 194.505 ;
        RECT 21.775 193.765 22.105 194.290 ;
        RECT 22.275 193.895 22.445 194.505 ;
        RECT 22.615 193.850 22.945 194.285 ;
        RECT 23.255 193.955 23.425 194.245 ;
        RECT 23.595 194.125 23.925 194.505 ;
        RECT 22.615 193.765 22.995 193.850 ;
        RECT 23.255 193.785 23.920 193.955 ;
        RECT 21.905 193.595 22.105 193.765 ;
        RECT 22.770 193.725 22.995 193.765 ;
        RECT 20.860 193.265 21.735 193.595 ;
        RECT 21.905 193.265 22.655 193.595 ;
        RECT 19.670 192.125 19.920 192.455 ;
        RECT 20.860 192.425 21.030 193.265 ;
        RECT 21.905 193.060 22.095 193.265 ;
        RECT 22.825 193.145 22.995 193.725 ;
        RECT 22.780 193.095 22.995 193.145 ;
        RECT 21.200 192.685 22.095 193.060 ;
        RECT 22.605 193.015 22.995 193.095 ;
        RECT 20.145 192.255 21.030 192.425 ;
        RECT 21.210 191.955 21.525 192.455 ;
        RECT 21.755 192.125 22.095 192.685 ;
        RECT 22.265 191.955 22.435 192.965 ;
        RECT 22.605 192.170 22.935 193.015 ;
        RECT 23.170 192.965 23.520 193.615 ;
        RECT 23.690 192.795 23.920 193.785 ;
        RECT 23.255 192.625 23.920 192.795 ;
        RECT 23.255 192.125 23.425 192.625 ;
        RECT 23.595 191.955 23.925 192.455 ;
        RECT 24.095 192.125 24.280 194.245 ;
        RECT 24.535 194.045 24.785 194.505 ;
        RECT 24.955 194.055 25.290 194.225 ;
        RECT 25.485 194.055 26.160 194.225 ;
        RECT 24.955 193.915 25.125 194.055 ;
        RECT 24.450 192.925 24.730 193.875 ;
        RECT 24.900 193.785 25.125 193.915 ;
        RECT 24.900 192.680 25.070 193.785 ;
        RECT 25.295 193.635 25.820 193.855 ;
        RECT 25.240 192.870 25.480 193.465 ;
        RECT 25.650 192.935 25.820 193.635 ;
        RECT 25.990 193.275 26.160 194.055 ;
        RECT 26.480 194.005 26.850 194.505 ;
        RECT 27.030 194.055 27.435 194.225 ;
        RECT 27.605 194.055 28.390 194.225 ;
        RECT 27.030 193.825 27.200 194.055 ;
        RECT 26.370 193.525 27.200 193.825 ;
        RECT 27.585 193.555 28.050 193.885 ;
        RECT 26.370 193.495 26.570 193.525 ;
        RECT 26.690 193.275 26.860 193.345 ;
        RECT 25.990 193.105 26.860 193.275 ;
        RECT 26.350 193.015 26.860 193.105 ;
        RECT 24.900 192.550 25.205 192.680 ;
        RECT 25.650 192.570 26.180 192.935 ;
        RECT 24.520 191.955 24.785 192.415 ;
        RECT 24.955 192.125 25.205 192.550 ;
        RECT 26.350 192.400 26.520 193.015 ;
        RECT 25.415 192.230 26.520 192.400 ;
        RECT 26.690 191.955 26.860 192.755 ;
        RECT 27.030 192.455 27.200 193.525 ;
        RECT 27.370 192.625 27.560 193.345 ;
        RECT 27.730 192.595 28.050 193.555 ;
        RECT 28.220 193.595 28.390 194.055 ;
        RECT 28.665 193.975 28.875 194.505 ;
        RECT 29.135 193.765 29.465 194.290 ;
        RECT 29.635 193.895 29.805 194.505 ;
        RECT 29.975 193.850 30.305 194.285 ;
        RECT 30.615 194.005 31.110 194.335 ;
        RECT 29.975 193.765 30.355 193.850 ;
        RECT 29.265 193.595 29.465 193.765 ;
        RECT 30.130 193.725 30.355 193.765 ;
        RECT 28.220 193.265 29.095 193.595 ;
        RECT 29.265 193.265 30.015 193.595 ;
        RECT 27.030 192.125 27.280 192.455 ;
        RECT 28.220 192.425 28.390 193.265 ;
        RECT 29.265 193.060 29.455 193.265 ;
        RECT 30.185 193.145 30.355 193.725 ;
        RECT 30.140 193.095 30.355 193.145 ;
        RECT 28.560 192.685 29.455 193.060 ;
        RECT 29.965 193.015 30.355 193.095 ;
        RECT 27.505 192.255 28.390 192.425 ;
        RECT 28.570 191.955 28.885 192.455 ;
        RECT 29.115 192.125 29.455 192.685 ;
        RECT 29.625 191.955 29.795 192.965 ;
        RECT 29.965 192.170 30.295 193.015 ;
        RECT 30.565 192.515 30.770 193.835 ;
        RECT 30.940 193.095 31.110 194.005 ;
        RECT 31.330 193.265 31.685 194.170 ;
        RECT 31.860 193.285 32.160 194.175 ;
        RECT 31.860 193.265 32.030 193.285 ;
        RECT 32.340 193.265 32.600 194.175 ;
        RECT 32.770 193.700 33.005 194.505 ;
        RECT 33.175 194.250 33.505 194.295 ;
        RECT 33.175 193.785 33.510 194.250 ;
        RECT 32.770 193.275 33.165 193.515 ;
        RECT 32.770 193.095 32.995 193.275 ;
        RECT 33.335 193.095 33.510 193.785 ;
        RECT 33.695 193.780 34.025 194.505 ;
        RECT 34.295 193.955 34.465 194.335 ;
        RECT 34.680 194.125 35.010 194.505 ;
        RECT 34.295 193.785 35.010 193.955 ;
        RECT 34.205 193.235 34.560 193.605 ;
        RECT 34.840 193.595 35.010 193.785 ;
        RECT 35.180 193.760 35.435 194.335 ;
        RECT 34.840 193.265 35.095 193.595 ;
        RECT 30.940 192.925 32.995 193.095 ;
        RECT 30.535 191.955 30.865 192.335 ;
        RECT 31.040 192.125 31.290 192.925 ;
        RECT 31.510 191.955 31.840 192.675 ;
        RECT 32.025 192.125 32.275 192.925 ;
        RECT 32.675 191.955 33.005 192.755 ;
        RECT 33.175 192.465 33.510 193.095 ;
        RECT 34.840 193.055 35.010 193.265 ;
        RECT 34.295 192.885 35.010 193.055 ;
        RECT 35.265 193.030 35.435 193.760 ;
        RECT 35.610 193.665 35.870 194.505 ;
        RECT 36.965 193.780 37.255 194.505 ;
        RECT 37.435 193.780 37.765 194.290 ;
        RECT 37.935 194.105 38.265 194.505 ;
        RECT 39.315 193.935 39.645 194.275 ;
        RECT 39.815 194.105 40.145 194.505 ;
        RECT 33.175 192.295 33.515 192.465 ;
        RECT 33.175 192.125 33.510 192.295 ;
        RECT 33.685 191.955 34.015 192.755 ;
        RECT 34.295 192.125 34.465 192.885 ;
        RECT 34.680 191.955 35.010 192.715 ;
        RECT 35.180 192.125 35.435 193.030 ;
        RECT 35.610 191.955 35.870 193.105 ;
        RECT 36.965 191.955 37.255 193.120 ;
        RECT 37.435 193.015 37.625 193.780 ;
        RECT 37.935 193.765 40.300 193.935 ;
        RECT 37.935 193.595 38.105 193.765 ;
        RECT 37.795 193.265 38.105 193.595 ;
        RECT 38.275 193.265 38.580 193.595 ;
        RECT 37.435 192.165 37.765 193.015 ;
        RECT 37.935 191.955 38.185 193.095 ;
        RECT 38.365 192.935 38.580 193.265 ;
        RECT 38.755 192.935 39.040 193.595 ;
        RECT 39.235 192.935 39.500 193.595 ;
        RECT 39.715 192.935 39.960 193.595 ;
        RECT 40.130 192.765 40.300 193.765 ;
        RECT 38.375 192.595 39.665 192.765 ;
        RECT 38.375 192.175 38.625 192.595 ;
        RECT 38.855 191.955 39.185 192.425 ;
        RECT 39.415 192.175 39.665 192.595 ;
        RECT 39.845 192.595 40.300 192.765 ;
        RECT 40.665 193.815 40.905 194.335 ;
        RECT 41.075 194.010 41.470 194.505 ;
        RECT 42.035 194.175 42.205 194.320 ;
        RECT 41.830 193.980 42.205 194.175 ;
        RECT 40.665 193.010 40.840 193.815 ;
        RECT 41.830 193.645 42.000 193.980 ;
        RECT 42.485 193.935 42.725 194.310 ;
        RECT 42.895 194.000 43.230 194.505 ;
        RECT 43.915 194.115 44.245 194.505 ;
        RECT 44.415 193.935 44.585 194.255 ;
        RECT 44.755 194.115 45.085 194.505 ;
        RECT 45.500 194.105 46.455 194.275 ;
        RECT 42.485 193.785 42.705 193.935 ;
        RECT 41.015 193.285 42.000 193.645 ;
        RECT 42.170 193.455 42.705 193.785 ;
        RECT 41.015 193.265 42.300 193.285 ;
        RECT 41.440 193.115 42.300 193.265 ;
        RECT 39.845 192.165 40.175 192.595 ;
        RECT 40.665 192.225 40.970 193.010 ;
        RECT 41.145 192.635 41.840 192.945 ;
        RECT 41.150 191.955 41.835 192.425 ;
        RECT 42.015 192.170 42.300 193.115 ;
        RECT 42.470 192.805 42.705 193.455 ;
        RECT 42.875 192.975 43.175 193.825 ;
        RECT 43.865 193.765 46.115 193.935 ;
        RECT 43.865 192.805 44.035 193.765 ;
        RECT 44.205 193.145 44.450 193.595 ;
        RECT 44.620 193.315 45.170 193.515 ;
        RECT 45.340 193.345 45.715 193.515 ;
        RECT 45.340 193.145 45.510 193.345 ;
        RECT 45.885 193.265 46.115 193.765 ;
        RECT 44.205 192.975 45.510 193.145 ;
        RECT 46.285 193.225 46.455 194.105 ;
        RECT 46.625 193.670 46.915 194.505 ;
        RECT 47.085 193.765 47.550 194.310 ;
        RECT 46.285 193.055 46.915 193.225 ;
        RECT 42.470 192.575 43.145 192.805 ;
        RECT 42.475 191.955 42.805 192.405 ;
        RECT 42.975 192.145 43.145 192.575 ;
        RECT 43.865 192.125 44.245 192.805 ;
        RECT 44.835 191.955 45.005 192.805 ;
        RECT 45.175 192.635 46.415 192.805 ;
        RECT 45.175 192.125 45.505 192.635 ;
        RECT 45.675 191.955 45.845 192.465 ;
        RECT 46.015 192.125 46.415 192.635 ;
        RECT 46.595 192.125 46.915 193.055 ;
        RECT 47.085 192.805 47.255 193.765 ;
        RECT 48.055 193.685 48.225 194.505 ;
        RECT 48.395 193.855 48.725 194.335 ;
        RECT 48.895 194.115 49.245 194.505 ;
        RECT 49.415 193.935 49.645 194.335 ;
        RECT 49.135 193.855 49.645 193.935 ;
        RECT 48.395 193.765 49.645 193.855 ;
        RECT 49.815 193.765 50.135 194.245 ;
        RECT 48.395 193.685 49.305 193.765 ;
        RECT 47.425 193.145 47.670 193.595 ;
        RECT 47.930 193.315 48.625 193.515 ;
        RECT 48.795 193.345 49.395 193.515 ;
        RECT 48.795 193.145 48.965 193.345 ;
        RECT 49.625 193.175 49.795 193.595 ;
        RECT 47.425 192.975 48.965 193.145 ;
        RECT 49.135 193.005 49.795 193.175 ;
        RECT 49.135 192.805 49.305 193.005 ;
        RECT 49.965 192.835 50.135 193.765 ;
        RECT 50.305 193.735 52.895 194.505 ;
        RECT 53.525 193.830 53.795 194.175 ;
        RECT 53.985 194.105 54.365 194.505 ;
        RECT 54.535 193.935 54.705 194.285 ;
        RECT 54.875 194.025 55.610 194.505 ;
        RECT 50.305 193.215 51.515 193.735 ;
        RECT 51.685 193.045 52.895 193.565 ;
        RECT 47.085 192.635 49.305 192.805 ;
        RECT 49.475 192.635 50.135 192.835 ;
        RECT 47.085 191.955 47.385 192.465 ;
        RECT 47.555 192.125 47.885 192.635 ;
        RECT 49.475 192.465 49.645 192.635 ;
        RECT 48.055 191.955 48.685 192.465 ;
        RECT 49.265 192.295 49.645 192.465 ;
        RECT 49.815 191.955 50.115 192.465 ;
        RECT 50.305 191.955 52.895 193.045 ;
        RECT 53.525 193.095 53.695 193.830 ;
        RECT 53.965 193.765 54.705 193.935 ;
        RECT 55.780 193.855 56.090 194.325 ;
        RECT 53.965 193.595 54.135 193.765 ;
        RECT 55.355 193.685 56.090 193.855 ;
        RECT 56.285 193.855 56.545 194.335 ;
        RECT 56.715 193.965 56.965 194.505 ;
        RECT 55.355 193.595 55.605 193.685 ;
        RECT 53.905 193.265 54.135 193.595 ;
        RECT 54.865 193.265 55.605 193.595 ;
        RECT 55.775 193.265 56.110 193.515 ;
        RECT 53.965 193.095 54.135 193.265 ;
        RECT 53.525 192.125 53.795 193.095 ;
        RECT 53.965 192.925 55.210 193.095 ;
        RECT 54.005 191.955 54.285 192.755 ;
        RECT 54.790 192.675 55.210 192.925 ;
        RECT 55.435 192.705 55.605 193.265 ;
        RECT 54.465 192.175 55.660 192.505 ;
        RECT 55.855 191.955 56.110 193.095 ;
        RECT 56.285 192.825 56.455 193.855 ;
        RECT 57.135 193.800 57.355 194.285 ;
        RECT 56.625 193.205 56.855 193.600 ;
        RECT 57.025 193.375 57.355 193.800 ;
        RECT 57.525 194.125 58.415 194.295 ;
        RECT 57.525 193.400 57.695 194.125 ;
        RECT 57.865 193.570 58.415 193.955 ;
        RECT 58.585 193.735 60.255 194.505 ;
        RECT 60.975 193.955 61.145 194.335 ;
        RECT 61.325 194.125 61.655 194.505 ;
        RECT 60.975 193.785 61.640 193.955 ;
        RECT 61.835 193.830 62.095 194.335 ;
        RECT 57.525 193.330 58.415 193.400 ;
        RECT 57.520 193.305 58.415 193.330 ;
        RECT 57.510 193.290 58.415 193.305 ;
        RECT 57.505 193.275 58.415 193.290 ;
        RECT 57.495 193.270 58.415 193.275 ;
        RECT 57.490 193.260 58.415 193.270 ;
        RECT 57.485 193.250 58.415 193.260 ;
        RECT 57.475 193.245 58.415 193.250 ;
        RECT 57.465 193.235 58.415 193.245 ;
        RECT 57.455 193.230 58.415 193.235 ;
        RECT 57.455 193.225 57.790 193.230 ;
        RECT 57.440 193.220 57.790 193.225 ;
        RECT 57.425 193.210 57.790 193.220 ;
        RECT 57.400 193.205 57.790 193.210 ;
        RECT 56.625 193.200 57.790 193.205 ;
        RECT 56.625 193.165 57.760 193.200 ;
        RECT 56.625 193.140 57.725 193.165 ;
        RECT 56.625 193.110 57.695 193.140 ;
        RECT 56.625 193.080 57.675 193.110 ;
        RECT 56.625 193.050 57.655 193.080 ;
        RECT 56.625 193.040 57.585 193.050 ;
        RECT 56.625 193.030 57.560 193.040 ;
        RECT 56.625 193.015 57.540 193.030 ;
        RECT 56.625 193.000 57.520 193.015 ;
        RECT 56.730 192.990 57.515 193.000 ;
        RECT 56.730 192.955 57.500 192.990 ;
        RECT 56.285 192.125 56.560 192.825 ;
        RECT 56.730 192.705 57.485 192.955 ;
        RECT 57.655 192.635 57.985 192.880 ;
        RECT 58.155 192.780 58.415 193.230 ;
        RECT 58.585 193.215 59.335 193.735 ;
        RECT 59.505 193.045 60.255 193.565 ;
        RECT 60.905 193.235 61.235 193.605 ;
        RECT 61.470 193.530 61.640 193.785 ;
        RECT 61.470 193.200 61.755 193.530 ;
        RECT 61.470 193.055 61.640 193.200 ;
        RECT 57.800 192.610 57.985 192.635 ;
        RECT 57.800 192.510 58.415 192.610 ;
        RECT 56.730 191.955 56.985 192.500 ;
        RECT 57.155 192.125 57.635 192.465 ;
        RECT 57.810 191.955 58.415 192.510 ;
        RECT 58.585 191.955 60.255 193.045 ;
        RECT 60.975 192.885 61.640 193.055 ;
        RECT 61.925 193.030 62.095 193.830 ;
        RECT 62.725 193.780 63.015 194.505 ;
        RECT 63.195 193.780 63.525 194.290 ;
        RECT 63.695 194.105 64.025 194.505 ;
        RECT 65.075 193.935 65.405 194.275 ;
        RECT 65.575 194.105 65.905 194.505 ;
        RECT 60.975 192.125 61.145 192.885 ;
        RECT 61.325 191.955 61.655 192.715 ;
        RECT 61.825 192.125 62.095 193.030 ;
        RECT 62.725 191.955 63.015 193.120 ;
        RECT 63.195 193.015 63.385 193.780 ;
        RECT 63.695 193.765 66.060 193.935 ;
        RECT 63.695 193.595 63.865 193.765 ;
        RECT 63.555 193.265 63.865 193.595 ;
        RECT 64.035 193.265 64.340 193.595 ;
        RECT 63.195 192.165 63.525 193.015 ;
        RECT 63.695 191.955 63.945 193.095 ;
        RECT 64.125 192.935 64.340 193.265 ;
        RECT 64.515 192.935 64.800 193.595 ;
        RECT 64.995 192.935 65.260 193.595 ;
        RECT 65.475 192.935 65.720 193.595 ;
        RECT 65.890 192.765 66.060 193.765 ;
        RECT 66.415 193.695 66.685 194.505 ;
        RECT 66.855 193.695 67.185 194.335 ;
        RECT 67.355 193.695 67.595 194.505 ;
        RECT 67.785 193.735 69.455 194.505 ;
        RECT 66.405 193.265 66.755 193.515 ;
        RECT 66.925 193.095 67.095 193.695 ;
        RECT 67.265 193.265 67.615 193.515 ;
        RECT 67.785 193.215 68.535 193.735 ;
        RECT 70.145 193.685 70.355 194.505 ;
        RECT 70.525 193.705 70.855 194.335 ;
        RECT 64.135 192.595 65.425 192.765 ;
        RECT 64.135 192.175 64.385 192.595 ;
        RECT 64.615 191.955 64.945 192.425 ;
        RECT 65.175 192.175 65.425 192.595 ;
        RECT 65.605 192.595 66.060 192.765 ;
        RECT 65.605 192.165 65.935 192.595 ;
        RECT 66.415 191.955 66.745 193.095 ;
        RECT 66.925 192.925 67.605 193.095 ;
        RECT 68.705 193.045 69.455 193.565 ;
        RECT 70.525 193.105 70.775 193.705 ;
        RECT 71.025 193.685 71.255 194.505 ;
        RECT 71.465 193.960 76.810 194.505 ;
        RECT 70.945 193.265 71.275 193.515 ;
        RECT 73.050 193.130 73.390 193.960 ;
        RECT 77.185 193.875 77.515 194.235 ;
        RECT 78.135 194.045 78.385 194.505 ;
        RECT 78.555 194.045 79.115 194.335 ;
        RECT 77.185 193.685 78.575 193.875 ;
        RECT 67.275 192.140 67.605 192.925 ;
        RECT 67.785 191.955 69.455 193.045 ;
        RECT 70.145 191.955 70.355 193.095 ;
        RECT 70.525 192.125 70.855 193.105 ;
        RECT 71.025 191.955 71.255 193.095 ;
        RECT 74.870 192.390 75.220 193.640 ;
        RECT 78.405 193.595 78.575 193.685 ;
        RECT 77.000 193.265 77.675 193.515 ;
        RECT 77.895 193.265 78.235 193.515 ;
        RECT 78.405 193.265 78.695 193.595 ;
        RECT 77.000 192.905 77.265 193.265 ;
        RECT 78.405 193.015 78.575 193.265 ;
        RECT 77.635 192.845 78.575 193.015 ;
        RECT 71.465 191.955 76.810 192.390 ;
        RECT 77.185 191.955 77.465 192.625 ;
        RECT 77.635 192.295 77.935 192.845 ;
        RECT 78.865 192.675 79.115 194.045 ;
        RECT 79.745 193.685 80.005 194.505 ;
        RECT 80.175 193.685 80.505 194.105 ;
        RECT 80.685 194.020 81.475 194.285 ;
        RECT 80.255 193.595 80.505 193.685 ;
        RECT 78.135 191.955 78.465 192.675 ;
        RECT 78.655 192.125 79.115 192.675 ;
        RECT 79.745 192.635 80.085 193.515 ;
        RECT 80.255 193.345 81.050 193.595 ;
        RECT 79.745 191.955 80.005 192.465 ;
        RECT 80.255 192.125 80.425 193.345 ;
        RECT 81.220 193.165 81.475 194.020 ;
        RECT 81.645 193.865 81.845 194.285 ;
        RECT 82.035 194.045 82.365 194.505 ;
        RECT 81.645 193.345 82.055 193.865 ;
        RECT 82.535 193.855 82.795 194.335 ;
        RECT 82.225 193.165 82.455 193.595 ;
        RECT 80.665 192.995 82.455 193.165 ;
        RECT 80.665 192.630 80.915 192.995 ;
        RECT 81.085 192.635 81.415 192.825 ;
        RECT 81.635 192.700 82.350 192.995 ;
        RECT 82.625 192.825 82.795 193.855 ;
        RECT 82.965 193.755 84.175 194.505 ;
        RECT 84.435 193.955 84.605 194.335 ;
        RECT 84.785 194.125 85.115 194.505 ;
        RECT 84.435 193.785 85.100 193.955 ;
        RECT 85.295 193.830 85.555 194.335 ;
        RECT 82.965 193.215 83.485 193.755 ;
        RECT 83.655 193.045 84.175 193.585 ;
        RECT 84.365 193.235 84.695 193.605 ;
        RECT 84.930 193.530 85.100 193.785 ;
        RECT 84.930 193.200 85.215 193.530 ;
        RECT 84.930 193.055 85.100 193.200 ;
        RECT 81.085 192.460 81.280 192.635 ;
        RECT 80.665 191.955 81.280 192.460 ;
        RECT 81.450 192.125 81.925 192.465 ;
        RECT 82.095 191.955 82.310 192.500 ;
        RECT 82.520 192.125 82.795 192.825 ;
        RECT 82.965 191.955 84.175 193.045 ;
        RECT 84.435 192.885 85.100 193.055 ;
        RECT 85.385 193.030 85.555 193.830 ;
        RECT 85.725 193.735 88.315 194.505 ;
        RECT 88.485 193.780 88.775 194.505 ;
        RECT 89.035 193.955 89.205 194.245 ;
        RECT 89.375 194.125 89.705 194.505 ;
        RECT 89.035 193.785 89.700 193.955 ;
        RECT 85.725 193.215 86.935 193.735 ;
        RECT 87.105 193.045 88.315 193.565 ;
        RECT 84.435 192.125 84.605 192.885 ;
        RECT 84.785 191.955 85.115 192.715 ;
        RECT 85.285 192.125 85.555 193.030 ;
        RECT 85.725 191.955 88.315 193.045 ;
        RECT 88.485 191.955 88.775 193.120 ;
        RECT 88.950 192.965 89.300 193.615 ;
        RECT 89.470 192.795 89.700 193.785 ;
        RECT 89.035 192.625 89.700 192.795 ;
        RECT 89.035 192.125 89.205 192.625 ;
        RECT 89.375 191.955 89.705 192.455 ;
        RECT 89.875 192.125 90.060 194.245 ;
        RECT 90.315 194.045 90.565 194.505 ;
        RECT 90.735 194.055 91.070 194.225 ;
        RECT 91.265 194.055 91.940 194.225 ;
        RECT 90.735 193.915 90.905 194.055 ;
        RECT 90.230 192.925 90.510 193.875 ;
        RECT 90.680 193.785 90.905 193.915 ;
        RECT 90.680 192.680 90.850 193.785 ;
        RECT 91.075 193.635 91.600 193.855 ;
        RECT 91.020 192.870 91.260 193.465 ;
        RECT 91.430 192.935 91.600 193.635 ;
        RECT 91.770 193.275 91.940 194.055 ;
        RECT 92.260 194.005 92.630 194.505 ;
        RECT 92.810 194.055 93.215 194.225 ;
        RECT 93.385 194.055 94.170 194.225 ;
        RECT 92.810 193.825 92.980 194.055 ;
        RECT 92.150 193.525 92.980 193.825 ;
        RECT 93.365 193.555 93.830 193.885 ;
        RECT 92.150 193.495 92.350 193.525 ;
        RECT 92.470 193.275 92.640 193.345 ;
        RECT 91.770 193.105 92.640 193.275 ;
        RECT 92.130 193.015 92.640 193.105 ;
        RECT 90.680 192.550 90.985 192.680 ;
        RECT 91.430 192.570 91.960 192.935 ;
        RECT 90.300 191.955 90.565 192.415 ;
        RECT 90.735 192.125 90.985 192.550 ;
        RECT 92.130 192.400 92.300 193.015 ;
        RECT 91.195 192.230 92.300 192.400 ;
        RECT 92.470 191.955 92.640 192.755 ;
        RECT 92.810 192.455 92.980 193.525 ;
        RECT 93.150 192.625 93.340 193.345 ;
        RECT 93.510 192.595 93.830 193.555 ;
        RECT 94.000 193.595 94.170 194.055 ;
        RECT 94.445 193.975 94.655 194.505 ;
        RECT 94.915 193.765 95.245 194.290 ;
        RECT 95.415 193.895 95.585 194.505 ;
        RECT 95.755 193.850 96.085 194.285 ;
        RECT 96.255 193.990 96.425 194.505 ;
        RECT 95.755 193.765 96.135 193.850 ;
        RECT 95.045 193.595 95.245 193.765 ;
        RECT 95.910 193.725 96.135 193.765 ;
        RECT 94.000 193.265 94.875 193.595 ;
        RECT 95.045 193.265 95.795 193.595 ;
        RECT 92.810 192.125 93.060 192.455 ;
        RECT 94.000 192.425 94.170 193.265 ;
        RECT 95.045 193.060 95.235 193.265 ;
        RECT 95.965 193.145 96.135 193.725 ;
        RECT 96.765 193.755 97.975 194.505 ;
        RECT 98.145 193.945 98.405 194.225 ;
        RECT 98.575 194.115 99.835 194.285 ;
        RECT 100.005 193.945 100.280 194.310 ;
        RECT 100.515 194.065 100.685 194.505 ;
        RECT 98.145 193.765 98.900 193.945 ;
        RECT 99.070 193.895 100.280 193.945 ;
        RECT 100.855 193.895 101.195 194.310 ;
        RECT 99.070 193.765 101.195 193.895 ;
        RECT 96.765 193.215 97.285 193.755 ;
        RECT 95.920 193.095 96.135 193.145 ;
        RECT 94.340 192.685 95.235 193.060 ;
        RECT 95.745 193.015 96.135 193.095 ;
        RECT 97.455 193.045 97.975 193.585 ;
        RECT 98.145 193.265 98.525 193.595 ;
        RECT 98.695 193.095 98.900 193.765 ;
        RECT 100.165 193.725 101.195 193.765 ;
        RECT 102.285 193.765 102.625 194.335 ;
        RECT 102.820 193.840 102.990 194.505 ;
        RECT 103.270 194.165 103.490 194.210 ;
        RECT 103.265 193.995 103.490 194.165 ;
        RECT 103.660 194.025 104.105 194.195 ;
        RECT 103.270 193.855 103.490 193.995 ;
        RECT 99.070 193.265 99.415 193.595 ;
        RECT 99.585 193.265 100.045 193.595 ;
        RECT 100.225 193.345 100.565 193.515 ;
        RECT 100.355 193.145 100.565 193.345 ;
        RECT 100.735 193.315 101.195 193.515 ;
        RECT 93.285 192.255 94.170 192.425 ;
        RECT 94.350 191.955 94.665 192.455 ;
        RECT 94.895 192.125 95.235 192.685 ;
        RECT 95.405 191.955 95.575 192.965 ;
        RECT 95.745 192.170 96.075 193.015 ;
        RECT 96.245 191.955 96.415 192.870 ;
        RECT 96.765 191.955 97.975 193.045 ;
        RECT 98.145 192.885 100.185 193.095 ;
        RECT 100.355 192.975 100.735 193.145 ;
        RECT 98.145 192.125 98.425 192.885 ;
        RECT 99.795 192.805 100.185 192.885 ;
        RECT 98.610 191.955 99.400 192.715 ;
        RECT 99.795 192.125 100.305 192.805 ;
        RECT 100.525 192.465 100.735 192.975 ;
        RECT 100.505 192.295 100.735 192.465 ;
        RECT 100.525 192.185 100.735 192.295 ;
        RECT 100.935 191.955 101.195 193.135 ;
        RECT 102.285 192.795 102.460 193.765 ;
        RECT 103.270 193.685 103.765 193.855 ;
        RECT 102.630 193.145 102.800 193.595 ;
        RECT 102.970 193.315 103.420 193.515 ;
        RECT 103.590 193.490 103.765 193.685 ;
        RECT 103.935 193.235 104.105 194.025 ;
        RECT 104.275 193.900 104.525 194.270 ;
        RECT 104.355 193.515 104.525 193.900 ;
        RECT 104.695 193.865 104.945 194.270 ;
        RECT 105.115 194.035 105.285 194.505 ;
        RECT 105.455 193.865 105.795 194.270 ;
        RECT 104.695 193.685 105.795 193.865 ;
        RECT 105.965 193.735 107.635 194.505 ;
        RECT 108.270 193.765 108.525 194.335 ;
        RECT 108.695 194.105 109.025 194.505 ;
        RECT 109.450 193.970 109.980 194.335 ;
        RECT 109.450 193.935 109.625 193.970 ;
        RECT 108.695 193.765 109.625 193.935 ;
        RECT 104.355 193.345 104.550 193.515 ;
        RECT 102.630 192.975 103.025 193.145 ;
        RECT 103.935 193.095 104.210 193.235 ;
        RECT 102.285 192.125 102.545 192.795 ;
        RECT 102.855 192.705 103.025 192.975 ;
        RECT 103.195 192.875 104.210 193.095 ;
        RECT 104.380 193.095 104.550 193.345 ;
        RECT 104.720 193.265 105.280 193.515 ;
        RECT 104.380 192.705 104.935 193.095 ;
        RECT 102.855 192.535 104.935 192.705 ;
        RECT 102.715 191.955 103.045 192.355 ;
        RECT 103.915 191.955 104.315 192.355 ;
        RECT 104.605 192.300 104.935 192.535 ;
        RECT 105.105 192.165 105.280 193.265 ;
        RECT 105.450 192.945 105.795 193.515 ;
        RECT 105.965 193.215 106.715 193.735 ;
        RECT 106.885 193.045 107.635 193.565 ;
        RECT 105.450 191.955 105.795 192.775 ;
        RECT 105.965 191.955 107.635 193.045 ;
        RECT 108.270 193.095 108.440 193.765 ;
        RECT 108.695 193.595 108.865 193.765 ;
        RECT 108.610 193.265 108.865 193.595 ;
        RECT 109.090 193.265 109.285 193.595 ;
        RECT 108.270 192.125 108.605 193.095 ;
        RECT 108.775 191.955 108.945 193.095 ;
        RECT 109.115 192.295 109.285 193.265 ;
        RECT 109.455 192.635 109.625 193.765 ;
        RECT 109.795 192.975 109.965 193.775 ;
        RECT 110.170 193.485 110.445 194.335 ;
        RECT 110.165 193.315 110.445 193.485 ;
        RECT 110.170 193.175 110.445 193.315 ;
        RECT 110.615 192.975 110.805 194.335 ;
        RECT 110.985 193.970 111.495 194.505 ;
        RECT 111.715 193.695 111.960 194.300 ;
        RECT 112.405 193.735 114.075 194.505 ;
        RECT 114.245 193.780 114.535 194.505 ;
        RECT 114.705 193.735 118.215 194.505 ;
        RECT 118.405 193.775 118.695 194.505 ;
        RECT 111.005 193.525 112.235 193.695 ;
        RECT 109.795 192.805 110.805 192.975 ;
        RECT 110.975 192.960 111.725 193.150 ;
        RECT 109.455 192.465 110.580 192.635 ;
        RECT 110.975 192.295 111.145 192.960 ;
        RECT 111.895 192.715 112.235 193.525 ;
        RECT 112.405 193.215 113.155 193.735 ;
        RECT 113.325 193.045 114.075 193.565 ;
        RECT 114.705 193.215 116.355 193.735 ;
        RECT 109.115 192.125 111.145 192.295 ;
        RECT 111.315 191.955 111.485 192.715 ;
        RECT 111.720 192.305 112.235 192.715 ;
        RECT 112.405 191.955 114.075 193.045 ;
        RECT 114.245 191.955 114.535 193.120 ;
        RECT 116.525 193.045 118.215 193.565 ;
        RECT 118.395 193.265 118.695 193.595 ;
        RECT 118.875 193.575 119.105 194.215 ;
        RECT 119.285 193.955 119.595 194.325 ;
        RECT 119.775 194.135 120.445 194.505 ;
        RECT 119.285 193.755 120.515 193.955 ;
        RECT 118.875 193.265 119.400 193.575 ;
        RECT 119.580 193.265 120.045 193.575 ;
        RECT 120.225 193.085 120.515 193.755 ;
        RECT 114.705 191.955 118.215 193.045 ;
        RECT 118.405 192.845 119.565 193.085 ;
        RECT 118.405 192.135 118.665 192.845 ;
        RECT 118.835 191.955 119.165 192.665 ;
        RECT 119.335 192.135 119.565 192.845 ;
        RECT 119.745 192.865 120.515 193.085 ;
        RECT 119.745 192.135 120.015 192.865 ;
        RECT 120.195 191.955 120.535 192.685 ;
        RECT 120.705 192.135 120.965 194.325 ;
        RECT 121.165 193.935 121.420 194.285 ;
        RECT 121.590 194.105 121.920 194.505 ;
        RECT 122.090 193.935 122.260 194.285 ;
        RECT 122.430 194.105 122.810 194.505 ;
        RECT 121.165 193.765 122.830 193.935 ;
        RECT 123.000 193.830 123.275 194.175 ;
        RECT 122.660 193.595 122.830 193.765 ;
        RECT 121.145 193.265 121.495 193.595 ;
        RECT 121.665 193.265 122.490 193.595 ;
        RECT 122.660 193.265 122.935 193.595 ;
        RECT 121.165 192.805 121.495 193.095 ;
        RECT 121.665 192.975 121.890 193.265 ;
        RECT 122.660 193.095 122.830 193.265 ;
        RECT 123.105 193.095 123.275 193.830 ;
        RECT 123.445 193.675 123.735 194.505 ;
        RECT 123.905 193.705 124.600 194.335 ;
        RECT 124.805 193.705 125.115 194.505 ;
        RECT 125.485 193.875 125.815 194.235 ;
        RECT 126.435 194.045 126.685 194.505 ;
        RECT 126.855 194.045 127.415 194.335 ;
        RECT 123.925 193.265 124.260 193.515 ;
        RECT 122.160 192.925 122.830 193.095 ;
        RECT 122.160 192.805 122.330 192.925 ;
        RECT 121.165 192.635 122.330 192.805 ;
        RECT 121.145 192.175 122.340 192.465 ;
        RECT 122.510 191.955 122.790 192.755 ;
        RECT 123.000 192.125 123.275 193.095 ;
        RECT 123.445 191.955 123.735 193.160 ;
        RECT 124.430 193.105 124.600 193.705 ;
        RECT 125.485 193.685 126.875 193.875 ;
        RECT 126.705 193.595 126.875 193.685 ;
        RECT 124.770 193.265 125.105 193.535 ;
        RECT 125.300 193.265 125.975 193.515 ;
        RECT 126.195 193.265 126.535 193.515 ;
        RECT 126.705 193.265 126.995 193.595 ;
        RECT 123.905 191.955 124.165 193.095 ;
        RECT 124.335 192.125 124.665 193.105 ;
        RECT 124.835 191.955 125.115 193.095 ;
        RECT 125.300 192.905 125.565 193.265 ;
        RECT 126.705 193.015 126.875 193.265 ;
        RECT 125.935 192.845 126.875 193.015 ;
        RECT 125.485 191.955 125.765 192.625 ;
        RECT 125.935 192.295 126.235 192.845 ;
        RECT 127.165 192.675 127.415 194.045 ;
        RECT 127.675 193.955 127.845 194.245 ;
        RECT 128.015 194.125 128.345 194.505 ;
        RECT 127.675 193.785 128.340 193.955 ;
        RECT 127.590 192.965 127.940 193.615 ;
        RECT 128.110 192.795 128.340 193.785 ;
        RECT 126.435 191.955 126.765 192.675 ;
        RECT 126.955 192.125 127.415 192.675 ;
        RECT 127.675 192.625 128.340 192.795 ;
        RECT 127.675 192.125 127.845 192.625 ;
        RECT 128.015 191.955 128.345 192.455 ;
        RECT 128.515 192.125 128.700 194.245 ;
        RECT 128.955 194.045 129.205 194.505 ;
        RECT 129.375 194.055 129.710 194.225 ;
        RECT 129.905 194.055 130.580 194.225 ;
        RECT 129.375 193.915 129.545 194.055 ;
        RECT 128.870 192.925 129.150 193.875 ;
        RECT 129.320 193.785 129.545 193.915 ;
        RECT 129.320 192.680 129.490 193.785 ;
        RECT 129.715 193.635 130.240 193.855 ;
        RECT 129.660 192.870 129.900 193.465 ;
        RECT 130.070 192.935 130.240 193.635 ;
        RECT 130.410 193.275 130.580 194.055 ;
        RECT 130.900 194.005 131.270 194.505 ;
        RECT 131.450 194.055 131.855 194.225 ;
        RECT 132.025 194.055 132.810 194.225 ;
        RECT 131.450 193.825 131.620 194.055 ;
        RECT 130.790 193.525 131.620 193.825 ;
        RECT 132.005 193.555 132.470 193.885 ;
        RECT 130.790 193.495 130.990 193.525 ;
        RECT 131.110 193.275 131.280 193.345 ;
        RECT 130.410 193.105 131.280 193.275 ;
        RECT 130.770 193.015 131.280 193.105 ;
        RECT 129.320 192.550 129.625 192.680 ;
        RECT 130.070 192.570 130.600 192.935 ;
        RECT 128.940 191.955 129.205 192.415 ;
        RECT 129.375 192.125 129.625 192.550 ;
        RECT 130.770 192.400 130.940 193.015 ;
        RECT 129.835 192.230 130.940 192.400 ;
        RECT 131.110 191.955 131.280 192.755 ;
        RECT 131.450 192.455 131.620 193.525 ;
        RECT 131.790 192.625 131.980 193.345 ;
        RECT 132.150 192.595 132.470 193.555 ;
        RECT 132.640 193.595 132.810 194.055 ;
        RECT 133.085 193.975 133.295 194.505 ;
        RECT 133.555 193.765 133.885 194.290 ;
        RECT 134.055 193.895 134.225 194.505 ;
        RECT 134.395 193.850 134.725 194.285 ;
        RECT 134.895 193.990 135.065 194.505 ;
        RECT 134.395 193.765 134.775 193.850 ;
        RECT 133.685 193.595 133.885 193.765 ;
        RECT 134.550 193.725 134.775 193.765 ;
        RECT 132.640 193.265 133.515 193.595 ;
        RECT 133.685 193.265 134.435 193.595 ;
        RECT 131.450 192.125 131.700 192.455 ;
        RECT 132.640 192.425 132.810 193.265 ;
        RECT 133.685 193.060 133.875 193.265 ;
        RECT 134.605 193.145 134.775 193.725 ;
        RECT 135.405 193.735 138.915 194.505 ;
        RECT 140.005 193.780 140.295 194.505 ;
        RECT 140.465 193.960 145.810 194.505 ;
        RECT 135.405 193.215 137.055 193.735 ;
        RECT 134.560 193.095 134.775 193.145 ;
        RECT 132.980 192.685 133.875 193.060 ;
        RECT 134.385 193.015 134.775 193.095 ;
        RECT 137.225 193.045 138.915 193.565 ;
        RECT 142.050 193.130 142.390 193.960 ;
        RECT 145.985 193.735 148.575 194.505 ;
        RECT 149.205 193.755 150.415 194.505 ;
        RECT 131.925 192.255 132.810 192.425 ;
        RECT 132.990 191.955 133.305 192.455 ;
        RECT 133.535 192.125 133.875 192.685 ;
        RECT 134.045 191.955 134.215 192.965 ;
        RECT 134.385 192.170 134.715 193.015 ;
        RECT 134.885 191.955 135.055 192.870 ;
        RECT 135.405 191.955 138.915 193.045 ;
        RECT 140.005 191.955 140.295 193.120 ;
        RECT 143.870 192.390 144.220 193.640 ;
        RECT 145.985 193.215 147.195 193.735 ;
        RECT 147.365 193.045 148.575 193.565 ;
        RECT 140.465 191.955 145.810 192.390 ;
        RECT 145.985 191.955 148.575 193.045 ;
        RECT 149.205 193.045 149.725 193.585 ;
        RECT 149.895 193.215 150.415 193.755 ;
        RECT 149.205 191.955 150.415 193.045 ;
        RECT 11.120 191.785 150.500 191.955 ;
        RECT 11.205 190.695 12.415 191.785 ;
        RECT 12.675 191.115 12.845 191.615 ;
        RECT 13.015 191.285 13.345 191.785 ;
        RECT 12.675 190.945 13.340 191.115 ;
        RECT 11.205 189.985 11.725 190.525 ;
        RECT 11.895 190.155 12.415 190.695 ;
        RECT 12.590 190.125 12.940 190.775 ;
        RECT 11.205 189.235 12.415 189.985 ;
        RECT 13.110 189.955 13.340 190.945 ;
        RECT 12.675 189.785 13.340 189.955 ;
        RECT 12.675 189.495 12.845 189.785 ;
        RECT 13.015 189.235 13.345 189.615 ;
        RECT 13.515 189.495 13.700 191.615 ;
        RECT 13.940 191.325 14.205 191.785 ;
        RECT 14.375 191.190 14.625 191.615 ;
        RECT 14.835 191.340 15.940 191.510 ;
        RECT 14.320 191.060 14.625 191.190 ;
        RECT 13.870 189.865 14.150 190.815 ;
        RECT 14.320 189.955 14.490 191.060 ;
        RECT 14.660 190.275 14.900 190.870 ;
        RECT 15.070 190.805 15.600 191.170 ;
        RECT 15.070 190.105 15.240 190.805 ;
        RECT 15.770 190.725 15.940 191.340 ;
        RECT 16.110 190.985 16.280 191.785 ;
        RECT 16.450 191.285 16.700 191.615 ;
        RECT 16.925 191.315 17.810 191.485 ;
        RECT 15.770 190.635 16.280 190.725 ;
        RECT 14.320 189.825 14.545 189.955 ;
        RECT 14.715 189.885 15.240 190.105 ;
        RECT 15.410 190.465 16.280 190.635 ;
        RECT 13.955 189.235 14.205 189.695 ;
        RECT 14.375 189.685 14.545 189.825 ;
        RECT 15.410 189.685 15.580 190.465 ;
        RECT 16.110 190.395 16.280 190.465 ;
        RECT 15.790 190.215 15.990 190.245 ;
        RECT 16.450 190.215 16.620 191.285 ;
        RECT 16.790 190.395 16.980 191.115 ;
        RECT 15.790 189.915 16.620 190.215 ;
        RECT 17.150 190.185 17.470 191.145 ;
        RECT 14.375 189.515 14.710 189.685 ;
        RECT 14.905 189.515 15.580 189.685 ;
        RECT 15.900 189.235 16.270 189.735 ;
        RECT 16.450 189.685 16.620 189.915 ;
        RECT 17.005 189.855 17.470 190.185 ;
        RECT 17.640 190.475 17.810 191.315 ;
        RECT 17.990 191.285 18.305 191.785 ;
        RECT 18.535 191.055 18.875 191.615 ;
        RECT 17.980 190.680 18.875 191.055 ;
        RECT 19.045 190.775 19.215 191.785 ;
        RECT 18.685 190.475 18.875 190.680 ;
        RECT 19.385 190.725 19.715 191.570 ;
        RECT 19.385 190.645 19.775 190.725 ;
        RECT 19.560 190.595 19.775 190.645 ;
        RECT 19.950 190.635 20.210 191.785 ;
        RECT 20.385 190.710 20.640 191.615 ;
        RECT 20.810 191.025 21.140 191.785 ;
        RECT 21.355 190.855 21.525 191.615 ;
        RECT 17.640 190.145 18.515 190.475 ;
        RECT 18.685 190.145 19.435 190.475 ;
        RECT 17.640 189.685 17.810 190.145 ;
        RECT 18.685 189.975 18.885 190.145 ;
        RECT 19.605 190.015 19.775 190.595 ;
        RECT 19.550 189.975 19.775 190.015 ;
        RECT 16.450 189.515 16.855 189.685 ;
        RECT 17.025 189.515 17.810 189.685 ;
        RECT 18.085 189.235 18.295 189.765 ;
        RECT 18.555 189.450 18.885 189.975 ;
        RECT 19.395 189.890 19.775 189.975 ;
        RECT 19.055 189.235 19.225 189.845 ;
        RECT 19.395 189.455 19.725 189.890 ;
        RECT 19.950 189.235 20.210 190.075 ;
        RECT 20.385 189.980 20.555 190.710 ;
        RECT 20.810 190.685 21.525 190.855 ;
        RECT 21.785 190.710 22.055 191.615 ;
        RECT 22.225 191.025 22.555 191.785 ;
        RECT 22.735 190.855 22.905 191.615 ;
        RECT 20.810 190.475 20.980 190.685 ;
        RECT 20.725 190.145 20.980 190.475 ;
        RECT 20.385 189.405 20.640 189.980 ;
        RECT 20.810 189.955 20.980 190.145 ;
        RECT 21.260 190.135 21.615 190.505 ;
        RECT 20.810 189.785 21.525 189.955 ;
        RECT 20.810 189.235 21.140 189.615 ;
        RECT 21.355 189.405 21.525 189.785 ;
        RECT 21.785 189.910 21.955 190.710 ;
        RECT 22.240 190.685 22.905 190.855 ;
        RECT 22.240 190.540 22.410 190.685 ;
        RECT 24.085 190.620 24.375 191.785 ;
        RECT 24.545 190.695 27.135 191.785 ;
        RECT 22.125 190.210 22.410 190.540 ;
        RECT 22.240 189.955 22.410 190.210 ;
        RECT 22.645 190.135 22.975 190.505 ;
        RECT 24.545 190.005 25.755 190.525 ;
        RECT 25.925 190.175 27.135 190.695 ;
        RECT 27.310 190.635 27.570 191.785 ;
        RECT 27.745 190.710 28.000 191.615 ;
        RECT 28.170 191.025 28.500 191.785 ;
        RECT 28.715 190.855 28.885 191.615 ;
        RECT 21.785 189.405 22.045 189.910 ;
        RECT 22.240 189.785 22.905 189.955 ;
        RECT 22.225 189.235 22.555 189.615 ;
        RECT 22.735 189.405 22.905 189.785 ;
        RECT 24.085 189.235 24.375 189.960 ;
        RECT 24.545 189.235 27.135 190.005 ;
        RECT 27.310 189.235 27.570 190.075 ;
        RECT 27.745 189.980 27.915 190.710 ;
        RECT 28.170 190.685 28.885 190.855 ;
        RECT 28.170 190.475 28.340 190.685 ;
        RECT 29.150 190.645 29.405 191.785 ;
        RECT 29.600 191.235 30.795 191.565 ;
        RECT 28.085 190.145 28.340 190.475 ;
        RECT 27.745 189.405 28.000 189.980 ;
        RECT 28.170 189.955 28.340 190.145 ;
        RECT 28.620 190.135 28.975 190.505 ;
        RECT 29.655 190.475 29.825 191.035 ;
        RECT 30.050 190.815 30.470 191.065 ;
        RECT 30.975 190.985 31.255 191.785 ;
        RECT 30.050 190.645 31.295 190.815 ;
        RECT 31.465 190.645 31.735 191.615 ;
        RECT 31.125 190.475 31.295 190.645 ;
        RECT 29.150 190.225 29.485 190.475 ;
        RECT 29.655 190.145 30.395 190.475 ;
        RECT 31.125 190.145 31.355 190.475 ;
        RECT 29.655 190.055 29.905 190.145 ;
        RECT 28.170 189.785 28.885 189.955 ;
        RECT 28.170 189.235 28.500 189.615 ;
        RECT 28.715 189.405 28.885 189.785 ;
        RECT 29.170 189.885 29.905 190.055 ;
        RECT 31.125 189.975 31.295 190.145 ;
        RECT 29.170 189.415 29.480 189.885 ;
        RECT 30.555 189.805 31.295 189.975 ;
        RECT 31.565 189.910 31.735 190.645 ;
        RECT 29.650 189.235 30.385 189.715 ;
        RECT 30.555 189.455 30.725 189.805 ;
        RECT 30.895 189.235 31.275 189.635 ;
        RECT 31.465 189.565 31.735 189.910 ;
        RECT 32.365 190.915 32.640 191.615 ;
        RECT 32.850 191.240 33.065 191.785 ;
        RECT 33.235 191.275 33.710 191.615 ;
        RECT 33.880 191.280 34.495 191.785 ;
        RECT 33.880 191.105 34.075 191.280 ;
        RECT 32.365 189.885 32.535 190.915 ;
        RECT 32.810 190.745 33.525 191.040 ;
        RECT 33.745 190.915 34.075 191.105 ;
        RECT 34.245 190.745 34.495 191.110 ;
        RECT 32.705 190.575 34.495 190.745 ;
        RECT 32.705 190.145 32.935 190.575 ;
        RECT 32.365 189.405 32.625 189.885 ;
        RECT 33.105 189.875 33.515 190.395 ;
        RECT 32.795 189.235 33.125 189.695 ;
        RECT 33.315 189.455 33.515 189.875 ;
        RECT 33.685 189.720 33.940 190.575 ;
        RECT 34.735 190.395 34.905 191.615 ;
        RECT 35.155 191.275 35.415 191.785 ;
        RECT 34.110 190.145 34.905 190.395 ;
        RECT 35.075 190.225 35.415 191.105 ;
        RECT 35.585 190.695 39.095 191.785 ;
        RECT 34.655 190.055 34.905 190.145 ;
        RECT 33.685 189.455 34.475 189.720 ;
        RECT 34.655 189.635 34.985 190.055 ;
        RECT 35.155 189.235 35.415 190.055 ;
        RECT 35.585 190.005 37.235 190.525 ;
        RECT 37.405 190.175 39.095 190.695 ;
        RECT 39.275 191.175 39.605 191.605 ;
        RECT 39.785 191.345 39.980 191.785 ;
        RECT 40.150 191.175 40.480 191.605 ;
        RECT 39.275 191.005 40.480 191.175 ;
        RECT 39.275 190.675 40.170 191.005 ;
        RECT 40.650 190.835 40.925 191.605 ;
        RECT 41.105 191.350 46.450 191.785 ;
        RECT 40.340 190.645 40.925 190.835 ;
        RECT 39.280 190.145 39.575 190.475 ;
        RECT 39.755 190.145 40.170 190.475 ;
        RECT 35.585 189.235 39.095 190.005 ;
        RECT 39.275 189.235 39.575 189.965 ;
        RECT 39.755 189.525 39.985 190.145 ;
        RECT 40.340 189.975 40.515 190.645 ;
        RECT 40.185 189.795 40.515 189.975 ;
        RECT 40.685 189.825 40.925 190.475 ;
        RECT 40.185 189.415 40.410 189.795 ;
        RECT 42.690 189.780 43.030 190.610 ;
        RECT 44.510 190.100 44.860 191.350 ;
        RECT 46.625 190.695 49.215 191.785 ;
        RECT 46.625 190.005 47.835 190.525 ;
        RECT 48.005 190.175 49.215 190.695 ;
        RECT 49.845 190.620 50.135 191.785 ;
        RECT 50.305 190.695 52.895 191.785 ;
        RECT 50.305 190.005 51.515 190.525 ;
        RECT 51.685 190.175 52.895 190.695 ;
        RECT 53.100 190.995 53.635 191.615 ;
        RECT 40.580 189.235 40.910 189.625 ;
        RECT 41.105 189.235 46.450 189.780 ;
        RECT 46.625 189.235 49.215 190.005 ;
        RECT 49.845 189.235 50.135 189.960 ;
        RECT 50.305 189.235 52.895 190.005 ;
        RECT 53.100 189.975 53.415 190.995 ;
        RECT 53.805 190.985 54.135 191.785 ;
        RECT 54.620 190.815 55.010 190.990 ;
        RECT 53.585 190.645 55.010 190.815 ;
        RECT 55.455 190.855 55.625 191.615 ;
        RECT 55.805 191.025 56.135 191.785 ;
        RECT 55.455 190.685 56.120 190.855 ;
        RECT 56.305 190.710 56.575 191.615 ;
        RECT 56.745 191.350 62.090 191.785 ;
        RECT 62.265 191.350 67.610 191.785 ;
        RECT 53.585 190.145 53.755 190.645 ;
        RECT 53.100 189.405 53.715 189.975 ;
        RECT 54.005 189.915 54.270 190.475 ;
        RECT 54.440 189.745 54.610 190.645 ;
        RECT 55.950 190.540 56.120 190.685 ;
        RECT 54.780 189.915 55.135 190.475 ;
        RECT 55.385 190.135 55.715 190.505 ;
        RECT 55.950 190.210 56.235 190.540 ;
        RECT 55.950 189.955 56.120 190.210 ;
        RECT 55.455 189.785 56.120 189.955 ;
        RECT 56.405 189.910 56.575 190.710 ;
        RECT 53.885 189.235 54.100 189.745 ;
        RECT 54.330 189.415 54.610 189.745 ;
        RECT 54.790 189.235 55.030 189.745 ;
        RECT 55.455 189.405 55.625 189.785 ;
        RECT 55.805 189.235 56.135 189.615 ;
        RECT 56.315 189.405 56.575 189.910 ;
        RECT 58.330 189.780 58.670 190.610 ;
        RECT 60.150 190.100 60.500 191.350 ;
        RECT 63.850 189.780 64.190 190.610 ;
        RECT 65.670 190.100 66.020 191.350 ;
        RECT 67.785 190.695 69.455 191.785 ;
        RECT 67.785 190.005 68.535 190.525 ;
        RECT 68.705 190.175 69.455 190.695 ;
        RECT 70.085 190.645 70.365 191.785 ;
        RECT 70.535 190.635 70.865 191.615 ;
        RECT 71.035 190.645 71.295 191.785 ;
        RECT 71.465 190.695 74.975 191.785 ;
        RECT 70.095 190.205 70.430 190.475 ;
        RECT 70.600 190.035 70.770 190.635 ;
        RECT 70.940 190.225 71.275 190.475 ;
        RECT 56.745 189.235 62.090 189.780 ;
        RECT 62.265 189.235 67.610 189.780 ;
        RECT 67.785 189.235 69.455 190.005 ;
        RECT 70.085 189.235 70.395 190.035 ;
        RECT 70.600 189.405 71.295 190.035 ;
        RECT 71.465 190.005 73.115 190.525 ;
        RECT 73.285 190.175 74.975 190.695 ;
        RECT 75.605 190.620 75.895 191.785 ;
        RECT 76.065 190.695 77.735 191.785 ;
        RECT 76.065 190.005 76.815 190.525 ;
        RECT 76.985 190.175 77.735 190.695 ;
        RECT 78.445 190.855 78.625 191.615 ;
        RECT 78.805 191.025 79.135 191.785 ;
        RECT 78.445 190.685 79.120 190.855 ;
        RECT 79.305 190.710 79.575 191.615 ;
        RECT 79.745 191.350 85.090 191.785 ;
        RECT 78.950 190.540 79.120 190.685 ;
        RECT 78.385 190.135 78.725 190.505 ;
        RECT 78.950 190.210 79.225 190.540 ;
        RECT 71.465 189.235 74.975 190.005 ;
        RECT 75.605 189.235 75.895 189.960 ;
        RECT 76.065 189.235 77.735 190.005 ;
        RECT 78.950 189.955 79.120 190.210 ;
        RECT 78.455 189.785 79.120 189.955 ;
        RECT 79.395 189.910 79.575 190.710 ;
        RECT 78.455 189.405 78.625 189.785 ;
        RECT 78.805 189.235 79.135 189.615 ;
        RECT 79.315 189.405 79.575 189.910 ;
        RECT 81.330 189.780 81.670 190.610 ;
        RECT 83.150 190.100 83.500 191.350 ;
        RECT 85.265 190.695 86.475 191.785 ;
        RECT 86.735 191.040 87.005 191.785 ;
        RECT 87.635 191.780 93.910 191.785 ;
        RECT 87.175 190.870 87.465 191.610 ;
        RECT 87.635 191.055 87.890 191.780 ;
        RECT 88.075 190.885 88.335 191.610 ;
        RECT 88.505 191.055 88.750 191.780 ;
        RECT 88.935 190.885 89.195 191.610 ;
        RECT 89.365 191.055 89.610 191.780 ;
        RECT 89.795 190.885 90.055 191.610 ;
        RECT 90.225 191.055 90.470 191.780 ;
        RECT 90.640 190.885 90.900 191.610 ;
        RECT 91.070 191.055 91.330 191.780 ;
        RECT 91.500 190.885 91.760 191.610 ;
        RECT 91.930 191.055 92.190 191.780 ;
        RECT 92.360 190.885 92.620 191.610 ;
        RECT 92.790 191.055 93.050 191.780 ;
        RECT 93.220 190.885 93.480 191.610 ;
        RECT 93.650 190.985 93.910 191.780 ;
        RECT 88.075 190.870 93.480 190.885 ;
        RECT 85.265 189.985 85.785 190.525 ;
        RECT 85.955 190.155 86.475 190.695 ;
        RECT 86.735 190.645 93.480 190.870 ;
        RECT 86.735 190.055 87.900 190.645 ;
        RECT 94.080 190.475 94.330 191.610 ;
        RECT 94.510 190.975 94.770 191.785 ;
        RECT 94.945 190.475 95.190 191.615 ;
        RECT 95.370 190.975 95.665 191.785 ;
        RECT 95.935 190.775 96.105 191.615 ;
        RECT 96.275 191.445 97.445 191.615 ;
        RECT 96.275 190.945 96.605 191.445 ;
        RECT 97.115 191.405 97.445 191.445 ;
        RECT 97.635 191.365 97.990 191.785 ;
        RECT 96.775 191.185 97.005 191.275 ;
        RECT 98.160 191.185 98.410 191.615 ;
        RECT 96.775 190.945 98.410 191.185 ;
        RECT 98.580 191.025 98.910 191.785 ;
        RECT 99.080 190.945 99.335 191.615 ;
        RECT 95.935 190.605 98.995 190.775 ;
        RECT 88.070 190.225 95.190 190.475 ;
        RECT 79.745 189.235 85.090 189.780 ;
        RECT 85.265 189.235 86.475 189.985 ;
        RECT 86.735 189.885 93.480 190.055 ;
        RECT 86.735 189.235 87.035 189.715 ;
        RECT 87.205 189.430 87.465 189.885 ;
        RECT 87.635 189.235 87.895 189.715 ;
        RECT 88.075 189.430 88.335 189.885 ;
        RECT 88.505 189.235 88.755 189.715 ;
        RECT 88.935 189.430 89.195 189.885 ;
        RECT 89.365 189.235 89.615 189.715 ;
        RECT 89.795 189.430 90.055 189.885 ;
        RECT 90.225 189.235 90.470 189.715 ;
        RECT 90.640 189.430 90.915 189.885 ;
        RECT 91.085 189.235 91.330 189.715 ;
        RECT 91.500 189.430 91.760 189.885 ;
        RECT 91.930 189.235 92.190 189.715 ;
        RECT 92.360 189.430 92.620 189.885 ;
        RECT 92.790 189.235 93.050 189.715 ;
        RECT 93.220 189.430 93.480 189.885 ;
        RECT 93.650 189.235 93.910 189.795 ;
        RECT 94.080 189.415 94.330 190.225 ;
        RECT 94.510 189.235 94.770 189.760 ;
        RECT 94.940 189.415 95.190 190.225 ;
        RECT 95.360 189.915 95.675 190.475 ;
        RECT 95.850 190.225 96.200 190.435 ;
        RECT 96.370 190.225 96.815 190.425 ;
        RECT 96.985 190.225 97.460 190.425 ;
        RECT 95.935 189.885 97.000 190.055 ;
        RECT 95.370 189.235 95.675 189.745 ;
        RECT 95.935 189.405 96.105 189.885 ;
        RECT 96.275 189.235 96.605 189.715 ;
        RECT 96.830 189.655 97.000 189.885 ;
        RECT 97.180 189.825 97.460 190.225 ;
        RECT 97.730 190.225 98.060 190.425 ;
        RECT 98.230 190.255 98.605 190.425 ;
        RECT 98.230 190.225 98.595 190.255 ;
        RECT 97.730 189.825 98.015 190.225 ;
        RECT 98.825 190.055 98.995 190.605 ;
        RECT 98.195 189.885 98.995 190.055 ;
        RECT 98.195 189.655 98.365 189.885 ;
        RECT 99.165 189.815 99.335 190.945 ;
        RECT 99.525 190.695 101.195 191.785 ;
        RECT 99.150 189.745 99.335 189.815 ;
        RECT 99.125 189.735 99.335 189.745 ;
        RECT 96.830 189.405 98.365 189.655 ;
        RECT 98.535 189.235 98.865 189.715 ;
        RECT 99.080 189.405 99.335 189.735 ;
        RECT 99.525 190.005 100.275 190.525 ;
        RECT 100.445 190.175 101.195 190.695 ;
        RECT 101.365 190.620 101.655 191.785 ;
        RECT 101.835 190.975 102.130 191.785 ;
        RECT 102.310 190.475 102.555 191.615 ;
        RECT 102.730 190.975 102.990 191.785 ;
        RECT 103.590 191.780 109.865 191.785 ;
        RECT 103.170 190.475 103.420 191.610 ;
        RECT 103.590 190.985 103.850 191.780 ;
        RECT 104.020 190.885 104.280 191.610 ;
        RECT 104.450 191.055 104.710 191.780 ;
        RECT 104.880 190.885 105.140 191.610 ;
        RECT 105.310 191.055 105.570 191.780 ;
        RECT 105.740 190.885 106.000 191.610 ;
        RECT 106.170 191.055 106.430 191.780 ;
        RECT 106.600 190.885 106.860 191.610 ;
        RECT 107.030 191.055 107.275 191.780 ;
        RECT 107.445 190.885 107.705 191.610 ;
        RECT 107.890 191.055 108.135 191.780 ;
        RECT 108.305 190.885 108.565 191.610 ;
        RECT 108.750 191.055 108.995 191.780 ;
        RECT 109.165 190.885 109.425 191.610 ;
        RECT 109.610 191.055 109.865 191.780 ;
        RECT 104.020 190.870 109.425 190.885 ;
        RECT 110.035 190.870 110.325 191.610 ;
        RECT 110.495 191.040 110.765 191.785 ;
        RECT 104.020 190.645 110.765 190.870 ;
        RECT 99.525 189.235 101.195 190.005 ;
        RECT 101.365 189.235 101.655 189.960 ;
        RECT 101.825 189.915 102.140 190.475 ;
        RECT 102.310 190.225 109.430 190.475 ;
        RECT 101.825 189.235 102.130 189.745 ;
        RECT 102.310 189.415 102.560 190.225 ;
        RECT 102.730 189.235 102.990 189.760 ;
        RECT 103.170 189.415 103.420 190.225 ;
        RECT 109.600 190.055 110.765 190.645 ;
        RECT 111.025 190.685 111.345 191.615 ;
        RECT 111.525 191.105 111.925 191.615 ;
        RECT 112.095 191.275 112.265 191.785 ;
        RECT 112.435 191.105 112.765 191.615 ;
        RECT 111.525 190.935 112.765 191.105 ;
        RECT 112.935 190.935 113.105 191.785 ;
        RECT 113.695 190.935 114.075 191.615 ;
        RECT 111.025 190.515 111.655 190.685 ;
        RECT 104.020 189.885 110.765 190.055 ;
        RECT 103.590 189.235 103.850 189.795 ;
        RECT 104.020 189.430 104.280 189.885 ;
        RECT 104.450 189.235 104.710 189.715 ;
        RECT 104.880 189.430 105.140 189.885 ;
        RECT 105.310 189.235 105.570 189.715 ;
        RECT 105.740 189.430 106.000 189.885 ;
        RECT 106.170 189.235 106.415 189.715 ;
        RECT 106.585 189.430 106.860 189.885 ;
        RECT 107.030 189.235 107.275 189.715 ;
        RECT 107.445 189.430 107.705 189.885 ;
        RECT 107.885 189.235 108.135 189.715 ;
        RECT 108.305 189.430 108.565 189.885 ;
        RECT 108.745 189.235 108.995 189.715 ;
        RECT 109.165 189.430 109.425 189.885 ;
        RECT 109.605 189.235 109.865 189.715 ;
        RECT 110.035 189.430 110.295 189.885 ;
        RECT 110.465 189.235 110.765 189.715 ;
        RECT 111.025 189.235 111.315 190.070 ;
        RECT 111.485 189.635 111.655 190.515 ;
        RECT 112.430 190.595 113.735 190.765 ;
        RECT 111.825 189.975 112.055 190.475 ;
        RECT 112.430 190.395 112.600 190.595 ;
        RECT 112.225 190.225 112.600 190.395 ;
        RECT 112.770 190.225 113.320 190.425 ;
        RECT 113.490 190.145 113.735 190.595 ;
        RECT 113.905 189.975 114.075 190.935 ;
        RECT 114.245 190.695 115.915 191.785 ;
        RECT 116.635 191.105 116.805 191.615 ;
        RECT 116.975 191.275 117.305 191.785 ;
        RECT 117.475 191.105 117.645 191.615 ;
        RECT 117.815 191.275 118.145 191.785 ;
        RECT 118.315 191.105 118.485 191.615 ;
        RECT 118.770 191.275 119.440 191.785 ;
        RECT 119.795 191.445 120.885 191.615 ;
        RECT 119.795 191.105 119.965 191.445 ;
        RECT 116.635 190.935 119.965 191.105 ;
        RECT 120.215 190.765 120.545 191.265 ;
        RECT 120.715 190.945 120.885 191.445 ;
        RECT 121.150 191.395 121.485 191.615 ;
        RECT 122.490 191.405 122.845 191.785 ;
        RECT 121.150 190.775 121.405 191.395 ;
        RECT 121.655 191.235 121.885 191.275 ;
        RECT 123.015 191.235 123.265 191.615 ;
        RECT 121.655 191.035 123.265 191.235 ;
        RECT 121.655 190.945 121.840 191.035 ;
        RECT 122.430 191.025 123.265 191.035 ;
        RECT 123.515 191.005 123.765 191.785 ;
        RECT 123.935 190.935 124.195 191.615 ;
        RECT 121.995 190.835 122.325 190.865 ;
        RECT 121.995 190.775 123.795 190.835 ;
        RECT 111.825 189.805 114.075 189.975 ;
        RECT 114.245 190.005 114.995 190.525 ;
        RECT 115.165 190.175 115.915 190.695 ;
        RECT 116.605 190.145 117.280 190.765 ;
        RECT 117.510 190.145 118.215 190.765 ;
        RECT 118.415 190.145 119.125 190.765 ;
        RECT 119.715 190.595 120.545 190.765 ;
        RECT 119.365 190.145 119.535 190.475 ;
        RECT 111.485 189.465 112.440 189.635 ;
        RECT 112.855 189.235 113.185 189.625 ;
        RECT 113.355 189.485 113.525 189.805 ;
        RECT 113.695 189.235 114.025 189.625 ;
        RECT 114.245 189.235 115.915 190.005 ;
        RECT 119.715 189.975 120.030 190.595 ;
        RECT 120.725 190.425 120.950 190.775 ;
        RECT 121.150 190.665 123.855 190.775 ;
        RECT 121.150 190.605 122.325 190.665 ;
        RECT 123.655 190.630 123.855 190.665 ;
        RECT 120.280 190.225 120.950 190.425 ;
        RECT 121.145 190.225 121.635 190.425 ;
        RECT 121.825 190.225 122.300 190.435 ;
        RECT 116.555 189.805 118.565 189.975 ;
        RECT 118.755 189.805 120.965 189.975 ;
        RECT 116.975 189.235 117.305 189.615 ;
        RECT 117.815 189.445 119.535 189.615 ;
        RECT 119.715 189.405 119.885 189.805 ;
        RECT 120.135 189.235 120.465 189.615 ;
        RECT 120.635 189.445 120.965 189.805 ;
        RECT 121.150 189.235 121.605 190.000 ;
        RECT 122.080 189.825 122.300 190.225 ;
        RECT 122.545 190.225 122.875 190.435 ;
        RECT 122.545 189.825 122.755 190.225 ;
        RECT 123.045 190.190 123.455 190.495 ;
        RECT 123.685 190.055 123.855 190.630 ;
        RECT 123.585 189.935 123.855 190.055 ;
        RECT 123.010 189.890 123.855 189.935 ;
        RECT 123.010 189.765 123.765 189.890 ;
        RECT 123.010 189.615 123.180 189.765 ;
        RECT 124.025 189.745 124.195 190.935 ;
        RECT 124.365 190.695 126.955 191.785 ;
        RECT 123.965 189.735 124.195 189.745 ;
        RECT 121.880 189.405 123.180 189.615 ;
        RECT 123.435 189.235 123.765 189.595 ;
        RECT 123.935 189.405 124.195 189.735 ;
        RECT 124.365 190.005 125.575 190.525 ;
        RECT 125.745 190.175 126.955 190.695 ;
        RECT 127.125 190.620 127.415 191.785 ;
        RECT 127.585 190.935 127.845 191.615 ;
        RECT 128.015 191.005 128.265 191.785 ;
        RECT 128.515 191.235 128.765 191.615 ;
        RECT 128.935 191.405 129.290 191.785 ;
        RECT 130.295 191.395 130.630 191.615 ;
        RECT 129.895 191.235 130.125 191.275 ;
        RECT 128.515 191.035 130.125 191.235 ;
        RECT 128.515 191.025 129.350 191.035 ;
        RECT 129.940 190.945 130.125 191.035 ;
        RECT 124.365 189.235 126.955 190.005 ;
        RECT 127.125 189.235 127.415 189.960 ;
        RECT 127.585 189.735 127.755 190.935 ;
        RECT 129.455 190.835 129.785 190.865 ;
        RECT 127.985 190.775 129.785 190.835 ;
        RECT 130.375 190.775 130.630 191.395 ;
        RECT 127.925 190.665 130.630 190.775 ;
        RECT 127.925 190.630 128.125 190.665 ;
        RECT 127.925 190.055 128.095 190.630 ;
        RECT 129.455 190.605 130.630 190.665 ;
        RECT 130.805 190.710 131.075 191.615 ;
        RECT 131.245 191.025 131.575 191.785 ;
        RECT 131.755 190.855 131.925 191.615 ;
        RECT 132.185 191.350 137.530 191.785 ;
        RECT 137.705 191.350 143.050 191.785 ;
        RECT 143.225 191.350 148.570 191.785 ;
        RECT 128.325 190.190 128.735 190.495 ;
        RECT 128.905 190.225 129.235 190.435 ;
        RECT 127.925 189.935 128.195 190.055 ;
        RECT 127.925 189.890 128.770 189.935 ;
        RECT 128.015 189.765 128.770 189.890 ;
        RECT 129.025 189.825 129.235 190.225 ;
        RECT 129.480 190.225 129.955 190.435 ;
        RECT 130.145 190.225 130.635 190.425 ;
        RECT 129.480 189.825 129.700 190.225 ;
        RECT 127.585 189.405 127.845 189.735 ;
        RECT 128.600 189.615 128.770 189.765 ;
        RECT 128.015 189.235 128.345 189.595 ;
        RECT 128.600 189.405 129.900 189.615 ;
        RECT 130.175 189.235 130.630 190.000 ;
        RECT 130.805 189.910 130.975 190.710 ;
        RECT 131.260 190.685 131.925 190.855 ;
        RECT 131.260 190.540 131.430 190.685 ;
        RECT 131.145 190.210 131.430 190.540 ;
        RECT 131.260 189.955 131.430 190.210 ;
        RECT 131.665 190.135 131.995 190.505 ;
        RECT 130.805 189.405 131.065 189.910 ;
        RECT 131.260 189.785 131.925 189.955 ;
        RECT 131.245 189.235 131.575 189.615 ;
        RECT 131.755 189.405 131.925 189.785 ;
        RECT 133.770 189.780 134.110 190.610 ;
        RECT 135.590 190.100 135.940 191.350 ;
        RECT 139.290 189.780 139.630 190.610 ;
        RECT 141.110 190.100 141.460 191.350 ;
        RECT 144.810 189.780 145.150 190.610 ;
        RECT 146.630 190.100 146.980 191.350 ;
        RECT 149.205 190.695 150.415 191.785 ;
        RECT 149.205 190.155 149.725 190.695 ;
        RECT 149.895 189.985 150.415 190.525 ;
        RECT 132.185 189.235 137.530 189.780 ;
        RECT 137.705 189.235 143.050 189.780 ;
        RECT 143.225 189.235 148.570 189.780 ;
        RECT 149.205 189.235 150.415 189.985 ;
        RECT 11.120 189.065 150.500 189.235 ;
        RECT 11.205 188.315 12.415 189.065 ;
        RECT 12.585 188.315 13.795 189.065 ;
        RECT 13.985 188.375 14.225 188.895 ;
        RECT 14.395 188.570 14.790 189.065 ;
        RECT 15.355 188.735 15.525 188.880 ;
        RECT 15.150 188.540 15.525 188.735 ;
        RECT 11.205 187.775 11.725 188.315 ;
        RECT 11.895 187.605 12.415 188.145 ;
        RECT 12.585 187.775 13.105 188.315 ;
        RECT 13.275 187.605 13.795 188.145 ;
        RECT 11.205 186.515 12.415 187.605 ;
        RECT 12.585 186.515 13.795 187.605 ;
        RECT 13.985 187.570 14.160 188.375 ;
        RECT 15.150 188.205 15.320 188.540 ;
        RECT 15.805 188.495 16.045 188.870 ;
        RECT 16.215 188.560 16.550 189.065 ;
        RECT 17.185 188.685 18.075 188.855 ;
        RECT 15.805 188.345 16.025 188.495 ;
        RECT 14.335 187.845 15.320 188.205 ;
        RECT 15.490 188.015 16.025 188.345 ;
        RECT 14.335 187.825 15.620 187.845 ;
        RECT 14.760 187.675 15.620 187.825 ;
        RECT 13.985 186.785 14.290 187.570 ;
        RECT 14.465 187.195 15.160 187.505 ;
        RECT 14.470 186.515 15.155 186.985 ;
        RECT 15.335 186.730 15.620 187.675 ;
        RECT 15.790 187.365 16.025 188.015 ;
        RECT 16.195 187.535 16.495 188.385 ;
        RECT 17.185 188.130 17.735 188.515 ;
        RECT 17.905 187.960 18.075 188.685 ;
        RECT 17.185 187.890 18.075 187.960 ;
        RECT 18.245 188.385 18.465 188.845 ;
        RECT 18.635 188.525 18.885 189.065 ;
        RECT 19.055 188.415 19.315 188.895 ;
        RECT 18.245 188.360 18.495 188.385 ;
        RECT 18.245 187.935 18.575 188.360 ;
        RECT 17.185 187.865 18.080 187.890 ;
        RECT 17.185 187.850 18.090 187.865 ;
        RECT 17.185 187.835 18.095 187.850 ;
        RECT 17.185 187.830 18.105 187.835 ;
        RECT 17.185 187.820 18.110 187.830 ;
        RECT 17.185 187.810 18.115 187.820 ;
        RECT 17.185 187.805 18.125 187.810 ;
        RECT 17.185 187.795 18.135 187.805 ;
        RECT 17.185 187.790 18.145 187.795 ;
        RECT 15.790 187.135 16.465 187.365 ;
        RECT 17.185 187.340 17.445 187.790 ;
        RECT 17.810 187.785 18.145 187.790 ;
        RECT 17.810 187.780 18.160 187.785 ;
        RECT 17.810 187.770 18.175 187.780 ;
        RECT 17.810 187.765 18.200 187.770 ;
        RECT 18.745 187.765 18.975 188.160 ;
        RECT 17.810 187.760 18.975 187.765 ;
        RECT 17.840 187.725 18.975 187.760 ;
        RECT 17.875 187.700 18.975 187.725 ;
        RECT 17.905 187.670 18.975 187.700 ;
        RECT 17.925 187.640 18.975 187.670 ;
        RECT 17.945 187.610 18.975 187.640 ;
        RECT 18.015 187.600 18.975 187.610 ;
        RECT 18.040 187.590 18.975 187.600 ;
        RECT 18.060 187.575 18.975 187.590 ;
        RECT 18.080 187.560 18.975 187.575 ;
        RECT 18.085 187.550 18.870 187.560 ;
        RECT 18.100 187.515 18.870 187.550 ;
        RECT 17.615 187.195 17.945 187.440 ;
        RECT 18.115 187.265 18.870 187.515 ;
        RECT 19.145 187.385 19.315 188.415 ;
        RECT 19.485 188.295 22.995 189.065 ;
        RECT 23.625 188.685 24.515 188.855 ;
        RECT 19.485 187.775 21.135 188.295 ;
        RECT 23.625 188.130 24.175 188.515 ;
        RECT 21.305 187.605 22.995 188.125 ;
        RECT 24.345 187.960 24.515 188.685 ;
        RECT 17.615 187.170 17.800 187.195 ;
        RECT 15.795 186.515 16.125 186.965 ;
        RECT 16.295 186.705 16.465 187.135 ;
        RECT 17.185 187.070 17.800 187.170 ;
        RECT 17.185 186.515 17.790 187.070 ;
        RECT 17.965 186.685 18.445 187.025 ;
        RECT 18.615 186.515 18.870 187.060 ;
        RECT 19.040 186.685 19.315 187.385 ;
        RECT 19.485 186.515 22.995 187.605 ;
        RECT 23.625 187.890 24.515 187.960 ;
        RECT 24.685 188.360 24.905 188.845 ;
        RECT 25.075 188.525 25.325 189.065 ;
        RECT 25.495 188.415 25.755 188.895 ;
        RECT 24.685 187.935 25.015 188.360 ;
        RECT 23.625 187.865 24.520 187.890 ;
        RECT 23.625 187.850 24.530 187.865 ;
        RECT 23.625 187.835 24.535 187.850 ;
        RECT 23.625 187.830 24.545 187.835 ;
        RECT 23.625 187.820 24.550 187.830 ;
        RECT 23.625 187.810 24.555 187.820 ;
        RECT 23.625 187.805 24.565 187.810 ;
        RECT 23.625 187.795 24.575 187.805 ;
        RECT 23.625 187.790 24.585 187.795 ;
        RECT 23.625 187.340 23.885 187.790 ;
        RECT 24.250 187.785 24.585 187.790 ;
        RECT 24.250 187.780 24.600 187.785 ;
        RECT 24.250 187.770 24.615 187.780 ;
        RECT 24.250 187.765 24.640 187.770 ;
        RECT 25.185 187.765 25.415 188.160 ;
        RECT 24.250 187.760 25.415 187.765 ;
        RECT 24.280 187.725 25.415 187.760 ;
        RECT 24.315 187.700 25.415 187.725 ;
        RECT 24.345 187.670 25.415 187.700 ;
        RECT 24.365 187.640 25.415 187.670 ;
        RECT 24.385 187.610 25.415 187.640 ;
        RECT 24.455 187.600 25.415 187.610 ;
        RECT 24.480 187.590 25.415 187.600 ;
        RECT 24.500 187.575 25.415 187.590 ;
        RECT 24.520 187.560 25.415 187.575 ;
        RECT 24.525 187.550 25.310 187.560 ;
        RECT 24.540 187.515 25.310 187.550 ;
        RECT 24.055 187.195 24.385 187.440 ;
        RECT 24.555 187.265 25.310 187.515 ;
        RECT 25.585 187.385 25.755 188.415 ;
        RECT 24.055 187.170 24.240 187.195 ;
        RECT 23.625 187.070 24.240 187.170 ;
        RECT 23.625 186.515 24.230 187.070 ;
        RECT 24.405 186.685 24.885 187.025 ;
        RECT 25.055 186.515 25.310 187.060 ;
        RECT 25.480 186.685 25.755 187.385 ;
        RECT 25.925 188.390 26.185 188.895 ;
        RECT 26.365 188.685 26.695 189.065 ;
        RECT 26.875 188.515 27.045 188.895 ;
        RECT 25.925 187.590 26.095 188.390 ;
        RECT 26.380 188.345 27.045 188.515 ;
        RECT 26.380 188.090 26.550 188.345 ;
        RECT 27.305 188.295 29.895 189.065 ;
        RECT 26.265 187.760 26.550 188.090 ;
        RECT 26.785 187.795 27.115 188.165 ;
        RECT 27.305 187.775 28.515 188.295 ;
        RECT 30.525 188.265 30.835 189.065 ;
        RECT 31.040 188.265 31.735 188.895 ;
        RECT 31.905 188.295 35.415 189.065 ;
        RECT 35.585 188.315 36.795 189.065 ;
        RECT 36.965 188.340 37.255 189.065 ;
        RECT 26.380 187.615 26.550 187.760 ;
        RECT 25.925 186.685 26.195 187.590 ;
        RECT 26.380 187.445 27.045 187.615 ;
        RECT 28.685 187.605 29.895 188.125 ;
        RECT 30.535 187.825 30.870 188.095 ;
        RECT 31.040 187.665 31.210 188.265 ;
        RECT 31.380 187.825 31.715 188.075 ;
        RECT 31.905 187.775 33.555 188.295 ;
        RECT 26.365 186.515 26.695 187.275 ;
        RECT 26.875 186.685 27.045 187.445 ;
        RECT 27.305 186.515 29.895 187.605 ;
        RECT 30.525 186.515 30.805 187.655 ;
        RECT 30.975 186.685 31.305 187.665 ;
        RECT 31.475 186.515 31.735 187.655 ;
        RECT 33.725 187.605 35.415 188.125 ;
        RECT 35.585 187.775 36.105 188.315 ;
        RECT 37.425 188.295 40.015 189.065 ;
        RECT 40.645 188.325 41.110 188.870 ;
        RECT 36.275 187.605 36.795 188.145 ;
        RECT 37.425 187.775 38.635 188.295 ;
        RECT 31.905 186.515 35.415 187.605 ;
        RECT 35.585 186.515 36.795 187.605 ;
        RECT 36.965 186.515 37.255 187.680 ;
        RECT 38.805 187.605 40.015 188.125 ;
        RECT 37.425 186.515 40.015 187.605 ;
        RECT 40.645 187.365 40.815 188.325 ;
        RECT 41.615 188.245 41.785 189.065 ;
        RECT 41.955 188.415 42.285 188.895 ;
        RECT 42.455 188.675 42.805 189.065 ;
        RECT 42.975 188.495 43.205 188.895 ;
        RECT 42.695 188.415 43.205 188.495 ;
        RECT 41.955 188.325 43.205 188.415 ;
        RECT 43.375 188.325 43.695 188.805 ;
        RECT 43.865 188.520 49.210 189.065 ;
        RECT 41.955 188.245 42.865 188.325 ;
        RECT 40.985 187.705 41.230 188.155 ;
        RECT 41.490 187.875 42.185 188.075 ;
        RECT 42.355 187.905 42.955 188.075 ;
        RECT 42.355 187.705 42.525 187.905 ;
        RECT 43.185 187.735 43.355 188.155 ;
        RECT 40.985 187.535 42.525 187.705 ;
        RECT 42.695 187.565 43.355 187.735 ;
        RECT 42.695 187.365 42.865 187.565 ;
        RECT 43.525 187.395 43.695 188.325 ;
        RECT 45.450 187.690 45.790 188.520 ;
        RECT 49.445 188.245 49.655 189.065 ;
        RECT 49.825 188.265 50.155 188.895 ;
        RECT 40.645 187.195 42.865 187.365 ;
        RECT 43.035 187.195 43.695 187.395 ;
        RECT 40.645 186.515 40.945 187.025 ;
        RECT 41.115 186.685 41.445 187.195 ;
        RECT 43.035 187.025 43.205 187.195 ;
        RECT 41.615 186.515 42.245 187.025 ;
        RECT 42.825 186.855 43.205 187.025 ;
        RECT 43.375 186.515 43.675 187.025 ;
        RECT 47.270 186.950 47.620 188.200 ;
        RECT 49.825 187.665 50.075 188.265 ;
        RECT 50.325 188.245 50.555 189.065 ;
        RECT 51.685 188.265 51.995 189.065 ;
        RECT 52.200 188.265 52.895 188.895 ;
        RECT 53.065 188.685 53.955 188.855 ;
        RECT 50.245 187.825 50.575 188.075 ;
        RECT 51.695 187.825 52.030 188.095 ;
        RECT 52.200 187.665 52.370 188.265 ;
        RECT 53.065 188.130 53.615 188.515 ;
        RECT 52.540 187.825 52.875 188.075 ;
        RECT 53.785 187.960 53.955 188.685 ;
        RECT 53.065 187.890 53.955 187.960 ;
        RECT 54.125 188.360 54.345 188.845 ;
        RECT 54.515 188.525 54.765 189.065 ;
        RECT 54.935 188.415 55.195 188.895 ;
        RECT 54.125 187.935 54.455 188.360 ;
        RECT 53.065 187.865 53.960 187.890 ;
        RECT 53.065 187.850 53.970 187.865 ;
        RECT 53.065 187.835 53.975 187.850 ;
        RECT 53.065 187.830 53.985 187.835 ;
        RECT 53.065 187.820 53.990 187.830 ;
        RECT 53.065 187.810 53.995 187.820 ;
        RECT 53.065 187.805 54.005 187.810 ;
        RECT 53.065 187.795 54.015 187.805 ;
        RECT 53.065 187.790 54.025 187.795 ;
        RECT 43.865 186.515 49.210 186.950 ;
        RECT 49.445 186.515 49.655 187.655 ;
        RECT 49.825 186.685 50.155 187.665 ;
        RECT 50.325 186.515 50.555 187.655 ;
        RECT 51.685 186.515 51.965 187.655 ;
        RECT 52.135 186.685 52.465 187.665 ;
        RECT 52.635 186.515 52.895 187.655 ;
        RECT 53.065 187.340 53.325 187.790 ;
        RECT 53.690 187.785 54.025 187.790 ;
        RECT 53.690 187.780 54.040 187.785 ;
        RECT 53.690 187.770 54.055 187.780 ;
        RECT 53.690 187.765 54.080 187.770 ;
        RECT 54.625 187.765 54.855 188.160 ;
        RECT 53.690 187.760 54.855 187.765 ;
        RECT 53.720 187.725 54.855 187.760 ;
        RECT 53.755 187.700 54.855 187.725 ;
        RECT 53.785 187.670 54.855 187.700 ;
        RECT 53.805 187.640 54.855 187.670 ;
        RECT 53.825 187.610 54.855 187.640 ;
        RECT 53.895 187.600 54.855 187.610 ;
        RECT 53.920 187.590 54.855 187.600 ;
        RECT 53.940 187.575 54.855 187.590 ;
        RECT 53.960 187.560 54.855 187.575 ;
        RECT 53.965 187.550 54.750 187.560 ;
        RECT 53.980 187.515 54.750 187.550 ;
        RECT 53.495 187.195 53.825 187.440 ;
        RECT 53.995 187.265 54.750 187.515 ;
        RECT 55.025 187.385 55.195 188.415 ;
        RECT 55.455 188.515 55.625 188.805 ;
        RECT 55.795 188.685 56.125 189.065 ;
        RECT 55.455 188.345 56.120 188.515 ;
        RECT 55.370 187.525 55.720 188.175 ;
        RECT 53.495 187.170 53.680 187.195 ;
        RECT 53.065 187.070 53.680 187.170 ;
        RECT 53.065 186.515 53.670 187.070 ;
        RECT 53.845 186.685 54.325 187.025 ;
        RECT 54.495 186.515 54.750 187.060 ;
        RECT 54.920 186.685 55.195 187.385 ;
        RECT 55.890 187.355 56.120 188.345 ;
        RECT 55.455 187.185 56.120 187.355 ;
        RECT 55.455 186.685 55.625 187.185 ;
        RECT 55.795 186.515 56.125 187.015 ;
        RECT 56.295 186.685 56.480 188.805 ;
        RECT 56.735 188.605 56.985 189.065 ;
        RECT 57.155 188.615 57.490 188.785 ;
        RECT 57.685 188.615 58.360 188.785 ;
        RECT 57.155 188.475 57.325 188.615 ;
        RECT 56.650 187.485 56.930 188.435 ;
        RECT 57.100 188.345 57.325 188.475 ;
        RECT 57.100 187.240 57.270 188.345 ;
        RECT 57.495 188.195 58.020 188.415 ;
        RECT 57.440 187.430 57.680 188.025 ;
        RECT 57.850 187.495 58.020 188.195 ;
        RECT 58.190 187.835 58.360 188.615 ;
        RECT 58.680 188.565 59.050 189.065 ;
        RECT 59.230 188.615 59.635 188.785 ;
        RECT 59.805 188.615 60.590 188.785 ;
        RECT 59.230 188.385 59.400 188.615 ;
        RECT 58.570 188.085 59.400 188.385 ;
        RECT 59.785 188.115 60.250 188.445 ;
        RECT 58.570 188.055 58.770 188.085 ;
        RECT 58.890 187.835 59.060 187.905 ;
        RECT 58.190 187.665 59.060 187.835 ;
        RECT 58.550 187.575 59.060 187.665 ;
        RECT 57.100 187.110 57.405 187.240 ;
        RECT 57.850 187.130 58.380 187.495 ;
        RECT 56.720 186.515 56.985 186.975 ;
        RECT 57.155 186.685 57.405 187.110 ;
        RECT 58.550 186.960 58.720 187.575 ;
        RECT 57.615 186.790 58.720 186.960 ;
        RECT 58.890 186.515 59.060 187.315 ;
        RECT 59.230 187.015 59.400 188.085 ;
        RECT 59.570 187.185 59.760 187.905 ;
        RECT 59.930 187.155 60.250 188.115 ;
        RECT 60.420 188.155 60.590 188.615 ;
        RECT 60.865 188.535 61.075 189.065 ;
        RECT 61.335 188.325 61.665 188.850 ;
        RECT 61.835 188.455 62.005 189.065 ;
        RECT 62.175 188.410 62.505 188.845 ;
        RECT 62.175 188.325 62.555 188.410 ;
        RECT 62.725 188.340 63.015 189.065 ;
        RECT 63.190 188.810 63.525 188.855 ;
        RECT 63.185 188.345 63.525 188.810 ;
        RECT 63.695 188.685 64.025 189.065 ;
        RECT 61.465 188.155 61.665 188.325 ;
        RECT 62.330 188.285 62.555 188.325 ;
        RECT 60.420 187.825 61.295 188.155 ;
        RECT 61.465 187.825 62.215 188.155 ;
        RECT 59.230 186.685 59.480 187.015 ;
        RECT 60.420 186.985 60.590 187.825 ;
        RECT 61.465 187.620 61.655 187.825 ;
        RECT 62.385 187.705 62.555 188.285 ;
        RECT 62.340 187.655 62.555 187.705 ;
        RECT 60.760 187.245 61.655 187.620 ;
        RECT 62.165 187.575 62.555 187.655 ;
        RECT 59.705 186.815 60.590 186.985 ;
        RECT 60.770 186.515 61.085 187.015 ;
        RECT 61.315 186.685 61.655 187.245 ;
        RECT 61.825 186.515 61.995 187.525 ;
        RECT 62.165 186.730 62.495 187.575 ;
        RECT 62.725 186.515 63.015 187.680 ;
        RECT 63.185 187.655 63.355 188.345 ;
        RECT 63.525 187.825 63.785 188.155 ;
        RECT 63.185 186.685 63.445 187.655 ;
        RECT 63.615 187.275 63.785 187.825 ;
        RECT 63.955 187.455 64.295 188.485 ;
        RECT 64.485 188.045 64.755 188.730 ;
        RECT 64.485 187.875 64.795 188.045 ;
        RECT 64.485 187.455 64.755 187.875 ;
        RECT 64.980 187.455 65.260 188.730 ;
        RECT 65.460 188.565 65.690 188.895 ;
        RECT 65.935 188.685 66.265 189.065 ;
        RECT 65.460 187.275 65.630 188.565 ;
        RECT 66.435 188.495 66.610 188.895 ;
        RECT 65.980 188.325 66.610 188.495 ;
        RECT 67.875 188.415 68.045 188.895 ;
        RECT 68.215 188.585 68.545 189.065 ;
        RECT 68.770 188.645 70.305 188.895 ;
        RECT 68.770 188.415 68.940 188.645 ;
        RECT 65.980 188.155 66.150 188.325 ;
        RECT 67.875 188.245 68.940 188.415 ;
        RECT 65.800 187.825 66.150 188.155 ;
        RECT 63.615 187.105 65.630 187.275 ;
        RECT 65.980 187.305 66.150 187.825 ;
        RECT 66.330 187.475 66.695 188.155 ;
        RECT 69.120 188.075 69.400 188.475 ;
        RECT 67.790 187.865 68.140 188.075 ;
        RECT 68.310 187.875 68.755 188.075 ;
        RECT 68.925 187.875 69.400 188.075 ;
        RECT 69.670 188.075 69.955 188.475 ;
        RECT 70.135 188.415 70.305 188.645 ;
        RECT 70.475 188.585 70.805 189.065 ;
        RECT 71.020 188.565 71.275 188.895 ;
        RECT 71.475 188.565 71.805 189.065 ;
        RECT 71.090 188.485 71.275 188.565 ;
        RECT 70.135 188.245 70.935 188.415 ;
        RECT 69.670 187.875 70.000 188.075 ;
        RECT 70.170 187.875 70.535 188.075 ;
        RECT 70.765 187.695 70.935 188.245 ;
        RECT 67.875 187.525 70.935 187.695 ;
        RECT 65.980 187.135 66.610 187.305 ;
        RECT 63.640 186.515 63.970 186.925 ;
        RECT 64.170 186.685 64.340 187.105 ;
        RECT 64.555 186.515 65.225 186.925 ;
        RECT 65.460 186.685 65.630 187.105 ;
        RECT 65.935 186.515 66.265 186.955 ;
        RECT 66.435 186.685 66.610 187.135 ;
        RECT 67.875 186.685 68.045 187.525 ;
        RECT 71.105 187.365 71.275 188.485 ;
        RECT 72.005 188.495 72.175 188.845 ;
        RECT 72.375 188.665 72.705 189.065 ;
        RECT 72.875 188.495 73.045 188.845 ;
        RECT 73.215 188.665 73.595 189.065 ;
        RECT 71.470 187.825 71.820 188.395 ;
        RECT 72.005 188.325 73.615 188.495 ;
        RECT 73.785 188.390 74.055 188.735 ;
        RECT 73.445 188.155 73.615 188.325 ;
        RECT 71.065 187.355 71.275 187.365 ;
        RECT 68.215 186.855 68.545 187.355 ;
        RECT 68.715 187.115 70.350 187.355 ;
        RECT 68.715 187.025 68.945 187.115 ;
        RECT 69.055 186.855 69.385 186.895 ;
        RECT 68.215 186.685 69.385 186.855 ;
        RECT 69.575 186.515 69.930 186.935 ;
        RECT 70.100 186.685 70.350 187.115 ;
        RECT 70.520 186.515 70.850 187.275 ;
        RECT 71.020 186.685 71.275 187.355 ;
        RECT 71.470 187.365 71.790 187.655 ;
        RECT 71.990 187.535 72.700 188.155 ;
        RECT 72.870 187.825 73.275 188.155 ;
        RECT 73.445 187.825 73.715 188.155 ;
        RECT 73.445 187.655 73.615 187.825 ;
        RECT 73.885 187.655 74.055 188.390 ;
        RECT 74.245 188.255 74.485 189.065 ;
        RECT 74.655 188.255 74.985 188.895 ;
        RECT 75.155 188.255 75.425 189.065 ;
        RECT 76.075 188.665 76.405 189.065 ;
        RECT 76.575 188.495 76.745 188.765 ;
        RECT 76.915 188.665 77.245 189.065 ;
        RECT 77.420 188.505 77.685 188.765 ;
        RECT 77.935 188.575 78.195 189.065 ;
        RECT 77.420 188.495 77.775 188.505 ;
        RECT 74.225 187.825 74.575 188.075 ;
        RECT 74.745 187.655 74.915 188.255 ;
        RECT 75.085 187.825 75.435 188.075 ;
        RECT 72.890 187.485 73.615 187.655 ;
        RECT 72.890 187.365 73.060 187.485 ;
        RECT 71.470 187.195 73.060 187.365 ;
        RECT 71.470 186.735 73.125 187.025 ;
        RECT 73.295 186.515 73.575 187.315 ;
        RECT 73.785 186.685 74.055 187.655 ;
        RECT 74.235 187.485 74.915 187.655 ;
        RECT 74.235 186.700 74.565 187.485 ;
        RECT 75.095 186.515 75.425 187.655 ;
        RECT 76.065 187.485 76.325 188.495 ;
        RECT 76.575 188.325 77.775 188.495 ;
        RECT 76.585 187.905 77.035 188.075 ;
        RECT 76.065 186.515 76.325 187.315 ;
        RECT 76.585 186.700 76.825 187.905 ;
        RECT 77.205 187.735 77.435 188.155 ;
        RECT 76.995 187.535 77.435 187.735 ;
        RECT 77.605 187.655 77.775 188.325 ;
        RECT 77.945 187.825 78.195 188.405 ;
        RECT 79.285 188.390 79.560 188.735 ;
        RECT 79.750 188.665 80.130 189.065 ;
        RECT 80.300 188.495 80.470 188.845 ;
        RECT 80.640 188.665 80.970 189.065 ;
        RECT 81.145 188.495 81.315 188.845 ;
        RECT 81.515 188.565 81.845 189.065 ;
        RECT 79.285 187.655 79.455 188.390 ;
        RECT 79.730 188.325 81.315 188.495 ;
        RECT 79.730 188.155 79.900 188.325 ;
        RECT 82.040 188.155 82.285 188.845 ;
        RECT 82.455 188.565 82.795 189.065 ;
        RECT 82.985 188.580 83.775 188.845 ;
        RECT 79.625 187.825 79.900 188.155 ;
        RECT 80.070 187.825 80.450 188.155 ;
        RECT 79.730 187.655 79.900 187.825 ;
        RECT 76.995 186.700 77.250 187.535 ;
        RECT 77.605 187.485 78.190 187.655 ;
        RECT 77.855 186.700 78.190 187.485 ;
        RECT 79.285 186.685 79.560 187.655 ;
        RECT 79.730 187.485 80.390 187.655 ;
        RECT 80.620 187.535 81.360 188.155 ;
        RECT 81.630 187.825 82.285 188.155 ;
        RECT 82.455 187.825 82.795 188.395 ;
        RECT 82.965 187.905 83.350 188.385 ;
        RECT 80.220 187.365 80.390 187.485 ;
        RECT 81.530 187.365 81.850 187.655 ;
        RECT 79.770 186.515 80.050 187.315 ;
        RECT 80.220 187.195 81.850 187.365 ;
        RECT 82.045 187.230 82.285 187.825 ;
        RECT 83.520 187.725 83.775 188.580 ;
        RECT 83.945 188.400 84.175 188.845 ;
        RECT 84.355 188.570 84.685 189.065 ;
        RECT 84.860 188.435 85.110 188.895 ;
        RECT 83.945 187.905 84.355 188.400 ;
        RECT 84.940 188.225 85.110 188.435 ;
        RECT 85.280 188.405 85.555 189.065 ;
        RECT 85.725 188.315 86.935 189.065 ;
        RECT 84.540 187.725 84.770 188.155 ;
        RECT 80.220 186.855 82.275 187.025 ;
        RECT 80.220 186.735 82.270 186.855 ;
        RECT 82.455 186.515 82.795 187.590 ;
        RECT 82.980 187.555 84.770 187.725 ;
        RECT 84.940 187.705 85.555 188.225 ;
        RECT 85.725 187.775 86.245 188.315 ;
        RECT 87.165 188.245 87.375 189.065 ;
        RECT 87.545 188.265 87.875 188.895 ;
        RECT 82.980 187.190 83.235 187.555 ;
        RECT 83.405 187.195 83.735 187.385 ;
        RECT 83.960 187.260 84.210 187.555 ;
        RECT 83.405 187.020 83.595 187.195 ;
        RECT 82.965 186.515 83.595 187.020 ;
        RECT 83.775 186.685 84.250 187.025 ;
        RECT 84.435 186.515 84.650 187.360 ;
        RECT 84.955 187.355 85.125 187.705 ;
        RECT 86.415 187.605 86.935 188.145 ;
        RECT 87.545 187.665 87.795 188.265 ;
        RECT 88.045 188.245 88.275 189.065 ;
        RECT 88.485 188.340 88.775 189.065 ;
        RECT 88.945 188.295 90.615 189.065 ;
        RECT 87.965 187.825 88.295 188.075 ;
        RECT 88.945 187.775 89.695 188.295 ;
        RECT 84.850 186.685 85.125 187.355 ;
        RECT 85.295 186.515 85.555 187.525 ;
        RECT 85.725 186.515 86.935 187.605 ;
        RECT 87.165 186.515 87.375 187.655 ;
        RECT 87.545 186.685 87.875 187.665 ;
        RECT 88.045 186.515 88.275 187.655 ;
        RECT 88.485 186.515 88.775 187.680 ;
        RECT 89.865 187.605 90.615 188.125 ;
        RECT 88.945 186.515 90.615 187.605 ;
        RECT 91.245 186.685 91.525 188.785 ;
        RECT 91.755 188.605 91.925 189.065 ;
        RECT 92.195 188.675 93.445 188.855 ;
        RECT 92.580 188.435 92.945 188.505 ;
        RECT 91.695 188.255 92.945 188.435 ;
        RECT 93.115 188.455 93.445 188.675 ;
        RECT 93.615 188.625 93.785 189.065 ;
        RECT 93.955 188.455 94.295 188.870 ;
        RECT 93.115 188.285 94.295 188.455 ;
        RECT 91.695 187.655 91.970 188.255 ;
        RECT 94.505 188.245 94.735 189.065 ;
        RECT 94.905 188.265 95.235 188.895 ;
        RECT 92.140 187.825 92.495 188.075 ;
        RECT 92.690 187.825 93.155 188.075 ;
        RECT 93.325 187.825 93.655 188.075 ;
        RECT 93.830 187.875 94.295 188.075 ;
        RECT 94.485 187.825 94.815 188.075 ;
        RECT 93.475 187.705 93.655 187.825 ;
        RECT 91.695 187.445 93.305 187.655 ;
        RECT 93.475 187.535 93.805 187.705 ;
        RECT 92.895 187.345 93.305 187.445 ;
        RECT 91.715 186.515 92.500 187.275 ;
        RECT 92.895 186.685 93.280 187.345 ;
        RECT 93.605 186.745 93.805 187.535 ;
        RECT 93.975 186.515 94.295 187.695 ;
        RECT 94.985 187.665 95.235 188.265 ;
        RECT 95.405 188.245 95.615 189.065 ;
        RECT 96.305 188.390 96.575 188.735 ;
        RECT 96.765 188.665 97.145 189.065 ;
        RECT 97.315 188.495 97.485 188.845 ;
        RECT 97.655 188.665 97.985 189.065 ;
        RECT 98.185 188.495 98.355 188.845 ;
        RECT 98.555 188.565 98.885 189.065 ;
        RECT 94.505 186.515 94.735 187.655 ;
        RECT 94.905 186.685 95.235 187.665 ;
        RECT 96.305 187.655 96.475 188.390 ;
        RECT 96.745 188.325 98.355 188.495 ;
        RECT 96.745 188.155 96.915 188.325 ;
        RECT 96.645 187.825 96.915 188.155 ;
        RECT 97.085 187.825 97.490 188.155 ;
        RECT 96.745 187.655 96.915 187.825 ;
        RECT 95.405 186.515 95.615 187.655 ;
        RECT 96.305 186.685 96.575 187.655 ;
        RECT 96.745 187.485 97.470 187.655 ;
        RECT 97.660 187.535 98.370 188.155 ;
        RECT 98.540 187.825 98.890 188.395 ;
        RECT 99.065 188.315 100.275 189.065 ;
        RECT 100.465 188.565 100.720 188.895 ;
        RECT 100.935 188.585 101.265 189.065 ;
        RECT 101.435 188.645 102.970 188.895 ;
        RECT 100.465 188.555 100.675 188.565 ;
        RECT 100.465 188.485 100.650 188.555 ;
        RECT 99.065 187.775 99.585 188.315 ;
        RECT 97.300 187.365 97.470 187.485 ;
        RECT 98.570 187.365 98.890 187.655 ;
        RECT 99.755 187.605 100.275 188.145 ;
        RECT 96.785 186.515 97.065 187.315 ;
        RECT 97.300 187.195 98.890 187.365 ;
        RECT 97.235 186.735 98.890 187.025 ;
        RECT 99.065 186.515 100.275 187.605 ;
        RECT 100.465 187.355 100.635 188.485 ;
        RECT 101.435 188.415 101.605 188.645 ;
        RECT 100.805 188.245 101.605 188.415 ;
        RECT 100.805 187.695 100.975 188.245 ;
        RECT 101.785 188.075 102.070 188.475 ;
        RECT 101.205 188.045 101.570 188.075 ;
        RECT 101.195 187.875 101.570 188.045 ;
        RECT 101.740 187.875 102.070 188.075 ;
        RECT 102.340 188.075 102.620 188.475 ;
        RECT 102.800 188.415 102.970 188.645 ;
        RECT 103.195 188.585 103.525 189.065 ;
        RECT 103.695 188.415 103.865 188.895 ;
        RECT 102.800 188.245 103.865 188.415 ;
        RECT 104.125 188.315 105.335 189.065 ;
        RECT 102.340 187.875 102.815 188.075 ;
        RECT 102.985 187.875 103.430 188.075 ;
        RECT 103.600 187.865 103.950 188.075 ;
        RECT 104.125 187.775 104.645 188.315 ;
        RECT 105.565 188.245 105.775 189.065 ;
        RECT 105.945 188.265 106.275 188.895 ;
        RECT 100.805 187.525 103.865 187.695 ;
        RECT 104.815 187.605 105.335 188.145 ;
        RECT 105.945 187.665 106.195 188.265 ;
        RECT 106.445 188.245 106.675 189.065 ;
        RECT 106.885 188.520 112.230 189.065 ;
        RECT 106.365 187.825 106.695 188.075 ;
        RECT 108.470 187.690 108.810 188.520 ;
        RECT 112.405 188.295 114.075 189.065 ;
        RECT 114.245 188.340 114.535 189.065 ;
        RECT 114.790 188.565 115.285 188.895 ;
        RECT 100.465 186.685 100.720 187.355 ;
        RECT 100.890 186.515 101.220 187.275 ;
        RECT 101.390 187.115 103.025 187.355 ;
        RECT 101.390 186.685 101.640 187.115 ;
        RECT 102.795 187.025 103.025 187.115 ;
        RECT 101.810 186.515 102.165 186.935 ;
        RECT 102.355 186.855 102.685 186.895 ;
        RECT 103.195 186.855 103.525 187.355 ;
        RECT 102.355 186.685 103.525 186.855 ;
        RECT 103.695 186.685 103.865 187.525 ;
        RECT 104.125 186.515 105.335 187.605 ;
        RECT 105.565 186.515 105.775 187.655 ;
        RECT 105.945 186.685 106.275 187.665 ;
        RECT 106.445 186.515 106.675 187.655 ;
        RECT 110.290 186.950 110.640 188.200 ;
        RECT 112.405 187.775 113.155 188.295 ;
        RECT 113.325 187.605 114.075 188.125 ;
        RECT 106.885 186.515 112.230 186.950 ;
        RECT 112.405 186.515 114.075 187.605 ;
        RECT 114.245 186.515 114.535 187.680 ;
        RECT 114.705 187.075 114.945 188.385 ;
        RECT 115.115 187.655 115.285 188.565 ;
        RECT 115.505 187.825 115.855 188.790 ;
        RECT 116.035 187.825 116.335 188.795 ;
        RECT 116.515 187.825 116.795 188.795 ;
        RECT 116.975 188.265 117.245 189.065 ;
        RECT 117.415 188.345 117.755 188.855 ;
        RECT 117.925 188.520 123.270 189.065 ;
        RECT 123.445 188.520 128.790 189.065 ;
        RECT 128.965 188.520 134.310 189.065 ;
        RECT 134.485 188.520 139.830 189.065 ;
        RECT 116.990 187.825 117.320 188.075 ;
        RECT 116.990 187.655 117.305 187.825 ;
        RECT 115.115 187.485 117.305 187.655 ;
        RECT 114.710 186.515 115.045 186.895 ;
        RECT 115.215 186.685 115.465 187.485 ;
        RECT 115.685 186.515 116.015 187.235 ;
        RECT 116.200 186.685 116.450 187.485 ;
        RECT 116.915 186.515 117.245 187.315 ;
        RECT 117.495 186.945 117.755 188.345 ;
        RECT 119.510 187.690 119.850 188.520 ;
        RECT 121.330 186.950 121.680 188.200 ;
        RECT 125.030 187.690 125.370 188.520 ;
        RECT 126.850 186.950 127.200 188.200 ;
        RECT 130.550 187.690 130.890 188.520 ;
        RECT 132.370 186.950 132.720 188.200 ;
        RECT 136.070 187.690 136.410 188.520 ;
        RECT 140.005 188.340 140.295 189.065 ;
        RECT 140.465 188.520 145.810 189.065 ;
        RECT 137.890 186.950 138.240 188.200 ;
        RECT 142.050 187.690 142.390 188.520 ;
        RECT 145.985 188.295 148.575 189.065 ;
        RECT 149.205 188.315 150.415 189.065 ;
        RECT 117.415 186.685 117.755 186.945 ;
        RECT 117.925 186.515 123.270 186.950 ;
        RECT 123.445 186.515 128.790 186.950 ;
        RECT 128.965 186.515 134.310 186.950 ;
        RECT 134.485 186.515 139.830 186.950 ;
        RECT 140.005 186.515 140.295 187.680 ;
        RECT 143.870 186.950 144.220 188.200 ;
        RECT 145.985 187.775 147.195 188.295 ;
        RECT 147.365 187.605 148.575 188.125 ;
        RECT 140.465 186.515 145.810 186.950 ;
        RECT 145.985 186.515 148.575 187.605 ;
        RECT 149.205 187.605 149.725 188.145 ;
        RECT 149.895 187.775 150.415 188.315 ;
        RECT 149.205 186.515 150.415 187.605 ;
        RECT 11.120 186.345 150.500 186.515 ;
        RECT 11.205 185.255 12.415 186.345 ;
        RECT 12.585 185.255 16.095 186.345 ;
        RECT 11.205 184.545 11.725 185.085 ;
        RECT 11.895 184.715 12.415 185.255 ;
        RECT 12.585 184.565 14.235 185.085 ;
        RECT 14.405 184.735 16.095 185.255 ;
        RECT 17.370 185.375 17.760 185.550 ;
        RECT 18.245 185.545 18.575 186.345 ;
        RECT 18.745 185.555 19.280 186.175 ;
        RECT 17.370 185.205 18.795 185.375 ;
        RECT 11.205 183.795 12.415 184.545 ;
        RECT 12.585 183.795 16.095 184.565 ;
        RECT 17.245 184.475 17.600 185.035 ;
        RECT 17.770 184.305 17.940 185.205 ;
        RECT 18.110 184.475 18.375 185.035 ;
        RECT 18.625 184.705 18.795 185.205 ;
        RECT 18.965 184.535 19.280 185.555 ;
        RECT 19.485 185.205 19.745 186.345 ;
        RECT 19.915 185.195 20.245 186.175 ;
        RECT 20.415 185.205 20.695 186.345 ;
        RECT 20.865 185.255 23.455 186.345 ;
        RECT 19.505 184.785 19.840 185.035 ;
        RECT 20.010 184.595 20.180 185.195 ;
        RECT 20.350 184.765 20.685 185.035 ;
        RECT 17.350 183.795 17.590 184.305 ;
        RECT 17.770 183.975 18.050 184.305 ;
        RECT 18.280 183.795 18.495 184.305 ;
        RECT 18.665 183.965 19.280 184.535 ;
        RECT 19.485 183.965 20.180 184.595 ;
        RECT 20.385 183.795 20.695 184.595 ;
        RECT 20.865 184.565 22.075 185.085 ;
        RECT 22.245 184.735 23.455 185.255 ;
        RECT 24.085 185.180 24.375 186.345 ;
        RECT 20.865 183.795 23.455 184.565 ;
        RECT 24.085 183.795 24.375 184.520 ;
        RECT 24.555 183.975 24.815 186.165 ;
        RECT 24.985 185.615 25.325 186.345 ;
        RECT 25.505 185.435 25.775 186.165 ;
        RECT 25.005 185.215 25.775 185.435 ;
        RECT 25.955 185.455 26.185 186.165 ;
        RECT 26.355 185.635 26.685 186.345 ;
        RECT 26.855 185.455 27.115 186.165 ;
        RECT 25.955 185.215 27.115 185.455 ;
        RECT 27.315 185.375 27.645 186.175 ;
        RECT 27.815 185.545 28.045 186.345 ;
        RECT 28.215 185.375 28.545 186.175 ;
        RECT 25.005 184.545 25.295 185.215 ;
        RECT 27.315 185.205 28.545 185.375 ;
        RECT 28.715 185.205 28.970 186.345 ;
        RECT 30.250 185.375 30.640 185.550 ;
        RECT 31.125 185.545 31.455 186.345 ;
        RECT 31.625 185.555 32.160 186.175 ;
        RECT 30.250 185.205 31.675 185.375 ;
        RECT 25.475 184.725 25.940 185.035 ;
        RECT 26.120 184.725 26.645 185.035 ;
        RECT 25.005 184.345 26.235 184.545 ;
        RECT 25.075 183.795 25.745 184.165 ;
        RECT 25.925 183.975 26.235 184.345 ;
        RECT 26.415 184.085 26.645 184.725 ;
        RECT 26.825 184.705 27.125 185.035 ;
        RECT 27.305 184.705 27.615 185.035 ;
        RECT 26.825 183.795 27.115 184.525 ;
        RECT 27.315 184.305 27.645 184.535 ;
        RECT 27.820 184.475 28.195 185.035 ;
        RECT 28.365 184.305 28.545 185.205 ;
        RECT 28.730 184.455 28.950 185.035 ;
        RECT 30.125 184.475 30.480 185.035 ;
        RECT 30.650 184.305 30.820 185.205 ;
        RECT 30.990 184.475 31.255 185.035 ;
        RECT 31.505 184.705 31.675 185.205 ;
        RECT 31.845 184.535 32.160 185.555 ;
        RECT 32.370 185.955 32.705 186.175 ;
        RECT 33.710 185.965 34.065 186.345 ;
        RECT 32.370 185.335 32.625 185.955 ;
        RECT 32.875 185.795 33.105 185.835 ;
        RECT 34.235 185.795 34.485 186.175 ;
        RECT 32.875 185.595 34.485 185.795 ;
        RECT 32.875 185.505 33.060 185.595 ;
        RECT 33.650 185.585 34.485 185.595 ;
        RECT 34.735 185.565 34.985 186.345 ;
        RECT 35.155 185.495 35.415 186.175 ;
        RECT 33.215 185.395 33.545 185.425 ;
        RECT 33.215 185.335 35.015 185.395 ;
        RECT 32.370 185.225 35.075 185.335 ;
        RECT 32.370 185.165 33.545 185.225 ;
        RECT 34.875 185.190 35.075 185.225 ;
        RECT 32.365 184.785 32.855 184.985 ;
        RECT 33.045 184.785 33.520 184.995 ;
        RECT 27.315 183.965 28.545 184.305 ;
        RECT 28.715 183.795 28.970 184.285 ;
        RECT 30.230 183.795 30.470 184.305 ;
        RECT 30.650 183.975 30.930 184.305 ;
        RECT 31.160 183.795 31.375 184.305 ;
        RECT 31.545 183.965 32.160 184.535 ;
        RECT 32.370 183.795 32.825 184.560 ;
        RECT 33.300 184.385 33.520 184.785 ;
        RECT 33.765 184.785 34.095 184.995 ;
        RECT 33.765 184.385 33.975 184.785 ;
        RECT 34.265 184.750 34.675 185.055 ;
        RECT 34.905 184.615 35.075 185.190 ;
        RECT 34.805 184.495 35.075 184.615 ;
        RECT 34.230 184.450 35.075 184.495 ;
        RECT 34.230 184.325 34.985 184.450 ;
        RECT 34.230 184.175 34.400 184.325 ;
        RECT 35.245 184.295 35.415 185.495 ;
        RECT 35.585 185.205 35.865 186.345 ;
        RECT 36.035 185.195 36.365 186.175 ;
        RECT 36.535 185.205 36.795 186.345 ;
        RECT 37.425 185.205 37.685 186.345 ;
        RECT 37.855 185.375 38.185 186.175 ;
        RECT 38.355 185.545 38.525 186.345 ;
        RECT 38.725 185.375 39.055 186.175 ;
        RECT 39.255 185.545 39.535 186.345 ;
        RECT 40.190 185.835 41.845 186.125 ;
        RECT 40.190 185.495 41.780 185.665 ;
        RECT 42.015 185.545 42.295 186.345 ;
        RECT 37.855 185.205 39.135 185.375 ;
        RECT 36.100 185.155 36.275 185.195 ;
        RECT 35.595 184.765 35.930 185.035 ;
        RECT 36.100 184.595 36.270 185.155 ;
        RECT 36.440 184.785 36.775 185.035 ;
        RECT 37.450 184.705 37.735 185.035 ;
        RECT 37.935 184.705 38.315 185.035 ;
        RECT 38.485 184.705 38.795 185.035 ;
        RECT 33.100 183.965 34.400 184.175 ;
        RECT 34.655 183.795 34.985 184.155 ;
        RECT 35.155 183.965 35.415 184.295 ;
        RECT 35.585 183.795 35.895 184.595 ;
        RECT 36.100 183.965 36.795 184.595 ;
        RECT 37.430 183.795 37.765 184.535 ;
        RECT 37.935 184.010 38.150 184.705 ;
        RECT 38.485 184.535 38.690 184.705 ;
        RECT 38.965 184.535 39.135 185.205 ;
        RECT 39.315 184.705 39.555 185.375 ;
        RECT 40.190 185.205 40.510 185.495 ;
        RECT 41.610 185.375 41.780 185.495 ;
        RECT 40.705 185.155 41.420 185.325 ;
        RECT 41.610 185.205 42.335 185.375 ;
        RECT 42.505 185.205 42.775 186.175 ;
        RECT 42.945 185.255 45.535 186.345 ;
        RECT 46.165 185.545 46.425 186.345 ;
        RECT 38.340 184.010 38.690 184.535 ;
        RECT 38.860 183.965 39.555 184.535 ;
        RECT 40.190 184.465 40.540 185.035 ;
        RECT 40.710 184.705 41.420 185.155 ;
        RECT 42.165 185.035 42.335 185.205 ;
        RECT 41.590 184.705 41.995 185.035 ;
        RECT 42.165 184.705 42.435 185.035 ;
        RECT 42.165 184.535 42.335 184.705 ;
        RECT 40.725 184.365 42.335 184.535 ;
        RECT 42.605 184.470 42.775 185.205 ;
        RECT 40.195 183.795 40.525 184.295 ;
        RECT 40.725 184.015 40.895 184.365 ;
        RECT 41.095 183.795 41.425 184.195 ;
        RECT 41.595 184.015 41.765 184.365 ;
        RECT 41.935 183.795 42.315 184.195 ;
        RECT 42.505 184.125 42.775 184.470 ;
        RECT 42.945 184.565 44.155 185.085 ;
        RECT 44.325 184.735 45.535 185.255 ;
        RECT 42.945 183.795 45.535 184.565 ;
        RECT 46.165 184.365 46.425 185.375 ;
        RECT 46.685 184.955 46.925 186.160 ;
        RECT 47.095 185.325 47.350 186.160 ;
        RECT 47.955 185.375 48.290 186.160 ;
        RECT 47.095 185.125 47.535 185.325 ;
        RECT 46.685 184.785 47.135 184.955 ;
        RECT 47.305 184.705 47.535 185.125 ;
        RECT 47.705 185.205 48.290 185.375 ;
        RECT 48.465 185.255 49.675 186.345 ;
        RECT 47.705 184.535 47.875 185.205 ;
        RECT 46.675 184.365 47.875 184.535 ;
        RECT 48.045 184.455 48.295 185.035 ;
        RECT 48.465 184.545 48.985 185.085 ;
        RECT 49.155 184.715 49.675 185.255 ;
        RECT 49.845 185.180 50.135 186.345 ;
        RECT 50.605 185.705 50.935 186.135 ;
        RECT 50.480 185.535 50.935 185.705 ;
        RECT 51.115 185.705 51.365 186.125 ;
        RECT 51.595 185.875 51.925 186.345 ;
        RECT 52.155 185.705 52.405 186.125 ;
        RECT 51.115 185.535 52.405 185.705 ;
        RECT 46.175 183.795 46.505 184.195 ;
        RECT 46.675 184.095 46.845 184.365 ;
        RECT 47.520 184.355 47.875 184.365 ;
        RECT 47.015 183.795 47.345 184.195 ;
        RECT 47.520 184.095 47.785 184.355 ;
        RECT 48.035 183.795 48.295 184.285 ;
        RECT 48.465 183.795 49.675 184.545 ;
        RECT 50.480 184.535 50.650 185.535 ;
        RECT 50.820 184.705 51.065 185.365 ;
        RECT 51.280 184.705 51.545 185.365 ;
        RECT 51.740 184.705 52.025 185.365 ;
        RECT 52.200 185.035 52.415 185.365 ;
        RECT 52.595 185.205 52.845 186.345 ;
        RECT 53.015 185.285 53.345 186.135 ;
        RECT 53.525 185.910 58.870 186.345 ;
        RECT 52.200 184.705 52.505 185.035 ;
        RECT 52.675 184.705 52.985 185.035 ;
        RECT 52.675 184.535 52.845 184.705 ;
        RECT 49.845 183.795 50.135 184.520 ;
        RECT 50.480 184.365 52.845 184.535 ;
        RECT 53.155 184.520 53.345 185.285 ;
        RECT 50.635 183.795 50.965 184.195 ;
        RECT 51.135 184.025 51.465 184.365 ;
        RECT 52.515 183.795 52.845 184.195 ;
        RECT 53.015 184.010 53.345 184.520 ;
        RECT 55.110 184.340 55.450 185.170 ;
        RECT 56.930 184.660 57.280 185.910 ;
        RECT 59.045 185.255 62.555 186.345 ;
        RECT 59.045 184.565 60.695 185.085 ;
        RECT 60.865 184.735 62.555 185.255 ;
        RECT 63.190 185.205 63.445 186.345 ;
        RECT 63.615 185.375 63.945 186.175 ;
        RECT 64.115 185.545 64.345 186.345 ;
        RECT 64.515 185.375 64.845 186.175 ;
        RECT 63.615 185.205 64.845 185.375 ;
        RECT 65.025 185.255 66.695 186.345 ;
        RECT 53.525 183.795 58.870 184.340 ;
        RECT 59.045 183.795 62.555 184.565 ;
        RECT 63.210 184.455 63.430 185.035 ;
        RECT 63.615 184.305 63.795 185.205 ;
        RECT 63.965 184.475 64.340 185.035 ;
        RECT 64.545 184.705 64.855 185.035 ;
        RECT 65.025 184.565 65.775 185.085 ;
        RECT 65.945 184.735 66.695 185.255 ;
        RECT 67.510 185.375 67.900 185.550 ;
        RECT 68.385 185.545 68.715 186.345 ;
        RECT 68.885 185.555 69.420 186.175 ;
        RECT 67.510 185.205 68.935 185.375 ;
        RECT 64.515 184.305 64.845 184.535 ;
        RECT 63.190 183.795 63.445 184.285 ;
        RECT 63.615 183.965 64.845 184.305 ;
        RECT 65.025 183.795 66.695 184.565 ;
        RECT 67.385 184.475 67.740 185.035 ;
        RECT 67.910 184.305 68.080 185.205 ;
        RECT 68.250 184.475 68.515 185.035 ;
        RECT 68.765 184.705 68.935 185.205 ;
        RECT 69.105 184.535 69.420 185.555 ;
        RECT 69.625 185.255 70.835 186.345 ;
        RECT 67.490 183.795 67.730 184.305 ;
        RECT 67.910 183.975 68.190 184.305 ;
        RECT 68.420 183.795 68.635 184.305 ;
        RECT 68.805 183.965 69.420 184.535 ;
        RECT 69.625 184.545 70.145 185.085 ;
        RECT 70.315 184.715 70.835 185.255 ;
        RECT 71.010 185.205 71.285 186.175 ;
        RECT 71.495 185.545 71.775 186.345 ;
        RECT 71.945 185.835 73.135 186.125 ;
        RECT 71.945 185.495 73.115 185.665 ;
        RECT 71.945 185.375 72.115 185.495 ;
        RECT 71.455 185.205 72.115 185.375 ;
        RECT 69.625 183.795 70.835 184.545 ;
        RECT 71.010 184.470 71.180 185.205 ;
        RECT 71.455 185.035 71.625 185.205 ;
        RECT 72.425 185.035 72.620 185.325 ;
        RECT 72.790 185.205 73.115 185.495 ;
        RECT 73.305 185.255 74.975 186.345 ;
        RECT 71.350 184.705 71.625 185.035 ;
        RECT 71.795 184.705 72.620 185.035 ;
        RECT 72.790 184.705 73.135 185.035 ;
        RECT 71.455 184.535 71.625 184.705 ;
        RECT 73.305 184.565 74.055 185.085 ;
        RECT 74.225 184.735 74.975 185.255 ;
        RECT 75.605 185.180 75.895 186.345 ;
        RECT 76.990 185.545 77.305 186.345 ;
        RECT 77.570 186.005 78.650 186.160 ;
        RECT 77.505 185.990 78.650 186.005 ;
        RECT 77.505 185.835 77.740 185.990 ;
        RECT 77.570 185.375 77.740 185.835 ;
        RECT 71.010 184.125 71.285 184.470 ;
        RECT 71.455 184.365 73.120 184.535 ;
        RECT 71.475 183.795 71.855 184.195 ;
        RECT 72.025 184.015 72.195 184.365 ;
        RECT 72.365 183.795 72.695 184.195 ;
        RECT 72.865 184.015 73.120 184.365 ;
        RECT 73.305 183.795 74.975 184.565 ;
        RECT 75.605 183.795 75.895 184.520 ;
        RECT 76.985 184.365 77.255 185.375 ;
        RECT 77.425 185.205 77.740 185.375 ;
        RECT 77.425 184.535 77.595 185.205 ;
        RECT 77.910 185.035 78.145 185.715 ;
        RECT 78.315 185.205 78.650 185.990 ;
        RECT 78.915 185.415 79.085 186.175 ;
        RECT 79.300 185.585 79.630 186.345 ;
        RECT 78.915 185.245 79.630 185.415 ;
        RECT 79.800 185.270 80.055 186.175 ;
        RECT 77.765 184.705 78.145 185.035 ;
        RECT 78.315 184.705 78.650 185.035 ;
        RECT 78.825 184.695 79.180 185.065 ;
        RECT 79.460 185.035 79.630 185.245 ;
        RECT 79.460 184.705 79.715 185.035 ;
        RECT 77.425 184.365 78.650 184.535 ;
        RECT 79.460 184.515 79.630 184.705 ;
        RECT 79.885 184.540 80.055 185.270 ;
        RECT 80.230 185.195 80.490 186.345 ;
        RECT 80.665 185.255 84.175 186.345 ;
        RECT 77.055 183.795 77.385 184.195 ;
        RECT 77.555 184.095 77.725 184.365 ;
        RECT 77.895 183.795 78.225 184.195 ;
        RECT 78.395 184.095 78.650 184.365 ;
        RECT 78.915 184.345 79.630 184.515 ;
        RECT 78.915 183.965 79.085 184.345 ;
        RECT 79.300 183.795 79.630 184.175 ;
        RECT 79.800 183.965 80.055 184.540 ;
        RECT 80.230 183.795 80.490 184.635 ;
        RECT 80.665 184.565 82.315 185.085 ;
        RECT 82.485 184.735 84.175 185.255 ;
        RECT 84.805 185.495 85.185 186.175 ;
        RECT 85.775 185.495 85.945 186.345 ;
        RECT 86.115 185.665 86.445 186.175 ;
        RECT 86.615 185.835 86.785 186.345 ;
        RECT 86.955 185.665 87.355 186.175 ;
        RECT 86.115 185.495 87.355 185.665 ;
        RECT 80.665 183.795 84.175 184.565 ;
        RECT 84.805 184.535 84.975 185.495 ;
        RECT 85.145 185.155 86.450 185.325 ;
        RECT 87.535 185.245 87.855 186.175 ;
        RECT 88.025 185.255 89.235 186.345 ;
        RECT 85.145 184.705 85.390 185.155 ;
        RECT 85.560 184.785 86.110 184.985 ;
        RECT 86.280 184.955 86.450 185.155 ;
        RECT 87.225 185.075 87.855 185.245 ;
        RECT 86.280 184.785 86.655 184.955 ;
        RECT 86.825 184.535 87.055 185.035 ;
        RECT 84.805 184.365 87.055 184.535 ;
        RECT 84.855 183.795 85.185 184.185 ;
        RECT 85.355 184.045 85.525 184.365 ;
        RECT 87.225 184.195 87.395 185.075 ;
        RECT 85.695 183.795 86.025 184.185 ;
        RECT 86.440 184.025 87.395 184.195 ;
        RECT 87.565 183.795 87.855 184.630 ;
        RECT 88.025 184.545 88.545 185.085 ;
        RECT 88.715 184.715 89.235 185.255 ;
        RECT 89.405 185.475 89.680 186.175 ;
        RECT 89.850 185.800 90.105 186.345 ;
        RECT 90.275 185.835 90.755 186.175 ;
        RECT 90.930 185.790 91.535 186.345 ;
        RECT 91.705 185.910 97.050 186.345 ;
        RECT 90.920 185.690 91.535 185.790 ;
        RECT 90.920 185.665 91.105 185.690 ;
        RECT 88.025 183.795 89.235 184.545 ;
        RECT 89.405 184.445 89.575 185.475 ;
        RECT 89.850 185.345 90.605 185.595 ;
        RECT 90.775 185.420 91.105 185.665 ;
        RECT 89.850 185.310 90.620 185.345 ;
        RECT 89.850 185.300 90.635 185.310 ;
        RECT 89.745 185.285 90.640 185.300 ;
        RECT 89.745 185.270 90.660 185.285 ;
        RECT 89.745 185.260 90.680 185.270 ;
        RECT 89.745 185.250 90.705 185.260 ;
        RECT 89.745 185.220 90.775 185.250 ;
        RECT 89.745 185.190 90.795 185.220 ;
        RECT 89.745 185.160 90.815 185.190 ;
        RECT 89.745 185.135 90.845 185.160 ;
        RECT 89.745 185.100 90.880 185.135 ;
        RECT 89.745 185.095 90.910 185.100 ;
        RECT 89.745 184.700 89.975 185.095 ;
        RECT 90.520 185.090 90.910 185.095 ;
        RECT 90.545 185.080 90.910 185.090 ;
        RECT 90.560 185.075 90.910 185.080 ;
        RECT 90.575 185.070 90.910 185.075 ;
        RECT 91.275 185.070 91.535 185.520 ;
        RECT 90.575 185.065 91.535 185.070 ;
        RECT 90.585 185.055 91.535 185.065 ;
        RECT 90.595 185.050 91.535 185.055 ;
        RECT 90.605 185.040 91.535 185.050 ;
        RECT 90.610 185.030 91.535 185.040 ;
        RECT 90.615 185.025 91.535 185.030 ;
        RECT 90.625 185.010 91.535 185.025 ;
        RECT 90.630 184.995 91.535 185.010 ;
        RECT 90.640 184.970 91.535 184.995 ;
        RECT 90.145 184.500 90.475 184.925 ;
        RECT 89.405 183.965 89.665 184.445 ;
        RECT 89.835 183.795 90.085 184.335 ;
        RECT 90.255 184.015 90.475 184.500 ;
        RECT 90.645 184.900 91.535 184.970 ;
        RECT 90.645 184.175 90.815 184.900 ;
        RECT 90.985 184.345 91.535 184.730 ;
        RECT 93.290 184.340 93.630 185.170 ;
        RECT 95.110 184.660 95.460 185.910 ;
        RECT 97.225 185.255 100.735 186.345 ;
        RECT 97.225 184.565 98.875 185.085 ;
        RECT 99.045 184.735 100.735 185.255 ;
        RECT 101.365 185.180 101.655 186.345 ;
        RECT 101.825 185.245 102.145 186.175 ;
        RECT 102.325 185.665 102.725 186.175 ;
        RECT 102.895 185.835 103.065 186.345 ;
        RECT 103.235 185.665 103.565 186.175 ;
        RECT 102.325 185.495 103.565 185.665 ;
        RECT 103.735 185.495 103.905 186.345 ;
        RECT 104.495 185.495 104.875 186.175 ;
        RECT 101.825 185.075 102.455 185.245 ;
        RECT 90.645 184.005 91.535 184.175 ;
        RECT 91.705 183.795 97.050 184.340 ;
        RECT 97.225 183.795 100.735 184.565 ;
        RECT 101.365 183.795 101.655 184.520 ;
        RECT 101.825 183.795 102.115 184.630 ;
        RECT 102.285 184.195 102.455 185.075 ;
        RECT 103.230 185.155 104.535 185.325 ;
        RECT 102.625 184.535 102.855 185.035 ;
        RECT 103.230 184.955 103.400 185.155 ;
        RECT 103.025 184.785 103.400 184.955 ;
        RECT 103.570 184.785 104.120 184.985 ;
        RECT 104.290 184.705 104.535 185.155 ;
        RECT 104.705 184.535 104.875 185.495 ;
        RECT 105.045 185.255 107.635 186.345 ;
        RECT 102.625 184.365 104.875 184.535 ;
        RECT 105.045 184.565 106.255 185.085 ;
        RECT 106.425 184.735 107.635 185.255 ;
        RECT 107.925 185.225 108.255 186.345 ;
        RECT 107.865 184.785 108.375 185.035 ;
        RECT 108.585 184.785 108.955 186.100 ;
        RECT 109.125 184.785 109.455 186.100 ;
        RECT 109.665 184.785 109.995 186.100 ;
        RECT 110.265 185.455 110.515 186.175 ;
        RECT 110.685 185.625 111.015 186.345 ;
        RECT 110.265 185.165 111.015 185.455 ;
        RECT 111.250 185.165 111.775 186.175 ;
        RECT 112.005 185.645 112.225 186.175 ;
        RECT 112.395 185.835 112.725 186.345 ;
        RECT 112.895 185.645 113.120 186.175 ;
        RECT 112.005 185.380 113.120 185.645 ;
        RECT 113.290 185.630 113.605 186.175 ;
        RECT 113.795 185.930 114.125 186.345 ;
        RECT 113.290 185.400 114.125 185.630 ;
        RECT 110.755 184.995 111.015 185.165 ;
        RECT 110.165 184.785 110.585 184.995 ;
        RECT 110.755 184.785 111.335 184.995 ;
        RECT 110.755 184.615 111.125 184.785 ;
        RECT 102.285 184.025 103.240 184.195 ;
        RECT 103.655 183.795 103.985 184.185 ;
        RECT 104.155 184.045 104.325 184.365 ;
        RECT 104.495 183.795 104.825 184.185 ;
        RECT 105.045 183.795 107.635 184.565 ;
        RECT 107.905 184.445 110.205 184.615 ;
        RECT 107.905 183.965 108.235 184.445 ;
        RECT 108.405 183.795 108.735 184.255 ;
        RECT 108.950 183.965 109.280 184.445 ;
        RECT 109.480 183.795 109.810 184.255 ;
        RECT 110.035 184.125 110.205 184.445 ;
        RECT 110.375 184.425 111.125 184.615 ;
        RECT 111.505 184.595 111.775 185.165 ;
        RECT 110.375 183.980 110.705 184.425 ;
        RECT 110.975 183.795 111.145 184.255 ;
        RECT 111.435 183.965 111.775 184.595 ;
        RECT 111.955 184.460 112.270 185.035 ;
        RECT 111.945 183.795 112.275 184.275 ;
        RECT 112.460 184.075 112.840 185.035 ;
        RECT 113.290 184.705 113.615 185.120 ;
        RECT 113.785 184.705 114.125 185.400 ;
        RECT 113.785 184.535 113.955 184.705 ;
        RECT 114.295 184.535 114.525 186.175 ;
        RECT 114.695 185.375 114.985 186.345 ;
        RECT 115.175 185.205 115.505 186.345 ;
        RECT 116.035 185.375 116.365 186.160 ;
        RECT 115.685 185.205 116.365 185.375 ;
        RECT 116.545 185.255 118.215 186.345 ;
        RECT 115.165 184.785 115.515 185.035 ;
        RECT 115.685 184.605 115.855 185.205 ;
        RECT 116.025 184.785 116.375 185.035 ;
        RECT 113.215 184.365 113.955 184.535 ;
        RECT 113.215 183.965 113.405 184.365 ;
        RECT 114.125 184.345 114.525 184.535 ;
        RECT 113.625 183.795 113.955 184.155 ;
        RECT 114.125 183.965 114.315 184.345 ;
        RECT 114.485 183.795 114.815 184.175 ;
        RECT 115.175 183.795 115.445 184.605 ;
        RECT 115.615 183.965 115.945 184.605 ;
        RECT 116.115 183.795 116.355 184.605 ;
        RECT 116.545 184.565 117.295 185.085 ;
        RECT 117.465 184.735 118.215 185.255 ;
        RECT 118.855 185.285 119.185 186.135 ;
        RECT 116.545 183.795 118.215 184.565 ;
        RECT 118.855 184.520 119.045 185.285 ;
        RECT 119.355 185.205 119.605 186.345 ;
        RECT 119.795 185.705 120.045 186.125 ;
        RECT 120.275 185.875 120.605 186.345 ;
        RECT 120.835 185.705 121.085 186.125 ;
        RECT 119.795 185.535 121.085 185.705 ;
        RECT 121.265 185.705 121.595 186.135 ;
        RECT 121.265 185.535 121.720 185.705 ;
        RECT 119.785 185.035 120.000 185.365 ;
        RECT 119.215 184.705 119.525 185.035 ;
        RECT 119.695 184.705 120.000 185.035 ;
        RECT 120.175 184.705 120.460 185.365 ;
        RECT 120.655 184.705 120.920 185.365 ;
        RECT 121.135 184.705 121.380 185.365 ;
        RECT 119.355 184.535 119.525 184.705 ;
        RECT 121.550 184.535 121.720 185.535 ;
        RECT 122.065 185.255 124.655 186.345 ;
        RECT 125.025 185.675 125.305 186.345 ;
        RECT 125.475 185.455 125.775 186.005 ;
        RECT 125.975 185.625 126.305 186.345 ;
        RECT 126.495 185.625 126.955 186.175 ;
        RECT 118.855 184.010 119.185 184.520 ;
        RECT 119.355 184.365 121.720 184.535 ;
        RECT 122.065 184.565 123.275 185.085 ;
        RECT 123.445 184.735 124.655 185.255 ;
        RECT 124.840 185.035 125.105 185.395 ;
        RECT 125.475 185.285 126.415 185.455 ;
        RECT 126.245 185.035 126.415 185.285 ;
        RECT 124.840 184.785 125.515 185.035 ;
        RECT 125.735 184.785 126.075 185.035 ;
        RECT 126.245 184.705 126.535 185.035 ;
        RECT 126.245 184.615 126.415 184.705 ;
        RECT 119.355 183.795 119.685 184.195 ;
        RECT 120.735 184.025 121.065 184.365 ;
        RECT 121.235 183.795 121.565 184.195 ;
        RECT 122.065 183.795 124.655 184.565 ;
        RECT 125.025 184.425 126.415 184.615 ;
        RECT 125.025 184.065 125.355 184.425 ;
        RECT 126.705 184.255 126.955 185.625 ;
        RECT 127.125 185.180 127.415 186.345 ;
        RECT 127.675 185.675 127.845 186.175 ;
        RECT 128.015 185.845 128.345 186.345 ;
        RECT 127.675 185.505 128.340 185.675 ;
        RECT 127.590 184.685 127.940 185.335 ;
        RECT 125.975 183.795 126.225 184.255 ;
        RECT 126.395 183.965 126.955 184.255 ;
        RECT 127.125 183.795 127.415 184.520 ;
        RECT 128.110 184.515 128.340 185.505 ;
        RECT 127.675 184.345 128.340 184.515 ;
        RECT 127.675 184.055 127.845 184.345 ;
        RECT 128.015 183.795 128.345 184.175 ;
        RECT 128.515 184.055 128.700 186.175 ;
        RECT 128.940 185.885 129.205 186.345 ;
        RECT 129.375 185.750 129.625 186.175 ;
        RECT 129.835 185.900 130.940 186.070 ;
        RECT 129.320 185.620 129.625 185.750 ;
        RECT 128.870 184.425 129.150 185.375 ;
        RECT 129.320 184.515 129.490 185.620 ;
        RECT 129.660 184.835 129.900 185.430 ;
        RECT 130.070 185.365 130.600 185.730 ;
        RECT 130.070 184.665 130.240 185.365 ;
        RECT 130.770 185.285 130.940 185.900 ;
        RECT 131.110 185.545 131.280 186.345 ;
        RECT 131.450 185.845 131.700 186.175 ;
        RECT 131.925 185.875 132.810 186.045 ;
        RECT 130.770 185.195 131.280 185.285 ;
        RECT 129.320 184.385 129.545 184.515 ;
        RECT 129.715 184.445 130.240 184.665 ;
        RECT 130.410 185.025 131.280 185.195 ;
        RECT 128.955 183.795 129.205 184.255 ;
        RECT 129.375 184.245 129.545 184.385 ;
        RECT 130.410 184.245 130.580 185.025 ;
        RECT 131.110 184.955 131.280 185.025 ;
        RECT 130.790 184.775 130.990 184.805 ;
        RECT 131.450 184.775 131.620 185.845 ;
        RECT 131.790 184.955 131.980 185.675 ;
        RECT 130.790 184.475 131.620 184.775 ;
        RECT 132.150 184.745 132.470 185.705 ;
        RECT 129.375 184.075 129.710 184.245 ;
        RECT 129.905 184.075 130.580 184.245 ;
        RECT 130.900 183.795 131.270 184.295 ;
        RECT 131.450 184.245 131.620 184.475 ;
        RECT 132.005 184.415 132.470 184.745 ;
        RECT 132.640 185.035 132.810 185.875 ;
        RECT 132.990 185.845 133.305 186.345 ;
        RECT 133.535 185.615 133.875 186.175 ;
        RECT 132.980 185.240 133.875 185.615 ;
        RECT 134.045 185.335 134.215 186.345 ;
        RECT 133.685 185.035 133.875 185.240 ;
        RECT 134.385 185.285 134.715 186.130 ;
        RECT 134.885 185.430 135.055 186.345 ;
        RECT 135.405 185.910 140.750 186.345 ;
        RECT 140.925 185.910 146.270 186.345 ;
        RECT 134.385 185.205 134.775 185.285 ;
        RECT 134.560 185.155 134.775 185.205 ;
        RECT 132.640 184.705 133.515 185.035 ;
        RECT 133.685 184.705 134.435 185.035 ;
        RECT 132.640 184.245 132.810 184.705 ;
        RECT 133.685 184.535 133.885 184.705 ;
        RECT 134.605 184.575 134.775 185.155 ;
        RECT 134.550 184.535 134.775 184.575 ;
        RECT 131.450 184.075 131.855 184.245 ;
        RECT 132.025 184.075 132.810 184.245 ;
        RECT 133.085 183.795 133.295 184.325 ;
        RECT 133.555 184.010 133.885 184.535 ;
        RECT 134.395 184.450 134.775 184.535 ;
        RECT 134.055 183.795 134.225 184.405 ;
        RECT 134.395 184.015 134.725 184.450 ;
        RECT 136.990 184.340 137.330 185.170 ;
        RECT 138.810 184.660 139.160 185.910 ;
        RECT 142.510 184.340 142.850 185.170 ;
        RECT 144.330 184.660 144.680 185.910 ;
        RECT 146.445 185.255 149.035 186.345 ;
        RECT 146.445 184.565 147.655 185.085 ;
        RECT 147.825 184.735 149.035 185.255 ;
        RECT 149.205 185.255 150.415 186.345 ;
        RECT 149.205 184.715 149.725 185.255 ;
        RECT 134.895 183.795 135.065 184.310 ;
        RECT 135.405 183.795 140.750 184.340 ;
        RECT 140.925 183.795 146.270 184.340 ;
        RECT 146.445 183.795 149.035 184.565 ;
        RECT 149.895 184.545 150.415 185.085 ;
        RECT 149.205 183.795 150.415 184.545 ;
        RECT 11.120 183.625 150.500 183.795 ;
        RECT 11.205 182.875 12.415 183.625 ;
        RECT 11.205 182.335 11.725 182.875 ;
        RECT 12.585 182.855 15.175 183.625 ;
        RECT 15.815 182.895 16.115 183.625 ;
        RECT 11.895 182.165 12.415 182.705 ;
        RECT 12.585 182.335 13.795 182.855 ;
        RECT 16.295 182.715 16.525 183.335 ;
        RECT 16.725 183.065 16.950 183.445 ;
        RECT 17.120 183.235 17.450 183.625 ;
        RECT 16.725 182.885 17.055 183.065 ;
        RECT 13.965 182.165 15.175 182.685 ;
        RECT 15.820 182.385 16.115 182.715 ;
        RECT 16.295 182.385 16.710 182.715 ;
        RECT 16.880 182.215 17.055 182.885 ;
        RECT 17.225 182.385 17.465 183.035 ;
        RECT 18.565 182.885 18.950 183.455 ;
        RECT 19.120 183.165 19.445 183.625 ;
        RECT 19.965 182.995 20.245 183.455 ;
        RECT 18.565 182.215 18.845 182.885 ;
        RECT 19.120 182.825 20.245 182.995 ;
        RECT 19.120 182.715 19.570 182.825 ;
        RECT 19.015 182.385 19.570 182.715 ;
        RECT 20.435 182.655 20.835 183.455 ;
        RECT 21.235 183.165 21.505 183.625 ;
        RECT 21.675 182.995 21.960 183.455 ;
        RECT 22.245 183.080 27.590 183.625 ;
        RECT 11.205 181.075 12.415 182.165 ;
        RECT 12.585 181.075 15.175 182.165 ;
        RECT 15.815 181.855 16.710 182.185 ;
        RECT 16.880 182.025 17.465 182.215 ;
        RECT 15.815 181.685 17.020 181.855 ;
        RECT 15.815 181.255 16.145 181.685 ;
        RECT 16.325 181.075 16.520 181.515 ;
        RECT 16.690 181.255 17.020 181.685 ;
        RECT 17.190 181.255 17.465 182.025 ;
        RECT 18.565 181.245 18.950 182.215 ;
        RECT 19.120 181.925 19.570 182.385 ;
        RECT 19.740 182.095 20.835 182.655 ;
        RECT 19.120 181.705 20.245 181.925 ;
        RECT 19.120 181.075 19.445 181.535 ;
        RECT 19.965 181.245 20.245 181.705 ;
        RECT 20.435 181.245 20.835 182.095 ;
        RECT 21.005 182.825 21.960 182.995 ;
        RECT 21.005 181.925 21.215 182.825 ;
        RECT 21.385 182.095 22.075 182.655 ;
        RECT 23.830 182.250 24.170 183.080 ;
        RECT 27.765 182.855 30.355 183.625 ;
        RECT 30.690 183.115 30.930 183.625 ;
        RECT 31.110 183.115 31.390 183.445 ;
        RECT 31.620 183.115 31.835 183.625 ;
        RECT 21.005 181.705 21.960 181.925 ;
        RECT 21.235 181.075 21.505 181.535 ;
        RECT 21.675 181.245 21.960 181.705 ;
        RECT 25.650 181.510 26.000 182.760 ;
        RECT 27.765 182.335 28.975 182.855 ;
        RECT 29.145 182.165 30.355 182.685 ;
        RECT 30.585 182.385 30.940 182.945 ;
        RECT 31.110 182.215 31.280 183.115 ;
        RECT 31.450 182.385 31.715 182.945 ;
        RECT 32.005 182.885 32.620 183.455 ;
        RECT 31.965 182.215 32.135 182.715 ;
        RECT 22.245 181.075 27.590 181.510 ;
        RECT 27.765 181.075 30.355 182.165 ;
        RECT 30.710 182.045 32.135 182.215 ;
        RECT 30.710 181.870 31.100 182.045 ;
        RECT 31.585 181.075 31.915 181.875 ;
        RECT 32.305 181.865 32.620 182.885 ;
        RECT 32.825 182.855 36.335 183.625 ;
        RECT 36.965 182.900 37.255 183.625 ;
        RECT 37.425 182.855 40.935 183.625 ;
        RECT 41.105 182.875 42.315 183.625 ;
        RECT 32.825 182.335 34.475 182.855 ;
        RECT 34.645 182.165 36.335 182.685 ;
        RECT 37.425 182.335 39.075 182.855 ;
        RECT 32.085 181.245 32.620 181.865 ;
        RECT 32.825 181.075 36.335 182.165 ;
        RECT 36.965 181.075 37.255 182.240 ;
        RECT 39.245 182.165 40.935 182.685 ;
        RECT 41.105 182.335 41.625 182.875 ;
        RECT 42.490 182.785 42.750 183.625 ;
        RECT 42.925 182.880 43.180 183.455 ;
        RECT 43.350 183.245 43.680 183.625 ;
        RECT 43.895 183.075 44.065 183.455 ;
        RECT 44.325 183.080 49.670 183.625 ;
        RECT 43.350 182.905 44.065 183.075 ;
        RECT 41.795 182.165 42.315 182.705 ;
        RECT 37.425 181.075 40.935 182.165 ;
        RECT 41.105 181.075 42.315 182.165 ;
        RECT 42.490 181.075 42.750 182.225 ;
        RECT 42.925 182.150 43.095 182.880 ;
        RECT 43.350 182.715 43.520 182.905 ;
        RECT 43.265 182.385 43.520 182.715 ;
        RECT 43.350 182.175 43.520 182.385 ;
        RECT 43.800 182.355 44.155 182.725 ;
        RECT 45.910 182.250 46.250 183.080 ;
        RECT 49.850 182.950 50.125 183.295 ;
        RECT 50.315 183.225 50.695 183.625 ;
        RECT 50.865 183.055 51.035 183.405 ;
        RECT 51.205 183.225 51.535 183.625 ;
        RECT 51.705 183.055 51.960 183.405 ;
        RECT 42.925 181.245 43.180 182.150 ;
        RECT 43.350 182.005 44.065 182.175 ;
        RECT 43.350 181.075 43.680 181.835 ;
        RECT 43.895 181.245 44.065 182.005 ;
        RECT 47.730 181.510 48.080 182.760 ;
        RECT 49.850 182.215 50.020 182.950 ;
        RECT 50.295 182.885 51.960 183.055 ;
        RECT 50.295 182.715 50.465 182.885 ;
        RECT 52.145 182.855 54.735 183.625 ;
        RECT 54.915 182.895 55.215 183.625 ;
        RECT 50.190 182.385 50.465 182.715 ;
        RECT 50.635 182.385 51.460 182.715 ;
        RECT 51.630 182.385 51.975 182.715 ;
        RECT 50.295 182.215 50.465 182.385 ;
        RECT 44.325 181.075 49.670 181.510 ;
        RECT 49.850 181.245 50.125 182.215 ;
        RECT 50.295 182.045 50.955 182.215 ;
        RECT 51.265 182.095 51.460 182.385 ;
        RECT 52.145 182.335 53.355 182.855 ;
        RECT 55.395 182.715 55.625 183.335 ;
        RECT 55.825 183.065 56.050 183.445 ;
        RECT 56.220 183.235 56.550 183.625 ;
        RECT 55.825 182.885 56.155 183.065 ;
        RECT 50.785 181.925 50.955 182.045 ;
        RECT 51.630 181.925 51.955 182.215 ;
        RECT 53.525 182.165 54.735 182.685 ;
        RECT 54.920 182.385 55.215 182.715 ;
        RECT 55.395 182.385 55.810 182.715 ;
        RECT 55.980 182.215 56.155 182.885 ;
        RECT 56.325 182.385 56.565 183.035 ;
        RECT 56.745 182.855 60.255 183.625 ;
        RECT 60.895 182.895 61.195 183.625 ;
        RECT 56.745 182.335 58.395 182.855 ;
        RECT 61.375 182.715 61.605 183.335 ;
        RECT 61.805 183.065 62.030 183.445 ;
        RECT 62.200 183.235 62.530 183.625 ;
        RECT 61.805 182.885 62.135 183.065 ;
        RECT 50.335 181.075 50.615 181.875 ;
        RECT 50.785 181.755 51.955 181.925 ;
        RECT 50.785 181.295 51.975 181.585 ;
        RECT 52.145 181.075 54.735 182.165 ;
        RECT 54.915 181.855 55.810 182.185 ;
        RECT 55.980 182.025 56.565 182.215 ;
        RECT 58.565 182.165 60.255 182.685 ;
        RECT 60.900 182.385 61.195 182.715 ;
        RECT 61.375 182.385 61.790 182.715 ;
        RECT 61.960 182.215 62.135 182.885 ;
        RECT 62.305 182.385 62.545 183.035 ;
        RECT 62.725 182.900 63.015 183.625 ;
        RECT 63.390 182.845 63.890 183.455 ;
        RECT 63.185 182.385 63.535 182.635 ;
        RECT 54.915 181.685 56.120 181.855 ;
        RECT 54.915 181.255 55.245 181.685 ;
        RECT 55.425 181.075 55.620 181.515 ;
        RECT 55.790 181.255 56.120 181.685 ;
        RECT 56.290 181.255 56.565 182.025 ;
        RECT 56.745 181.075 60.255 182.165 ;
        RECT 60.895 181.855 61.790 182.185 ;
        RECT 61.960 182.025 62.545 182.215 ;
        RECT 60.895 181.685 62.100 181.855 ;
        RECT 60.895 181.255 61.225 181.685 ;
        RECT 61.405 181.075 61.600 181.515 ;
        RECT 61.770 181.255 62.100 181.685 ;
        RECT 62.270 181.255 62.545 182.025 ;
        RECT 62.725 181.075 63.015 182.240 ;
        RECT 63.720 182.215 63.890 182.845 ;
        RECT 64.520 182.975 64.850 183.455 ;
        RECT 65.020 183.165 65.245 183.625 ;
        RECT 65.415 182.975 65.745 183.455 ;
        RECT 64.520 182.805 65.745 182.975 ;
        RECT 65.935 182.825 66.185 183.625 ;
        RECT 66.355 182.825 66.695 183.455 ;
        RECT 66.865 183.080 72.210 183.625 ;
        RECT 64.060 182.435 64.390 182.635 ;
        RECT 64.560 182.435 64.890 182.635 ;
        RECT 65.060 182.435 65.480 182.635 ;
        RECT 65.655 182.465 66.350 182.635 ;
        RECT 65.655 182.215 65.825 182.465 ;
        RECT 66.520 182.265 66.695 182.825 ;
        RECT 66.465 182.215 66.695 182.265 ;
        RECT 68.450 182.250 68.790 183.080 ;
        RECT 72.385 182.855 74.975 183.625 ;
        RECT 75.180 182.885 75.795 183.455 ;
        RECT 75.965 183.115 76.180 183.625 ;
        RECT 76.410 183.115 76.690 183.445 ;
        RECT 76.870 183.115 77.110 183.625 ;
        RECT 63.390 182.045 65.825 182.215 ;
        RECT 63.390 181.245 63.720 182.045 ;
        RECT 63.890 181.075 64.220 181.875 ;
        RECT 64.520 181.245 64.850 182.045 ;
        RECT 65.495 181.075 65.745 181.875 ;
        RECT 66.015 181.075 66.185 182.215 ;
        RECT 66.355 181.245 66.695 182.215 ;
        RECT 70.270 181.510 70.620 182.760 ;
        RECT 72.385 182.335 73.595 182.855 ;
        RECT 73.765 182.165 74.975 182.685 ;
        RECT 66.865 181.075 72.210 181.510 ;
        RECT 72.385 181.075 74.975 182.165 ;
        RECT 75.180 181.865 75.495 182.885 ;
        RECT 75.665 182.215 75.835 182.715 ;
        RECT 76.085 182.385 76.350 182.945 ;
        RECT 76.520 182.215 76.690 183.115 ;
        RECT 77.445 183.080 82.790 183.625 ;
        RECT 82.965 183.080 88.310 183.625 ;
        RECT 76.860 182.385 77.215 182.945 ;
        RECT 79.030 182.250 79.370 183.080 ;
        RECT 75.665 182.045 77.090 182.215 ;
        RECT 75.180 181.245 75.715 181.865 ;
        RECT 75.885 181.075 76.215 181.875 ;
        RECT 76.700 181.870 77.090 182.045 ;
        RECT 80.850 181.510 81.200 182.760 ;
        RECT 84.550 182.250 84.890 183.080 ;
        RECT 88.485 182.900 88.775 183.625 ;
        RECT 89.455 183.235 89.785 183.625 ;
        RECT 89.955 183.055 90.125 183.375 ;
        RECT 90.295 183.235 90.625 183.625 ;
        RECT 91.040 183.225 91.995 183.395 ;
        RECT 89.405 182.885 91.655 183.055 ;
        RECT 86.370 181.510 86.720 182.760 ;
        RECT 77.445 181.075 82.790 181.510 ;
        RECT 82.965 181.075 88.310 181.510 ;
        RECT 88.485 181.075 88.775 182.240 ;
        RECT 89.405 181.925 89.575 182.885 ;
        RECT 89.745 182.265 89.990 182.715 ;
        RECT 90.160 182.435 90.710 182.635 ;
        RECT 90.880 182.465 91.255 182.635 ;
        RECT 90.880 182.265 91.050 182.465 ;
        RECT 91.425 182.385 91.655 182.885 ;
        RECT 89.745 182.095 91.050 182.265 ;
        RECT 91.825 182.345 91.995 183.225 ;
        RECT 92.165 182.790 92.455 183.625 ;
        RECT 92.625 183.080 97.970 183.625 ;
        RECT 91.825 182.175 92.455 182.345 ;
        RECT 94.210 182.250 94.550 183.080 ;
        RECT 98.145 182.855 101.655 183.625 ;
        RECT 102.375 183.075 102.545 183.365 ;
        RECT 102.715 183.245 103.045 183.625 ;
        RECT 102.375 182.905 103.040 183.075 ;
        RECT 89.405 181.245 89.785 181.925 ;
        RECT 90.375 181.075 90.545 181.925 ;
        RECT 90.715 181.755 91.955 181.925 ;
        RECT 90.715 181.245 91.045 181.755 ;
        RECT 91.215 181.075 91.385 181.585 ;
        RECT 91.555 181.245 91.955 181.755 ;
        RECT 92.135 181.245 92.455 182.175 ;
        RECT 96.030 181.510 96.380 182.760 ;
        RECT 98.145 182.335 99.795 182.855 ;
        RECT 99.965 182.165 101.655 182.685 ;
        RECT 92.625 181.075 97.970 181.510 ;
        RECT 98.145 181.075 101.655 182.165 ;
        RECT 102.290 182.085 102.640 182.735 ;
        RECT 102.810 181.915 103.040 182.905 ;
        RECT 102.375 181.745 103.040 181.915 ;
        RECT 102.375 181.245 102.545 181.745 ;
        RECT 102.715 181.075 103.045 181.575 ;
        RECT 103.215 181.245 103.400 183.365 ;
        RECT 103.655 183.165 103.905 183.625 ;
        RECT 104.075 183.175 104.410 183.345 ;
        RECT 104.605 183.175 105.280 183.345 ;
        RECT 104.075 183.035 104.245 183.175 ;
        RECT 103.570 182.045 103.850 182.995 ;
        RECT 104.020 182.905 104.245 183.035 ;
        RECT 104.020 181.800 104.190 182.905 ;
        RECT 104.415 182.755 104.940 182.975 ;
        RECT 104.360 181.990 104.600 182.585 ;
        RECT 104.770 182.055 104.940 182.755 ;
        RECT 105.110 182.395 105.280 183.175 ;
        RECT 105.600 183.125 105.970 183.625 ;
        RECT 106.150 183.175 106.555 183.345 ;
        RECT 106.725 183.175 107.510 183.345 ;
        RECT 106.150 182.945 106.320 183.175 ;
        RECT 105.490 182.645 106.320 182.945 ;
        RECT 106.705 182.675 107.170 183.005 ;
        RECT 105.490 182.615 105.690 182.645 ;
        RECT 105.810 182.395 105.980 182.465 ;
        RECT 105.110 182.225 105.980 182.395 ;
        RECT 105.470 182.135 105.980 182.225 ;
        RECT 104.020 181.670 104.325 181.800 ;
        RECT 104.770 181.690 105.300 182.055 ;
        RECT 103.640 181.075 103.905 181.535 ;
        RECT 104.075 181.245 104.325 181.670 ;
        RECT 105.470 181.520 105.640 182.135 ;
        RECT 104.535 181.350 105.640 181.520 ;
        RECT 105.810 181.075 105.980 181.875 ;
        RECT 106.150 181.575 106.320 182.645 ;
        RECT 106.490 181.745 106.680 182.465 ;
        RECT 106.850 181.715 107.170 182.675 ;
        RECT 107.340 182.715 107.510 183.175 ;
        RECT 107.785 183.095 107.995 183.625 ;
        RECT 108.255 182.885 108.585 183.410 ;
        RECT 108.755 183.015 108.925 183.625 ;
        RECT 109.095 182.970 109.425 183.405 ;
        RECT 109.595 183.110 109.765 183.625 ;
        RECT 109.095 182.885 109.475 182.970 ;
        RECT 110.115 182.895 110.415 183.625 ;
        RECT 108.385 182.715 108.585 182.885 ;
        RECT 109.250 182.845 109.475 182.885 ;
        RECT 107.340 182.385 108.215 182.715 ;
        RECT 108.385 182.385 109.135 182.715 ;
        RECT 106.150 181.245 106.400 181.575 ;
        RECT 107.340 181.545 107.510 182.385 ;
        RECT 108.385 182.180 108.575 182.385 ;
        RECT 109.305 182.265 109.475 182.845 ;
        RECT 110.595 182.715 110.825 183.335 ;
        RECT 111.025 183.065 111.250 183.445 ;
        RECT 111.420 183.235 111.750 183.625 ;
        RECT 111.025 182.885 111.355 183.065 ;
        RECT 110.120 182.385 110.415 182.715 ;
        RECT 110.595 182.385 111.010 182.715 ;
        RECT 109.260 182.215 109.475 182.265 ;
        RECT 107.680 181.805 108.575 182.180 ;
        RECT 109.085 182.135 109.475 182.215 ;
        RECT 111.180 182.215 111.355 182.885 ;
        RECT 111.525 182.385 111.765 183.035 ;
        RECT 111.945 182.855 113.615 183.625 ;
        RECT 114.245 182.900 114.535 183.625 ;
        RECT 114.705 182.855 116.375 183.625 ;
        RECT 116.585 183.115 116.985 183.625 ;
        RECT 117.560 183.010 117.730 183.455 ;
        RECT 117.900 183.225 118.620 183.625 ;
        RECT 118.790 183.055 118.960 183.455 ;
        RECT 119.195 183.180 119.625 183.625 ;
        RECT 111.945 182.335 112.695 182.855 ;
        RECT 106.625 181.375 107.510 181.545 ;
        RECT 107.690 181.075 108.005 181.575 ;
        RECT 108.235 181.245 108.575 181.805 ;
        RECT 108.745 181.075 108.915 182.085 ;
        RECT 109.085 181.290 109.415 182.135 ;
        RECT 109.585 181.075 109.755 181.990 ;
        RECT 110.115 181.855 111.010 182.185 ;
        RECT 111.180 182.025 111.765 182.215 ;
        RECT 112.865 182.165 113.615 182.685 ;
        RECT 114.705 182.335 115.455 182.855 ;
        RECT 110.115 181.685 111.320 181.855 ;
        RECT 110.115 181.255 110.445 181.685 ;
        RECT 110.625 181.075 110.820 181.515 ;
        RECT 110.990 181.255 111.320 181.685 ;
        RECT 111.490 181.255 111.765 182.025 ;
        RECT 111.945 181.075 113.615 182.165 ;
        RECT 114.245 181.075 114.535 182.240 ;
        RECT 115.625 182.165 116.375 182.685 ;
        RECT 114.705 181.075 116.375 182.165 ;
        RECT 116.600 182.055 116.860 182.945 ;
        RECT 117.060 182.355 117.320 182.945 ;
        RECT 117.560 182.840 117.910 183.010 ;
        RECT 117.060 182.055 117.540 182.355 ;
        RECT 116.625 181.705 117.565 181.875 ;
        RECT 116.625 181.245 116.805 181.705 ;
        RECT 116.975 181.075 117.225 181.535 ;
        RECT 117.395 181.455 117.565 181.705 ;
        RECT 117.740 181.815 117.910 182.840 ;
        RECT 118.080 182.885 118.960 183.055 ;
        RECT 119.795 182.900 120.055 183.455 ;
        RECT 118.080 182.165 118.250 182.885 ;
        RECT 118.440 182.335 118.730 182.715 ;
        RECT 118.080 181.995 118.600 182.165 ;
        RECT 118.900 182.095 119.230 182.715 ;
        RECT 119.455 182.385 119.710 182.715 ;
        RECT 117.740 181.645 118.150 181.815 ;
        RECT 118.430 181.805 118.600 181.995 ;
        RECT 119.455 181.905 119.625 182.385 ;
        RECT 119.880 182.185 120.055 182.900 ;
        RECT 117.895 181.510 118.150 181.645 ;
        RECT 118.865 181.735 119.625 181.905 ;
        RECT 118.865 181.510 119.035 181.735 ;
        RECT 117.395 181.285 117.725 181.455 ;
        RECT 117.895 181.340 119.035 181.510 ;
        RECT 117.895 181.245 118.150 181.340 ;
        RECT 119.295 181.075 119.625 181.475 ;
        RECT 119.795 181.245 120.055 182.185 ;
        RECT 120.230 182.025 120.565 183.445 ;
        RECT 120.745 183.255 121.490 183.625 ;
        RECT 122.055 183.085 122.310 183.445 ;
        RECT 122.490 183.255 122.820 183.625 ;
        RECT 123.000 183.085 123.225 183.445 ;
        RECT 120.740 182.895 123.225 183.085 ;
        RECT 120.740 182.205 120.965 182.895 ;
        RECT 123.910 182.860 124.365 183.625 ;
        RECT 124.640 183.245 125.940 183.455 ;
        RECT 126.195 183.265 126.525 183.625 ;
        RECT 125.770 183.095 125.940 183.245 ;
        RECT 126.695 183.125 126.955 183.455 ;
        RECT 121.165 182.385 121.445 182.715 ;
        RECT 121.625 182.385 122.200 182.715 ;
        RECT 122.380 182.385 122.815 182.715 ;
        RECT 122.995 182.385 123.265 182.715 ;
        RECT 124.840 182.635 125.060 183.035 ;
        RECT 123.905 182.435 124.395 182.635 ;
        RECT 124.585 182.425 125.060 182.635 ;
        RECT 125.305 182.635 125.515 183.035 ;
        RECT 125.770 182.970 126.525 183.095 ;
        RECT 125.770 182.925 126.615 182.970 ;
        RECT 126.345 182.805 126.615 182.925 ;
        RECT 125.305 182.425 125.635 182.635 ;
        RECT 125.805 182.365 126.215 182.670 ;
        RECT 120.740 182.025 123.235 182.205 ;
        RECT 120.230 181.255 120.495 182.025 ;
        RECT 120.665 181.075 120.995 181.795 ;
        RECT 121.185 181.615 122.375 181.845 ;
        RECT 121.185 181.255 121.445 181.615 ;
        RECT 121.615 181.075 121.945 181.445 ;
        RECT 122.115 181.255 122.375 181.615 ;
        RECT 122.945 181.255 123.235 182.025 ;
        RECT 123.910 182.195 125.085 182.255 ;
        RECT 126.445 182.230 126.615 182.805 ;
        RECT 126.415 182.195 126.615 182.230 ;
        RECT 123.910 182.085 126.615 182.195 ;
        RECT 123.910 181.465 124.165 182.085 ;
        RECT 124.755 182.025 126.555 182.085 ;
        RECT 124.755 181.995 125.085 182.025 ;
        RECT 126.785 181.925 126.955 183.125 ;
        RECT 127.125 182.855 129.715 183.625 ;
        RECT 129.885 182.950 130.145 183.455 ;
        RECT 130.325 183.245 130.655 183.625 ;
        RECT 130.835 183.075 131.005 183.455 ;
        RECT 131.265 183.080 136.610 183.625 ;
        RECT 127.125 182.335 128.335 182.855 ;
        RECT 128.505 182.165 129.715 182.685 ;
        RECT 124.415 181.825 124.600 181.915 ;
        RECT 125.190 181.825 126.025 181.835 ;
        RECT 124.415 181.625 126.025 181.825 ;
        RECT 124.415 181.585 124.645 181.625 ;
        RECT 123.910 181.245 124.245 181.465 ;
        RECT 125.250 181.075 125.605 181.455 ;
        RECT 125.775 181.245 126.025 181.625 ;
        RECT 126.275 181.075 126.525 181.855 ;
        RECT 126.695 181.245 126.955 181.925 ;
        RECT 127.125 181.075 129.715 182.165 ;
        RECT 129.885 182.150 130.055 182.950 ;
        RECT 130.340 182.905 131.005 183.075 ;
        RECT 130.340 182.650 130.510 182.905 ;
        RECT 130.225 182.320 130.510 182.650 ;
        RECT 130.745 182.355 131.075 182.725 ;
        RECT 130.340 182.175 130.510 182.320 ;
        RECT 132.850 182.250 133.190 183.080 ;
        RECT 136.785 182.855 139.375 183.625 ;
        RECT 140.005 182.900 140.295 183.625 ;
        RECT 140.465 183.080 145.810 183.625 ;
        RECT 129.885 181.245 130.155 182.150 ;
        RECT 130.340 182.005 131.005 182.175 ;
        RECT 130.325 181.075 130.655 181.835 ;
        RECT 130.835 181.245 131.005 182.005 ;
        RECT 134.670 181.510 135.020 182.760 ;
        RECT 136.785 182.335 137.995 182.855 ;
        RECT 138.165 182.165 139.375 182.685 ;
        RECT 142.050 182.250 142.390 183.080 ;
        RECT 145.985 182.855 148.575 183.625 ;
        RECT 149.205 182.875 150.415 183.625 ;
        RECT 131.265 181.075 136.610 181.510 ;
        RECT 136.785 181.075 139.375 182.165 ;
        RECT 140.005 181.075 140.295 182.240 ;
        RECT 143.870 181.510 144.220 182.760 ;
        RECT 145.985 182.335 147.195 182.855 ;
        RECT 147.365 182.165 148.575 182.685 ;
        RECT 140.465 181.075 145.810 181.510 ;
        RECT 145.985 181.075 148.575 182.165 ;
        RECT 149.205 182.165 149.725 182.705 ;
        RECT 149.895 182.335 150.415 182.875 ;
        RECT 149.205 181.075 150.415 182.165 ;
        RECT 11.120 180.905 150.500 181.075 ;
        RECT 11.205 179.815 12.415 180.905 ;
        RECT 13.595 180.235 13.765 180.735 ;
        RECT 13.935 180.405 14.265 180.905 ;
        RECT 13.595 180.065 14.260 180.235 ;
        RECT 11.205 179.105 11.725 179.645 ;
        RECT 11.895 179.275 12.415 179.815 ;
        RECT 13.510 179.245 13.860 179.895 ;
        RECT 11.205 178.355 12.415 179.105 ;
        RECT 14.030 179.075 14.260 180.065 ;
        RECT 13.595 178.905 14.260 179.075 ;
        RECT 13.595 178.615 13.765 178.905 ;
        RECT 13.935 178.355 14.265 178.735 ;
        RECT 14.435 178.615 14.620 180.735 ;
        RECT 14.860 180.445 15.125 180.905 ;
        RECT 15.295 180.310 15.545 180.735 ;
        RECT 15.755 180.460 16.860 180.630 ;
        RECT 15.240 180.180 15.545 180.310 ;
        RECT 14.790 178.985 15.070 179.935 ;
        RECT 15.240 179.075 15.410 180.180 ;
        RECT 15.580 179.395 15.820 179.990 ;
        RECT 15.990 179.925 16.520 180.290 ;
        RECT 15.990 179.225 16.160 179.925 ;
        RECT 16.690 179.845 16.860 180.460 ;
        RECT 17.030 180.105 17.200 180.905 ;
        RECT 17.370 180.405 17.620 180.735 ;
        RECT 17.845 180.435 18.730 180.605 ;
        RECT 16.690 179.755 17.200 179.845 ;
        RECT 15.240 178.945 15.465 179.075 ;
        RECT 15.635 179.005 16.160 179.225 ;
        RECT 16.330 179.585 17.200 179.755 ;
        RECT 14.875 178.355 15.125 178.815 ;
        RECT 15.295 178.805 15.465 178.945 ;
        RECT 16.330 178.805 16.500 179.585 ;
        RECT 17.030 179.515 17.200 179.585 ;
        RECT 16.710 179.335 16.910 179.365 ;
        RECT 17.370 179.335 17.540 180.405 ;
        RECT 17.710 179.515 17.900 180.235 ;
        RECT 16.710 179.035 17.540 179.335 ;
        RECT 18.070 179.305 18.390 180.265 ;
        RECT 15.295 178.635 15.630 178.805 ;
        RECT 15.825 178.635 16.500 178.805 ;
        RECT 16.820 178.355 17.190 178.855 ;
        RECT 17.370 178.805 17.540 179.035 ;
        RECT 17.925 178.975 18.390 179.305 ;
        RECT 18.560 179.595 18.730 180.435 ;
        RECT 18.910 180.405 19.225 180.905 ;
        RECT 19.455 180.175 19.795 180.735 ;
        RECT 18.900 179.800 19.795 180.175 ;
        RECT 19.965 179.895 20.135 180.905 ;
        RECT 19.605 179.595 19.795 179.800 ;
        RECT 20.305 179.845 20.635 180.690 ;
        RECT 20.805 179.990 20.975 180.905 ;
        RECT 22.255 180.295 22.585 180.725 ;
        RECT 22.765 180.465 22.960 180.905 ;
        RECT 23.130 180.295 23.460 180.725 ;
        RECT 22.255 180.125 23.460 180.295 ;
        RECT 20.305 179.765 20.695 179.845 ;
        RECT 22.255 179.795 23.150 180.125 ;
        RECT 23.630 179.955 23.905 180.725 ;
        RECT 20.480 179.715 20.695 179.765 ;
        RECT 18.560 179.265 19.435 179.595 ;
        RECT 19.605 179.265 20.355 179.595 ;
        RECT 18.560 178.805 18.730 179.265 ;
        RECT 19.605 179.095 19.805 179.265 ;
        RECT 20.525 179.135 20.695 179.715 ;
        RECT 23.320 179.765 23.905 179.955 ;
        RECT 22.260 179.265 22.555 179.595 ;
        RECT 22.735 179.265 23.150 179.595 ;
        RECT 20.470 179.095 20.695 179.135 ;
        RECT 17.370 178.635 17.775 178.805 ;
        RECT 17.945 178.635 18.730 178.805 ;
        RECT 19.005 178.355 19.215 178.885 ;
        RECT 19.475 178.570 19.805 179.095 ;
        RECT 20.315 179.010 20.695 179.095 ;
        RECT 19.975 178.355 20.145 178.965 ;
        RECT 20.315 178.575 20.645 179.010 ;
        RECT 20.815 178.355 20.985 178.870 ;
        RECT 22.255 178.355 22.555 179.085 ;
        RECT 22.735 178.645 22.965 179.265 ;
        RECT 23.320 179.095 23.495 179.765 ;
        RECT 24.085 179.740 24.375 180.905 ;
        RECT 24.635 180.235 24.805 180.735 ;
        RECT 24.975 180.405 25.305 180.905 ;
        RECT 24.635 180.065 25.300 180.235 ;
        RECT 23.165 178.915 23.495 179.095 ;
        RECT 23.665 178.945 23.905 179.595 ;
        RECT 24.550 179.245 24.900 179.895 ;
        RECT 23.165 178.535 23.390 178.915 ;
        RECT 23.560 178.355 23.890 178.745 ;
        RECT 24.085 178.355 24.375 179.080 ;
        RECT 25.070 179.075 25.300 180.065 ;
        RECT 24.635 178.905 25.300 179.075 ;
        RECT 24.635 178.615 24.805 178.905 ;
        RECT 24.975 178.355 25.305 178.735 ;
        RECT 25.475 178.615 25.660 180.735 ;
        RECT 25.900 180.445 26.165 180.905 ;
        RECT 26.335 180.310 26.585 180.735 ;
        RECT 26.795 180.460 27.900 180.630 ;
        RECT 26.280 180.180 26.585 180.310 ;
        RECT 25.830 178.985 26.110 179.935 ;
        RECT 26.280 179.075 26.450 180.180 ;
        RECT 26.620 179.395 26.860 179.990 ;
        RECT 27.030 179.925 27.560 180.290 ;
        RECT 27.030 179.225 27.200 179.925 ;
        RECT 27.730 179.845 27.900 180.460 ;
        RECT 28.070 180.105 28.240 180.905 ;
        RECT 28.410 180.405 28.660 180.735 ;
        RECT 28.885 180.435 29.770 180.605 ;
        RECT 27.730 179.755 28.240 179.845 ;
        RECT 26.280 178.945 26.505 179.075 ;
        RECT 26.675 179.005 27.200 179.225 ;
        RECT 27.370 179.585 28.240 179.755 ;
        RECT 25.915 178.355 26.165 178.815 ;
        RECT 26.335 178.805 26.505 178.945 ;
        RECT 27.370 178.805 27.540 179.585 ;
        RECT 28.070 179.515 28.240 179.585 ;
        RECT 27.750 179.335 27.950 179.365 ;
        RECT 28.410 179.335 28.580 180.405 ;
        RECT 28.750 179.515 28.940 180.235 ;
        RECT 27.750 179.035 28.580 179.335 ;
        RECT 29.110 179.305 29.430 180.265 ;
        RECT 26.335 178.635 26.670 178.805 ;
        RECT 26.865 178.635 27.540 178.805 ;
        RECT 27.860 178.355 28.230 178.855 ;
        RECT 28.410 178.805 28.580 179.035 ;
        RECT 28.965 178.975 29.430 179.305 ;
        RECT 29.600 179.595 29.770 180.435 ;
        RECT 29.950 180.405 30.265 180.905 ;
        RECT 30.495 180.175 30.835 180.735 ;
        RECT 29.940 179.800 30.835 180.175 ;
        RECT 31.005 179.895 31.175 180.905 ;
        RECT 30.645 179.595 30.835 179.800 ;
        RECT 31.345 179.845 31.675 180.690 ;
        RECT 31.345 179.765 31.735 179.845 ;
        RECT 31.520 179.715 31.735 179.765 ;
        RECT 31.910 179.755 32.170 180.905 ;
        RECT 32.345 179.830 32.600 180.735 ;
        RECT 32.770 180.145 33.100 180.905 ;
        RECT 33.315 179.975 33.485 180.735 ;
        RECT 29.600 179.265 30.475 179.595 ;
        RECT 30.645 179.265 31.395 179.595 ;
        RECT 29.600 178.805 29.770 179.265 ;
        RECT 30.645 179.095 30.845 179.265 ;
        RECT 31.565 179.135 31.735 179.715 ;
        RECT 31.510 179.095 31.735 179.135 ;
        RECT 28.410 178.635 28.815 178.805 ;
        RECT 28.985 178.635 29.770 178.805 ;
        RECT 30.045 178.355 30.255 178.885 ;
        RECT 30.515 178.570 30.845 179.095 ;
        RECT 31.355 179.010 31.735 179.095 ;
        RECT 31.015 178.355 31.185 178.965 ;
        RECT 31.355 178.575 31.685 179.010 ;
        RECT 31.910 178.355 32.170 179.195 ;
        RECT 32.345 179.100 32.515 179.830 ;
        RECT 32.770 179.805 33.485 179.975 ;
        RECT 32.770 179.595 32.940 179.805 ;
        RECT 34.675 179.765 35.005 180.905 ;
        RECT 35.535 179.935 35.865 180.720 ;
        RECT 36.135 180.235 36.305 180.735 ;
        RECT 36.475 180.405 36.805 180.905 ;
        RECT 36.135 180.065 36.800 180.235 ;
        RECT 35.185 179.765 35.865 179.935 ;
        RECT 32.685 179.265 32.940 179.595 ;
        RECT 32.345 178.525 32.600 179.100 ;
        RECT 32.770 179.075 32.940 179.265 ;
        RECT 33.220 179.255 33.575 179.625 ;
        RECT 34.665 179.345 35.015 179.595 ;
        RECT 35.185 179.165 35.355 179.765 ;
        RECT 35.525 179.345 35.875 179.595 ;
        RECT 36.050 179.245 36.400 179.895 ;
        RECT 32.770 178.905 33.485 179.075 ;
        RECT 32.770 178.355 33.100 178.735 ;
        RECT 33.315 178.525 33.485 178.905 ;
        RECT 34.675 178.355 34.945 179.165 ;
        RECT 35.115 178.525 35.445 179.165 ;
        RECT 35.615 178.355 35.855 179.165 ;
        RECT 36.570 179.075 36.800 180.065 ;
        RECT 36.135 178.905 36.800 179.075 ;
        RECT 36.135 178.615 36.305 178.905 ;
        RECT 36.475 178.355 36.805 178.735 ;
        RECT 36.975 178.615 37.160 180.735 ;
        RECT 37.400 180.445 37.665 180.905 ;
        RECT 37.835 180.310 38.085 180.735 ;
        RECT 38.295 180.460 39.400 180.630 ;
        RECT 37.780 180.180 38.085 180.310 ;
        RECT 37.330 178.985 37.610 179.935 ;
        RECT 37.780 179.075 37.950 180.180 ;
        RECT 38.120 179.395 38.360 179.990 ;
        RECT 38.530 179.925 39.060 180.290 ;
        RECT 38.530 179.225 38.700 179.925 ;
        RECT 39.230 179.845 39.400 180.460 ;
        RECT 39.570 180.105 39.740 180.905 ;
        RECT 39.910 180.405 40.160 180.735 ;
        RECT 40.385 180.435 41.270 180.605 ;
        RECT 39.230 179.755 39.740 179.845 ;
        RECT 37.780 178.945 38.005 179.075 ;
        RECT 38.175 179.005 38.700 179.225 ;
        RECT 38.870 179.585 39.740 179.755 ;
        RECT 37.415 178.355 37.665 178.815 ;
        RECT 37.835 178.805 38.005 178.945 ;
        RECT 38.870 178.805 39.040 179.585 ;
        RECT 39.570 179.515 39.740 179.585 ;
        RECT 39.250 179.335 39.450 179.365 ;
        RECT 39.910 179.335 40.080 180.405 ;
        RECT 40.250 179.515 40.440 180.235 ;
        RECT 39.250 179.035 40.080 179.335 ;
        RECT 40.610 179.305 40.930 180.265 ;
        RECT 37.835 178.635 38.170 178.805 ;
        RECT 38.365 178.635 39.040 178.805 ;
        RECT 39.360 178.355 39.730 178.855 ;
        RECT 39.910 178.805 40.080 179.035 ;
        RECT 40.465 178.975 40.930 179.305 ;
        RECT 41.100 179.595 41.270 180.435 ;
        RECT 41.450 180.405 41.765 180.905 ;
        RECT 41.995 180.175 42.335 180.735 ;
        RECT 41.440 179.800 42.335 180.175 ;
        RECT 42.505 179.895 42.675 180.905 ;
        RECT 42.145 179.595 42.335 179.800 ;
        RECT 42.845 179.845 43.175 180.690 ;
        RECT 42.845 179.765 43.235 179.845 ;
        RECT 43.410 179.765 43.665 180.905 ;
        RECT 43.835 179.935 44.165 180.735 ;
        RECT 44.335 180.105 44.505 180.905 ;
        RECT 44.675 179.935 45.005 180.735 ;
        RECT 45.175 180.105 45.505 180.905 ;
        RECT 45.675 179.935 46.005 180.735 ;
        RECT 46.315 180.105 46.645 180.905 ;
        RECT 46.915 179.935 47.245 180.735 ;
        RECT 43.020 179.715 43.235 179.765 ;
        RECT 43.835 179.715 47.245 179.935 ;
        RECT 47.415 179.715 47.745 180.905 ;
        RECT 48.005 179.815 49.675 180.905 ;
        RECT 41.100 179.265 41.975 179.595 ;
        RECT 42.145 179.265 42.895 179.595 ;
        RECT 41.100 178.805 41.270 179.265 ;
        RECT 42.145 179.095 42.345 179.265 ;
        RECT 43.065 179.135 43.235 179.715 ;
        RECT 46.690 179.545 47.245 179.715 ;
        RECT 43.430 179.345 44.165 179.545 ;
        RECT 44.385 179.375 45.020 179.545 ;
        RECT 44.390 179.345 45.020 179.375 ;
        RECT 45.555 179.345 46.400 179.545 ;
        RECT 46.690 179.375 47.315 179.545 ;
        RECT 46.690 179.325 47.245 179.375 ;
        RECT 47.485 179.345 47.815 179.545 ;
        RECT 43.010 179.095 43.235 179.135 ;
        RECT 39.910 178.635 40.315 178.805 ;
        RECT 40.485 178.635 41.270 178.805 ;
        RECT 41.545 178.355 41.755 178.885 ;
        RECT 42.015 178.570 42.345 179.095 ;
        RECT 42.855 179.010 43.235 179.095 ;
        RECT 42.515 178.355 42.685 178.965 ;
        RECT 42.855 178.575 43.185 179.010 ;
        RECT 43.410 179.005 44.505 179.175 ;
        RECT 43.410 178.525 43.745 179.005 ;
        RECT 43.915 178.355 44.085 178.815 ;
        RECT 44.255 178.735 44.505 179.005 ;
        RECT 44.675 178.905 46.405 179.175 ;
        RECT 46.575 178.735 46.745 179.155 ;
        RECT 46.915 178.905 47.245 179.325 ;
        RECT 47.415 178.735 47.745 179.175 ;
        RECT 44.255 178.525 45.445 178.735 ;
        RECT 45.635 178.525 47.745 178.735 ;
        RECT 48.005 179.125 48.755 179.645 ;
        RECT 48.925 179.295 49.675 179.815 ;
        RECT 49.845 179.740 50.135 180.905 ;
        RECT 50.305 179.765 50.580 180.735 ;
        RECT 50.790 180.105 51.070 180.905 ;
        RECT 51.240 180.395 52.855 180.725 ;
        RECT 51.240 180.055 52.415 180.225 ;
        RECT 51.240 179.935 51.410 180.055 ;
        RECT 50.750 179.765 51.410 179.935 ;
        RECT 48.005 178.355 49.675 179.125 ;
        RECT 49.845 178.355 50.135 179.080 ;
        RECT 50.305 179.030 50.475 179.765 ;
        RECT 50.750 179.595 50.920 179.765 ;
        RECT 51.670 179.595 51.915 179.885 ;
        RECT 52.085 179.765 52.415 180.055 ;
        RECT 52.675 179.595 52.845 180.155 ;
        RECT 53.095 179.765 53.355 180.905 ;
        RECT 53.525 179.815 55.195 180.905 ;
        RECT 50.645 179.265 50.920 179.595 ;
        RECT 51.090 179.265 51.915 179.595 ;
        RECT 52.130 179.265 52.845 179.595 ;
        RECT 53.015 179.345 53.350 179.595 ;
        RECT 50.750 179.095 50.920 179.265 ;
        RECT 52.595 179.175 52.845 179.265 ;
        RECT 50.305 178.685 50.580 179.030 ;
        RECT 50.750 178.925 52.415 179.095 ;
        RECT 50.770 178.355 51.145 178.755 ;
        RECT 51.315 178.575 51.485 178.925 ;
        RECT 51.655 178.355 51.985 178.755 ;
        RECT 52.155 178.525 52.415 178.925 ;
        RECT 52.595 178.755 52.925 179.175 ;
        RECT 53.095 178.355 53.355 179.175 ;
        RECT 53.525 179.125 54.275 179.645 ;
        RECT 54.445 179.295 55.195 179.815 ;
        RECT 55.385 180.065 55.640 180.735 ;
        RECT 55.810 180.145 56.140 180.905 ;
        RECT 56.310 180.305 56.560 180.735 ;
        RECT 56.730 180.485 57.085 180.905 ;
        RECT 57.275 180.565 58.445 180.735 ;
        RECT 57.275 180.525 57.605 180.565 ;
        RECT 57.715 180.305 57.945 180.395 ;
        RECT 56.310 180.065 57.945 180.305 ;
        RECT 58.115 180.065 58.445 180.565 ;
        RECT 53.525 178.355 55.195 179.125 ;
        RECT 55.385 178.935 55.555 180.065 ;
        RECT 58.615 179.895 58.785 180.735 ;
        RECT 55.725 179.725 58.785 179.895 ;
        RECT 59.975 179.765 60.305 180.905 ;
        RECT 60.835 179.935 61.165 180.720 ;
        RECT 60.485 179.765 61.165 179.935 ;
        RECT 61.345 179.815 64.855 180.905 ;
        RECT 65.025 179.815 66.235 180.905 ;
        RECT 66.510 180.105 66.765 180.905 ;
        RECT 66.935 179.935 67.265 180.735 ;
        RECT 67.435 180.105 67.605 180.905 ;
        RECT 67.775 179.935 68.105 180.735 ;
        RECT 55.725 179.175 55.895 179.725 ;
        RECT 56.115 179.375 56.490 179.545 ;
        RECT 56.125 179.345 56.490 179.375 ;
        RECT 56.660 179.345 56.990 179.545 ;
        RECT 55.725 179.005 56.525 179.175 ;
        RECT 55.385 178.855 55.570 178.935 ;
        RECT 55.385 178.525 55.640 178.855 ;
        RECT 55.855 178.355 56.185 178.835 ;
        RECT 56.355 178.775 56.525 179.005 ;
        RECT 56.705 178.945 56.990 179.345 ;
        RECT 57.260 179.345 57.735 179.545 ;
        RECT 57.905 179.345 58.350 179.545 ;
        RECT 58.520 179.345 58.870 179.555 ;
        RECT 59.965 179.345 60.315 179.595 ;
        RECT 57.260 178.945 57.540 179.345 ;
        RECT 57.720 179.005 58.785 179.175 ;
        RECT 60.485 179.165 60.655 179.765 ;
        RECT 60.825 179.345 61.175 179.595 ;
        RECT 57.720 178.775 57.890 179.005 ;
        RECT 56.355 178.525 57.890 178.775 ;
        RECT 58.115 178.355 58.445 178.835 ;
        RECT 58.615 178.525 58.785 179.005 ;
        RECT 59.975 178.355 60.245 179.165 ;
        RECT 60.415 178.525 60.745 179.165 ;
        RECT 60.915 178.355 61.155 179.165 ;
        RECT 61.345 179.125 62.995 179.645 ;
        RECT 63.165 179.295 64.855 179.815 ;
        RECT 61.345 178.355 64.855 179.125 ;
        RECT 65.025 179.105 65.545 179.645 ;
        RECT 65.715 179.275 66.235 179.815 ;
        RECT 66.405 179.765 68.105 179.935 ;
        RECT 68.275 179.765 68.535 180.905 ;
        RECT 68.705 180.470 74.050 180.905 ;
        RECT 66.405 179.175 66.685 179.765 ;
        RECT 66.855 179.345 67.605 179.595 ;
        RECT 67.775 179.345 68.535 179.595 ;
        RECT 65.025 178.355 66.235 179.105 ;
        RECT 66.405 178.925 67.265 179.175 ;
        RECT 67.435 178.985 68.535 179.155 ;
        RECT 66.515 178.735 66.845 178.755 ;
        RECT 67.435 178.735 67.685 178.985 ;
        RECT 66.515 178.525 67.685 178.735 ;
        RECT 67.855 178.355 68.025 178.815 ;
        RECT 68.195 178.525 68.535 178.985 ;
        RECT 70.290 178.900 70.630 179.730 ;
        RECT 72.110 179.220 72.460 180.470 ;
        RECT 74.225 179.815 75.435 180.905 ;
        RECT 74.225 179.105 74.745 179.645 ;
        RECT 74.915 179.275 75.435 179.815 ;
        RECT 75.605 179.740 75.895 180.905 ;
        RECT 76.065 179.815 77.735 180.905 ;
        RECT 76.065 179.125 76.815 179.645 ;
        RECT 76.985 179.295 77.735 179.815 ;
        RECT 78.375 179.765 78.705 180.905 ;
        RECT 79.235 179.935 79.565 180.720 ;
        RECT 80.295 180.235 80.465 180.735 ;
        RECT 80.635 180.405 80.965 180.905 ;
        RECT 80.295 180.065 80.960 180.235 ;
        RECT 78.885 179.765 79.565 179.935 ;
        RECT 78.365 179.345 78.715 179.595 ;
        RECT 78.885 179.165 79.055 179.765 ;
        RECT 79.225 179.345 79.575 179.595 ;
        RECT 80.210 179.245 80.560 179.895 ;
        RECT 68.705 178.355 74.050 178.900 ;
        RECT 74.225 178.355 75.435 179.105 ;
        RECT 75.605 178.355 75.895 179.080 ;
        RECT 76.065 178.355 77.735 179.125 ;
        RECT 78.375 178.355 78.645 179.165 ;
        RECT 78.815 178.525 79.145 179.165 ;
        RECT 79.315 178.355 79.555 179.165 ;
        RECT 80.730 179.075 80.960 180.065 ;
        RECT 80.295 178.905 80.960 179.075 ;
        RECT 80.295 178.615 80.465 178.905 ;
        RECT 80.635 178.355 80.965 178.735 ;
        RECT 81.135 178.615 81.320 180.735 ;
        RECT 81.560 180.445 81.825 180.905 ;
        RECT 81.995 180.310 82.245 180.735 ;
        RECT 82.455 180.460 83.560 180.630 ;
        RECT 81.940 180.180 82.245 180.310 ;
        RECT 81.490 178.985 81.770 179.935 ;
        RECT 81.940 179.075 82.110 180.180 ;
        RECT 82.280 179.395 82.520 179.990 ;
        RECT 82.690 179.925 83.220 180.290 ;
        RECT 82.690 179.225 82.860 179.925 ;
        RECT 83.390 179.845 83.560 180.460 ;
        RECT 83.730 180.105 83.900 180.905 ;
        RECT 84.070 180.405 84.320 180.735 ;
        RECT 84.545 180.435 85.430 180.605 ;
        RECT 83.390 179.755 83.900 179.845 ;
        RECT 81.940 178.945 82.165 179.075 ;
        RECT 82.335 179.005 82.860 179.225 ;
        RECT 83.030 179.585 83.900 179.755 ;
        RECT 81.575 178.355 81.825 178.815 ;
        RECT 81.995 178.805 82.165 178.945 ;
        RECT 83.030 178.805 83.200 179.585 ;
        RECT 83.730 179.515 83.900 179.585 ;
        RECT 83.410 179.335 83.610 179.365 ;
        RECT 84.070 179.335 84.240 180.405 ;
        RECT 84.410 179.515 84.600 180.235 ;
        RECT 83.410 179.035 84.240 179.335 ;
        RECT 84.770 179.305 85.090 180.265 ;
        RECT 81.995 178.635 82.330 178.805 ;
        RECT 82.525 178.635 83.200 178.805 ;
        RECT 83.520 178.355 83.890 178.855 ;
        RECT 84.070 178.805 84.240 179.035 ;
        RECT 84.625 178.975 85.090 179.305 ;
        RECT 85.260 179.595 85.430 180.435 ;
        RECT 85.610 180.405 85.925 180.905 ;
        RECT 86.155 180.175 86.495 180.735 ;
        RECT 85.600 179.800 86.495 180.175 ;
        RECT 86.665 179.895 86.835 180.905 ;
        RECT 86.305 179.595 86.495 179.800 ;
        RECT 87.005 179.845 87.335 180.690 ;
        RECT 87.005 179.765 87.395 179.845 ;
        RECT 87.180 179.715 87.395 179.765 ;
        RECT 85.260 179.265 86.135 179.595 ;
        RECT 86.305 179.265 87.055 179.595 ;
        RECT 85.260 178.805 85.430 179.265 ;
        RECT 86.305 179.095 86.505 179.265 ;
        RECT 87.225 179.135 87.395 179.715 ;
        RECT 87.170 179.095 87.395 179.135 ;
        RECT 84.070 178.635 84.475 178.805 ;
        RECT 84.645 178.635 85.430 178.805 ;
        RECT 85.705 178.355 85.915 178.885 ;
        RECT 86.175 178.570 86.505 179.095 ;
        RECT 87.015 179.010 87.395 179.095 ;
        RECT 87.565 179.725 88.090 180.735 ;
        RECT 88.325 180.185 88.655 180.905 ;
        RECT 88.825 180.015 89.075 180.735 ;
        RECT 88.325 179.725 89.075 180.015 ;
        RECT 87.565 179.155 87.835 179.725 ;
        RECT 88.325 179.555 88.585 179.725 ;
        RECT 88.005 179.345 88.585 179.555 ;
        RECT 88.755 179.345 89.175 179.555 ;
        RECT 89.345 179.345 89.675 180.660 ;
        RECT 89.885 179.345 90.215 180.660 ;
        RECT 90.385 179.345 90.755 180.660 ;
        RECT 91.085 179.785 91.415 180.905 ;
        RECT 91.705 179.765 92.090 180.735 ;
        RECT 92.260 180.445 92.585 180.905 ;
        RECT 93.105 180.275 93.385 180.735 ;
        RECT 92.260 180.055 93.385 180.275 ;
        RECT 90.965 179.345 91.475 179.595 ;
        RECT 88.215 179.175 88.585 179.345 ;
        RECT 86.675 178.355 86.845 178.965 ;
        RECT 87.015 178.575 87.345 179.010 ;
        RECT 87.565 178.525 87.905 179.155 ;
        RECT 88.215 178.985 88.965 179.175 ;
        RECT 88.195 178.355 88.365 178.815 ;
        RECT 88.635 178.540 88.965 178.985 ;
        RECT 89.135 179.005 91.435 179.175 ;
        RECT 89.135 178.685 89.305 179.005 ;
        RECT 89.530 178.355 89.860 178.815 ;
        RECT 90.060 178.525 90.390 179.005 ;
        RECT 90.605 178.355 90.935 178.815 ;
        RECT 91.105 178.525 91.435 179.005 ;
        RECT 91.705 179.095 91.985 179.765 ;
        RECT 92.260 179.595 92.710 180.055 ;
        RECT 93.575 179.885 93.975 180.735 ;
        RECT 94.375 180.445 94.645 180.905 ;
        RECT 94.815 180.275 95.100 180.735 ;
        RECT 95.405 180.395 95.705 180.905 ;
        RECT 95.875 180.395 96.255 180.565 ;
        RECT 96.835 180.395 97.465 180.905 ;
        RECT 92.155 179.265 92.710 179.595 ;
        RECT 92.880 179.325 93.975 179.885 ;
        RECT 92.260 179.155 92.710 179.265 ;
        RECT 91.705 178.525 92.090 179.095 ;
        RECT 92.260 178.985 93.385 179.155 ;
        RECT 92.260 178.355 92.585 178.815 ;
        RECT 93.105 178.525 93.385 178.985 ;
        RECT 93.575 178.525 93.975 179.325 ;
        RECT 94.145 180.055 95.100 180.275 ;
        RECT 95.875 180.225 96.045 180.395 ;
        RECT 97.635 180.225 97.965 180.735 ;
        RECT 98.135 180.395 98.435 180.905 ;
        RECT 94.145 179.155 94.355 180.055 ;
        RECT 95.385 180.025 96.045 180.225 ;
        RECT 96.215 180.055 98.435 180.225 ;
        RECT 94.525 179.325 95.215 179.885 ;
        RECT 94.145 178.985 95.100 179.155 ;
        RECT 94.375 178.355 94.645 178.815 ;
        RECT 94.815 178.525 95.100 178.985 ;
        RECT 95.385 179.095 95.555 180.025 ;
        RECT 96.215 179.855 96.385 180.055 ;
        RECT 95.725 179.685 96.385 179.855 ;
        RECT 96.555 179.715 98.095 179.885 ;
        RECT 95.725 179.265 95.895 179.685 ;
        RECT 96.555 179.515 96.725 179.715 ;
        RECT 96.125 179.345 96.725 179.515 ;
        RECT 96.895 179.345 97.590 179.545 ;
        RECT 97.850 179.265 98.095 179.715 ;
        RECT 96.215 179.095 97.125 179.175 ;
        RECT 95.385 178.615 95.705 179.095 ;
        RECT 95.875 179.005 97.125 179.095 ;
        RECT 95.875 178.925 96.385 179.005 ;
        RECT 95.875 178.525 96.105 178.925 ;
        RECT 96.275 178.355 96.625 178.745 ;
        RECT 96.795 178.525 97.125 179.005 ;
        RECT 97.295 178.355 97.465 179.175 ;
        RECT 98.265 179.095 98.435 180.055 ;
        RECT 98.605 179.765 98.865 180.905 ;
        RECT 99.035 179.755 99.365 180.735 ;
        RECT 99.535 179.765 99.815 180.905 ;
        RECT 99.985 179.815 101.195 180.905 ;
        RECT 98.625 179.345 98.960 179.595 ;
        RECT 99.130 179.205 99.300 179.755 ;
        RECT 99.470 179.325 99.805 179.595 ;
        RECT 99.125 179.155 99.300 179.205 ;
        RECT 97.970 178.550 98.435 179.095 ;
        RECT 98.605 178.525 99.300 179.155 ;
        RECT 99.505 178.355 99.815 179.155 ;
        RECT 99.985 179.105 100.505 179.645 ;
        RECT 100.675 179.275 101.195 179.815 ;
        RECT 101.365 179.740 101.655 180.905 ;
        RECT 101.825 179.815 103.035 180.905 ;
        RECT 101.825 179.105 102.345 179.645 ;
        RECT 102.515 179.275 103.035 179.815 ;
        RECT 103.295 179.975 103.465 180.735 ;
        RECT 103.645 180.145 103.975 180.905 ;
        RECT 103.295 179.805 103.960 179.975 ;
        RECT 104.145 179.830 104.415 180.735 ;
        RECT 104.585 180.470 109.930 180.905 ;
        RECT 103.790 179.660 103.960 179.805 ;
        RECT 103.225 179.255 103.555 179.625 ;
        RECT 103.790 179.330 104.075 179.660 ;
        RECT 99.985 178.355 101.195 179.105 ;
        RECT 101.365 178.355 101.655 179.080 ;
        RECT 101.825 178.355 103.035 179.105 ;
        RECT 103.790 179.075 103.960 179.330 ;
        RECT 103.295 178.905 103.960 179.075 ;
        RECT 104.245 179.030 104.415 179.830 ;
        RECT 103.295 178.525 103.465 178.905 ;
        RECT 103.645 178.355 103.975 178.735 ;
        RECT 104.155 178.525 104.415 179.030 ;
        RECT 106.170 178.900 106.510 179.730 ;
        RECT 107.990 179.220 108.340 180.470 ;
        RECT 110.105 179.815 111.775 180.905 ;
        RECT 112.415 180.185 112.745 180.905 ;
        RECT 110.105 179.125 110.855 179.645 ;
        RECT 111.025 179.295 111.775 179.815 ;
        RECT 112.405 179.545 112.635 179.885 ;
        RECT 112.925 179.545 113.140 180.660 ;
        RECT 113.335 179.960 113.665 180.735 ;
        RECT 113.835 180.130 114.545 180.905 ;
        RECT 113.335 179.745 114.485 179.960 ;
        RECT 112.405 179.345 112.735 179.545 ;
        RECT 112.925 179.365 113.375 179.545 ;
        RECT 113.045 179.345 113.375 179.365 ;
        RECT 113.545 179.345 114.015 179.575 ;
        RECT 114.200 179.175 114.485 179.745 ;
        RECT 114.715 179.300 114.995 180.735 ;
        RECT 115.170 179.935 115.445 180.735 ;
        RECT 115.615 180.105 115.945 180.905 ;
        RECT 116.115 180.565 117.255 180.735 ;
        RECT 116.115 179.935 116.285 180.565 ;
        RECT 115.170 179.725 116.285 179.935 ;
        RECT 116.455 179.935 116.785 180.395 ;
        RECT 116.955 180.105 117.255 180.565 ;
        RECT 118.385 180.185 118.845 180.735 ;
        RECT 119.035 180.185 119.365 180.905 ;
        RECT 116.455 179.715 117.215 179.935 ;
        RECT 115.170 179.345 115.890 179.545 ;
        RECT 116.060 179.345 116.830 179.545 ;
        RECT 104.585 178.355 109.930 178.900 ;
        RECT 110.105 178.355 111.775 179.125 ;
        RECT 112.405 178.985 113.585 179.175 ;
        RECT 112.405 178.525 112.745 178.985 ;
        RECT 113.255 178.905 113.585 178.985 ;
        RECT 113.775 178.985 114.485 179.175 ;
        RECT 113.775 178.845 114.075 178.985 ;
        RECT 113.760 178.835 114.075 178.845 ;
        RECT 113.750 178.825 114.075 178.835 ;
        RECT 113.740 178.820 114.075 178.825 ;
        RECT 112.915 178.355 113.085 178.815 ;
        RECT 113.735 178.810 114.075 178.820 ;
        RECT 113.730 178.805 114.075 178.810 ;
        RECT 113.725 178.795 114.075 178.805 ;
        RECT 113.720 178.790 114.075 178.795 ;
        RECT 113.715 178.525 114.075 178.790 ;
        RECT 114.315 178.355 114.485 178.815 ;
        RECT 114.655 178.525 114.995 179.300 ;
        RECT 117.000 179.175 117.215 179.715 ;
        RECT 115.170 178.355 115.445 179.175 ;
        RECT 115.615 179.005 117.215 179.175 ;
        RECT 115.615 178.995 116.785 179.005 ;
        RECT 115.615 178.525 115.945 178.995 ;
        RECT 116.115 178.355 116.285 178.825 ;
        RECT 116.455 178.525 116.785 178.995 ;
        RECT 116.955 178.355 117.245 178.825 ;
        RECT 118.385 178.815 118.635 180.185 ;
        RECT 119.565 180.015 119.865 180.565 ;
        RECT 120.035 180.235 120.315 180.905 ;
        RECT 118.925 179.845 119.865 180.015 ;
        RECT 118.925 179.595 119.095 179.845 ;
        RECT 120.235 179.595 120.500 179.955 ;
        RECT 120.685 179.815 123.275 180.905 ;
        RECT 118.805 179.265 119.095 179.595 ;
        RECT 119.265 179.345 119.605 179.595 ;
        RECT 119.825 179.345 120.500 179.595 ;
        RECT 118.925 179.175 119.095 179.265 ;
        RECT 118.925 178.985 120.315 179.175 ;
        RECT 118.385 178.525 118.945 178.815 ;
        RECT 119.115 178.355 119.365 178.815 ;
        RECT 119.985 178.625 120.315 178.985 ;
        RECT 120.685 179.125 121.895 179.645 ;
        RECT 122.065 179.295 123.275 179.815 ;
        RECT 123.450 179.765 123.725 180.735 ;
        RECT 123.935 180.105 124.215 180.905 ;
        RECT 124.385 180.395 125.575 180.685 ;
        RECT 124.385 180.055 125.555 180.225 ;
        RECT 124.385 179.935 124.555 180.055 ;
        RECT 123.895 179.765 124.555 179.935 ;
        RECT 120.685 178.355 123.275 179.125 ;
        RECT 123.450 179.030 123.620 179.765 ;
        RECT 123.895 179.595 124.065 179.765 ;
        RECT 124.865 179.595 125.060 179.885 ;
        RECT 125.230 179.765 125.555 180.055 ;
        RECT 125.745 179.815 126.955 180.905 ;
        RECT 123.790 179.265 124.065 179.595 ;
        RECT 124.235 179.265 125.060 179.595 ;
        RECT 125.230 179.265 125.575 179.595 ;
        RECT 123.895 179.095 124.065 179.265 ;
        RECT 125.745 179.105 126.265 179.645 ;
        RECT 126.435 179.275 126.955 179.815 ;
        RECT 127.125 179.740 127.415 180.905 ;
        RECT 127.590 180.105 127.845 180.905 ;
        RECT 128.045 180.055 128.375 180.735 ;
        RECT 127.590 179.565 127.835 179.925 ;
        RECT 128.025 179.775 128.375 180.055 ;
        RECT 128.025 179.395 128.195 179.775 ;
        RECT 128.555 179.595 128.750 180.645 ;
        RECT 128.930 179.765 129.250 180.905 ;
        RECT 129.425 180.470 134.770 180.905 ;
        RECT 134.945 180.470 140.290 180.905 ;
        RECT 140.465 180.470 145.810 180.905 ;
        RECT 127.675 179.225 128.195 179.395 ;
        RECT 128.365 179.265 128.750 179.595 ;
        RECT 128.930 179.545 129.190 179.595 ;
        RECT 128.930 179.375 129.195 179.545 ;
        RECT 128.930 179.265 129.190 179.375 ;
        RECT 123.450 178.685 123.725 179.030 ;
        RECT 123.895 178.925 125.560 179.095 ;
        RECT 123.915 178.355 124.295 178.755 ;
        RECT 124.465 178.575 124.635 178.925 ;
        RECT 124.805 178.355 125.135 178.755 ;
        RECT 125.305 178.575 125.560 178.925 ;
        RECT 125.745 178.355 126.955 179.105 ;
        RECT 127.125 178.355 127.415 179.080 ;
        RECT 127.675 178.865 127.845 179.225 ;
        RECT 127.645 178.695 127.845 178.865 ;
        RECT 127.675 178.660 127.845 178.695 ;
        RECT 128.035 178.885 129.250 179.055 ;
        RECT 131.010 178.900 131.350 179.730 ;
        RECT 132.830 179.220 133.180 180.470 ;
        RECT 136.530 178.900 136.870 179.730 ;
        RECT 138.350 179.220 138.700 180.470 ;
        RECT 142.050 178.900 142.390 179.730 ;
        RECT 143.870 179.220 144.220 180.470 ;
        RECT 145.985 179.815 148.575 180.905 ;
        RECT 145.985 179.125 147.195 179.645 ;
        RECT 147.365 179.295 148.575 179.815 ;
        RECT 149.205 179.815 150.415 180.905 ;
        RECT 149.205 179.275 149.725 179.815 ;
        RECT 128.035 178.580 128.265 178.885 ;
        RECT 128.435 178.355 128.765 178.715 ;
        RECT 128.960 178.535 129.250 178.885 ;
        RECT 129.425 178.355 134.770 178.900 ;
        RECT 134.945 178.355 140.290 178.900 ;
        RECT 140.465 178.355 145.810 178.900 ;
        RECT 145.985 178.355 148.575 179.125 ;
        RECT 149.895 179.105 150.415 179.645 ;
        RECT 149.205 178.355 150.415 179.105 ;
        RECT 11.120 178.185 150.500 178.355 ;
        RECT 11.205 177.435 12.415 178.185 ;
        RECT 11.205 176.895 11.725 177.435 ;
        RECT 12.585 177.415 16.095 178.185 ;
        RECT 17.275 177.845 17.445 177.880 ;
        RECT 17.245 177.675 17.445 177.845 ;
        RECT 11.895 176.725 12.415 177.265 ;
        RECT 12.585 176.895 14.235 177.415 ;
        RECT 17.275 177.315 17.445 177.675 ;
        RECT 17.635 177.655 17.865 177.960 ;
        RECT 18.035 177.825 18.365 178.185 ;
        RECT 18.560 177.655 18.850 178.005 ;
        RECT 17.635 177.485 18.850 177.655 ;
        RECT 19.025 177.640 24.370 178.185 ;
        RECT 24.635 177.845 24.805 177.880 ;
        RECT 24.605 177.675 24.805 177.845 ;
        RECT 14.405 176.725 16.095 177.245 ;
        RECT 17.275 177.145 17.795 177.315 ;
        RECT 11.205 175.635 12.415 176.725 ;
        RECT 12.585 175.635 16.095 176.725 ;
        RECT 17.190 176.615 17.435 176.975 ;
        RECT 17.625 176.765 17.795 177.145 ;
        RECT 17.965 176.945 18.350 177.275 ;
        RECT 18.530 177.165 18.790 177.275 ;
        RECT 18.530 176.995 18.795 177.165 ;
        RECT 18.530 176.945 18.790 176.995 ;
        RECT 17.625 176.485 17.975 176.765 ;
        RECT 17.190 175.635 17.445 176.435 ;
        RECT 17.645 175.805 17.975 176.485 ;
        RECT 18.155 175.895 18.350 176.945 ;
        RECT 20.610 176.810 20.950 177.640 ;
        RECT 18.530 175.635 18.850 176.775 ;
        RECT 22.430 176.070 22.780 177.320 ;
        RECT 24.635 177.315 24.805 177.675 ;
        RECT 24.995 177.655 25.225 177.960 ;
        RECT 25.395 177.825 25.725 178.185 ;
        RECT 25.920 177.655 26.210 178.005 ;
        RECT 24.995 177.485 26.210 177.655 ;
        RECT 26.385 177.640 31.730 178.185 ;
        RECT 32.365 177.725 32.925 178.015 ;
        RECT 33.095 177.725 33.345 178.185 ;
        RECT 24.635 177.145 25.155 177.315 ;
        RECT 24.550 176.615 24.795 176.975 ;
        RECT 24.985 176.765 25.155 177.145 ;
        RECT 25.325 176.945 25.710 177.275 ;
        RECT 25.890 177.165 26.150 177.275 ;
        RECT 25.890 176.995 26.155 177.165 ;
        RECT 25.890 176.945 26.150 176.995 ;
        RECT 24.985 176.485 25.335 176.765 ;
        RECT 19.025 175.635 24.370 176.070 ;
        RECT 24.550 175.635 24.805 176.435 ;
        RECT 25.005 175.805 25.335 176.485 ;
        RECT 25.515 175.895 25.710 176.945 ;
        RECT 27.970 176.810 28.310 177.640 ;
        RECT 25.890 175.635 26.210 176.775 ;
        RECT 29.790 176.070 30.140 177.320 ;
        RECT 32.365 176.355 32.615 177.725 ;
        RECT 33.965 177.555 34.295 177.915 ;
        RECT 32.905 177.365 34.295 177.555 ;
        RECT 34.670 177.655 34.960 178.005 ;
        RECT 35.155 177.825 35.485 178.185 ;
        RECT 35.655 177.655 35.885 177.960 ;
        RECT 34.670 177.485 35.885 177.655 ;
        RECT 32.905 177.275 33.075 177.365 ;
        RECT 36.075 177.315 36.245 177.880 ;
        RECT 36.965 177.460 37.255 178.185 ;
        RECT 37.515 177.705 37.815 178.185 ;
        RECT 37.985 177.535 38.245 177.990 ;
        RECT 38.415 177.705 38.675 178.185 ;
        RECT 38.855 177.535 39.115 177.990 ;
        RECT 39.285 177.705 39.535 178.185 ;
        RECT 39.715 177.535 39.975 177.990 ;
        RECT 40.145 177.705 40.395 178.185 ;
        RECT 40.575 177.535 40.835 177.990 ;
        RECT 41.005 177.705 41.250 178.185 ;
        RECT 41.420 177.535 41.695 177.990 ;
        RECT 41.865 177.705 42.110 178.185 ;
        RECT 42.280 177.535 42.540 177.990 ;
        RECT 42.710 177.705 42.970 178.185 ;
        RECT 43.140 177.535 43.400 177.990 ;
        RECT 43.570 177.705 43.830 178.185 ;
        RECT 44.000 177.535 44.260 177.990 ;
        RECT 44.430 177.625 44.690 178.185 ;
        RECT 32.785 176.945 33.075 177.275 ;
        RECT 33.245 176.945 33.585 177.195 ;
        RECT 33.805 176.945 34.480 177.195 ;
        RECT 34.730 177.165 34.990 177.275 ;
        RECT 34.725 176.995 34.990 177.165 ;
        RECT 34.730 176.945 34.990 176.995 ;
        RECT 35.170 176.945 35.555 177.275 ;
        RECT 35.725 177.145 36.245 177.315 ;
        RECT 37.515 177.365 44.260 177.535 ;
        RECT 37.515 177.165 38.680 177.365 ;
        RECT 44.860 177.195 45.110 178.005 ;
        RECT 45.290 177.660 45.550 178.185 ;
        RECT 45.720 177.195 45.970 178.005 ;
        RECT 46.150 177.675 46.455 178.185 ;
        RECT 47.545 177.675 47.850 178.185 ;
        RECT 32.905 176.695 33.075 176.945 ;
        RECT 32.905 176.525 33.845 176.695 ;
        RECT 34.215 176.585 34.480 176.945 ;
        RECT 26.385 175.635 31.730 176.070 ;
        RECT 32.365 175.805 32.825 176.355 ;
        RECT 33.015 175.635 33.345 176.355 ;
        RECT 33.545 175.975 33.845 176.525 ;
        RECT 34.015 175.635 34.295 176.305 ;
        RECT 34.670 175.635 34.990 176.775 ;
        RECT 35.170 175.895 35.365 176.945 ;
        RECT 35.725 176.765 35.895 177.145 ;
        RECT 37.485 176.995 38.680 177.165 ;
        RECT 35.545 176.485 35.895 176.765 ;
        RECT 36.085 176.615 36.330 176.975 ;
        RECT 35.545 175.805 35.875 176.485 ;
        RECT 36.075 175.635 36.330 176.435 ;
        RECT 36.965 175.635 37.255 176.800 ;
        RECT 37.515 176.775 38.680 176.995 ;
        RECT 38.850 176.945 45.970 177.195 ;
        RECT 46.140 176.945 46.455 177.505 ;
        RECT 47.545 176.945 47.860 177.505 ;
        RECT 48.030 177.195 48.280 178.005 ;
        RECT 48.450 177.660 48.710 178.185 ;
        RECT 48.890 177.195 49.140 178.005 ;
        RECT 49.310 177.625 49.570 178.185 ;
        RECT 49.740 177.535 50.000 177.990 ;
        RECT 50.170 177.705 50.430 178.185 ;
        RECT 50.600 177.535 50.860 177.990 ;
        RECT 51.030 177.705 51.290 178.185 ;
        RECT 51.460 177.535 51.720 177.990 ;
        RECT 51.890 177.705 52.135 178.185 ;
        RECT 52.305 177.535 52.580 177.990 ;
        RECT 52.750 177.705 52.995 178.185 ;
        RECT 53.165 177.535 53.425 177.990 ;
        RECT 53.605 177.705 53.855 178.185 ;
        RECT 54.025 177.535 54.285 177.990 ;
        RECT 54.465 177.705 54.715 178.185 ;
        RECT 54.885 177.535 55.145 177.990 ;
        RECT 55.325 177.705 55.585 178.185 ;
        RECT 55.755 177.535 56.015 177.990 ;
        RECT 56.185 177.705 56.485 178.185 ;
        RECT 49.740 177.365 56.485 177.535 ;
        RECT 48.030 176.945 55.150 177.195 ;
        RECT 37.515 176.550 44.260 176.775 ;
        RECT 37.515 175.635 37.785 176.380 ;
        RECT 37.955 175.810 38.245 176.550 ;
        RECT 38.855 176.535 44.260 176.550 ;
        RECT 38.415 175.640 38.670 176.365 ;
        RECT 38.855 175.810 39.115 176.535 ;
        RECT 39.285 175.640 39.530 176.365 ;
        RECT 39.715 175.810 39.975 176.535 ;
        RECT 40.145 175.640 40.390 176.365 ;
        RECT 40.575 175.810 40.835 176.535 ;
        RECT 41.005 175.640 41.250 176.365 ;
        RECT 41.420 175.810 41.680 176.535 ;
        RECT 41.850 175.640 42.110 176.365 ;
        RECT 42.280 175.810 42.540 176.535 ;
        RECT 42.710 175.640 42.970 176.365 ;
        RECT 43.140 175.810 43.400 176.535 ;
        RECT 43.570 175.640 43.830 176.365 ;
        RECT 44.000 175.810 44.260 176.535 ;
        RECT 44.430 175.640 44.690 176.435 ;
        RECT 44.860 175.810 45.110 176.945 ;
        RECT 38.415 175.635 44.690 175.640 ;
        RECT 45.290 175.635 45.550 176.445 ;
        RECT 45.725 175.805 45.970 176.945 ;
        RECT 46.150 175.635 46.445 176.445 ;
        RECT 47.555 175.635 47.850 176.445 ;
        RECT 48.030 175.805 48.275 176.945 ;
        RECT 48.450 175.635 48.710 176.445 ;
        RECT 48.890 175.810 49.140 176.945 ;
        RECT 55.320 176.775 56.485 177.365 ;
        RECT 49.740 176.550 56.485 176.775 ;
        RECT 49.740 176.535 55.145 176.550 ;
        RECT 49.310 175.640 49.570 176.435 ;
        RECT 49.740 175.810 50.000 176.535 ;
        RECT 50.170 175.640 50.430 176.365 ;
        RECT 50.600 175.810 50.860 176.535 ;
        RECT 51.030 175.640 51.290 176.365 ;
        RECT 51.460 175.810 51.720 176.535 ;
        RECT 51.890 175.640 52.150 176.365 ;
        RECT 52.320 175.810 52.580 176.535 ;
        RECT 52.750 175.640 52.995 176.365 ;
        RECT 53.165 175.810 53.425 176.535 ;
        RECT 53.610 175.640 53.855 176.365 ;
        RECT 54.025 175.810 54.285 176.535 ;
        RECT 54.470 175.640 54.715 176.365 ;
        RECT 54.885 175.810 55.145 176.535 ;
        RECT 55.330 175.640 55.585 176.365 ;
        RECT 55.755 175.810 56.045 176.550 ;
        RECT 49.310 175.635 55.585 175.640 ;
        RECT 56.215 175.635 56.485 176.380 ;
        RECT 56.745 175.805 57.005 178.015 ;
        RECT 57.175 177.805 57.505 178.185 ;
        RECT 57.715 177.275 57.910 177.850 ;
        RECT 58.180 177.275 58.365 177.855 ;
        RECT 57.175 176.355 57.345 177.275 ;
        RECT 57.655 176.945 57.910 177.275 ;
        RECT 58.135 176.945 58.365 177.275 ;
        RECT 58.615 177.845 60.095 178.015 ;
        RECT 58.615 176.945 58.785 177.845 ;
        RECT 58.955 177.345 59.505 177.675 ;
        RECT 59.695 177.515 60.095 177.845 ;
        RECT 60.275 177.805 60.605 178.185 ;
        RECT 60.915 177.685 61.175 178.015 ;
        RECT 57.715 176.635 57.910 176.945 ;
        RECT 58.180 176.635 58.365 176.945 ;
        RECT 58.955 176.355 59.125 177.345 ;
        RECT 59.695 177.035 59.865 177.515 ;
        RECT 60.445 177.325 60.655 177.505 ;
        RECT 60.035 177.155 60.655 177.325 ;
        RECT 57.175 176.185 59.125 176.355 ;
        RECT 59.295 176.865 59.865 177.035 ;
        RECT 61.005 176.985 61.175 177.685 ;
        RECT 59.295 176.355 59.465 176.865 ;
        RECT 60.045 176.815 61.175 176.985 ;
        RECT 61.345 177.435 62.555 178.185 ;
        RECT 62.725 177.460 63.015 178.185 ;
        RECT 63.185 177.535 63.445 178.015 ;
        RECT 63.615 177.725 63.945 178.185 ;
        RECT 64.135 177.545 64.335 177.965 ;
        RECT 61.345 176.895 61.865 177.435 ;
        RECT 60.045 176.695 60.215 176.815 ;
        RECT 59.635 176.525 60.215 176.695 ;
        RECT 59.295 176.185 60.035 176.355 ;
        RECT 60.485 176.315 60.835 176.645 ;
        RECT 57.175 175.635 57.505 176.015 ;
        RECT 57.930 175.805 58.100 176.185 ;
        RECT 58.360 175.635 58.690 176.015 ;
        RECT 58.885 175.805 59.055 176.185 ;
        RECT 59.265 175.635 59.595 176.015 ;
        RECT 59.845 175.805 60.035 176.185 ;
        RECT 61.005 176.135 61.175 176.815 ;
        RECT 62.035 176.725 62.555 177.265 ;
        RECT 60.275 175.635 60.605 176.015 ;
        RECT 60.915 175.805 61.175 176.135 ;
        RECT 61.345 175.635 62.555 176.725 ;
        RECT 62.725 175.635 63.015 176.800 ;
        RECT 63.185 176.505 63.355 177.535 ;
        RECT 63.525 176.845 63.755 177.275 ;
        RECT 63.925 177.025 64.335 177.545 ;
        RECT 64.505 177.700 65.295 177.965 ;
        RECT 64.505 176.845 64.760 177.700 ;
        RECT 65.475 177.365 65.805 177.785 ;
        RECT 65.975 177.365 66.235 178.185 ;
        RECT 65.475 177.275 65.725 177.365 ;
        RECT 64.930 177.025 65.725 177.275 ;
        RECT 63.525 176.675 65.315 176.845 ;
        RECT 63.185 175.805 63.460 176.505 ;
        RECT 63.630 176.380 64.345 176.675 ;
        RECT 64.565 176.315 64.895 176.505 ;
        RECT 63.670 175.635 63.885 176.180 ;
        RECT 64.055 175.805 64.530 176.145 ;
        RECT 64.700 176.140 64.895 176.315 ;
        RECT 65.065 176.310 65.315 176.675 ;
        RECT 64.700 175.635 65.315 176.140 ;
        RECT 65.555 175.805 65.725 177.025 ;
        RECT 65.895 176.315 66.235 177.195 ;
        RECT 65.975 175.635 66.235 176.145 ;
        RECT 66.415 175.815 66.675 178.005 ;
        RECT 66.935 177.815 67.605 178.185 ;
        RECT 67.785 177.635 68.095 178.005 ;
        RECT 66.865 177.435 68.095 177.635 ;
        RECT 66.865 176.765 67.155 177.435 ;
        RECT 68.275 177.255 68.505 177.895 ;
        RECT 68.685 177.455 68.975 178.185 ;
        RECT 69.165 177.415 70.835 178.185 ;
        RECT 71.095 177.635 71.265 177.925 ;
        RECT 71.435 177.805 71.765 178.185 ;
        RECT 71.095 177.465 71.760 177.635 ;
        RECT 67.335 176.945 67.800 177.255 ;
        RECT 67.980 176.945 68.505 177.255 ;
        RECT 68.685 176.945 68.985 177.275 ;
        RECT 69.165 176.895 69.915 177.415 ;
        RECT 66.865 176.545 67.635 176.765 ;
        RECT 66.845 175.635 67.185 176.365 ;
        RECT 67.365 175.815 67.635 176.545 ;
        RECT 67.815 176.525 68.975 176.765 ;
        RECT 70.085 176.725 70.835 177.245 ;
        RECT 67.815 175.815 68.045 176.525 ;
        RECT 68.215 175.635 68.545 176.345 ;
        RECT 68.715 175.815 68.975 176.525 ;
        RECT 69.165 175.635 70.835 176.725 ;
        RECT 71.010 176.645 71.360 177.295 ;
        RECT 71.530 176.475 71.760 177.465 ;
        RECT 71.095 176.305 71.760 176.475 ;
        RECT 71.095 175.805 71.265 176.305 ;
        RECT 71.435 175.635 71.765 176.135 ;
        RECT 71.935 175.805 72.120 177.925 ;
        RECT 72.375 177.725 72.625 178.185 ;
        RECT 72.795 177.735 73.130 177.905 ;
        RECT 73.325 177.735 74.000 177.905 ;
        RECT 72.795 177.595 72.965 177.735 ;
        RECT 72.290 176.605 72.570 177.555 ;
        RECT 72.740 177.465 72.965 177.595 ;
        RECT 72.740 176.360 72.910 177.465 ;
        RECT 73.135 177.315 73.660 177.535 ;
        RECT 73.080 176.550 73.320 177.145 ;
        RECT 73.490 176.615 73.660 177.315 ;
        RECT 73.830 176.955 74.000 177.735 ;
        RECT 74.320 177.685 74.690 178.185 ;
        RECT 74.870 177.735 75.275 177.905 ;
        RECT 75.445 177.735 76.230 177.905 ;
        RECT 74.870 177.505 75.040 177.735 ;
        RECT 74.210 177.205 75.040 177.505 ;
        RECT 75.425 177.235 75.890 177.565 ;
        RECT 74.210 177.175 74.410 177.205 ;
        RECT 74.530 176.955 74.700 177.025 ;
        RECT 73.830 176.785 74.700 176.955 ;
        RECT 74.190 176.695 74.700 176.785 ;
        RECT 72.740 176.230 73.045 176.360 ;
        RECT 73.490 176.250 74.020 176.615 ;
        RECT 72.360 175.635 72.625 176.095 ;
        RECT 72.795 175.805 73.045 176.230 ;
        RECT 74.190 176.080 74.360 176.695 ;
        RECT 73.255 175.910 74.360 176.080 ;
        RECT 74.530 175.635 74.700 176.435 ;
        RECT 74.870 176.135 75.040 177.205 ;
        RECT 75.210 176.305 75.400 177.025 ;
        RECT 75.570 176.275 75.890 177.235 ;
        RECT 76.060 177.275 76.230 177.735 ;
        RECT 76.505 177.655 76.715 178.185 ;
        RECT 76.975 177.445 77.305 177.970 ;
        RECT 77.475 177.575 77.645 178.185 ;
        RECT 77.815 177.530 78.145 177.965 ;
        RECT 77.815 177.445 78.195 177.530 ;
        RECT 77.105 177.275 77.305 177.445 ;
        RECT 77.970 177.405 78.195 177.445 ;
        RECT 76.060 176.945 76.935 177.275 ;
        RECT 77.105 176.945 77.855 177.275 ;
        RECT 74.870 175.805 75.120 176.135 ;
        RECT 76.060 176.105 76.230 176.945 ;
        RECT 77.105 176.740 77.295 176.945 ;
        RECT 78.025 176.825 78.195 177.405 ;
        RECT 77.980 176.775 78.195 176.825 ;
        RECT 76.400 176.365 77.295 176.740 ;
        RECT 77.805 176.695 78.195 176.775 ;
        RECT 78.370 177.510 78.645 177.855 ;
        RECT 78.835 177.785 79.215 178.185 ;
        RECT 79.385 177.615 79.555 177.965 ;
        RECT 79.725 177.785 80.055 178.185 ;
        RECT 80.225 177.615 80.480 177.965 ;
        RECT 78.370 176.775 78.540 177.510 ;
        RECT 78.815 177.445 80.480 177.615 ;
        RECT 78.815 177.275 78.985 177.445 ;
        RECT 80.665 177.415 82.335 178.185 ;
        RECT 78.710 176.945 78.985 177.275 ;
        RECT 79.155 176.945 79.980 177.275 ;
        RECT 80.150 176.945 80.495 177.275 ;
        RECT 78.815 176.775 78.985 176.945 ;
        RECT 75.345 175.935 76.230 176.105 ;
        RECT 76.410 175.635 76.725 176.135 ;
        RECT 76.955 175.805 77.295 176.365 ;
        RECT 77.465 175.635 77.635 176.645 ;
        RECT 77.805 175.850 78.135 176.695 ;
        RECT 78.370 175.805 78.645 176.775 ;
        RECT 78.815 176.605 79.475 176.775 ;
        RECT 79.785 176.655 79.980 176.945 ;
        RECT 80.665 176.895 81.415 177.415 ;
        RECT 79.305 176.485 79.475 176.605 ;
        RECT 80.150 176.485 80.475 176.775 ;
        RECT 81.585 176.725 82.335 177.245 ;
        RECT 78.855 175.635 79.135 176.435 ;
        RECT 79.305 176.315 80.475 176.485 ;
        RECT 79.305 175.855 80.495 176.145 ;
        RECT 80.665 175.635 82.335 176.725 ;
        RECT 82.505 177.240 82.845 178.015 ;
        RECT 83.015 177.725 83.185 178.185 ;
        RECT 83.425 177.750 83.785 178.015 ;
        RECT 83.425 177.745 83.780 177.750 ;
        RECT 83.425 177.735 83.775 177.745 ;
        RECT 83.425 177.730 83.770 177.735 ;
        RECT 83.425 177.720 83.765 177.730 ;
        RECT 84.415 177.725 84.585 178.185 ;
        RECT 83.425 177.715 83.760 177.720 ;
        RECT 83.425 177.705 83.750 177.715 ;
        RECT 83.425 177.695 83.740 177.705 ;
        RECT 83.425 177.555 83.725 177.695 ;
        RECT 83.015 177.365 83.725 177.555 ;
        RECT 83.915 177.555 84.245 177.635 ;
        RECT 84.755 177.555 85.095 178.015 ;
        RECT 83.915 177.365 85.095 177.555 ;
        RECT 85.265 177.415 87.855 178.185 ;
        RECT 88.485 177.460 88.775 178.185 ;
        RECT 88.945 177.415 90.615 178.185 ;
        RECT 91.250 177.930 91.585 177.975 ;
        RECT 91.245 177.465 91.585 177.930 ;
        RECT 91.755 177.805 92.085 178.185 ;
        RECT 82.505 175.805 82.785 177.240 ;
        RECT 83.015 176.795 83.300 177.365 ;
        RECT 83.485 176.965 83.955 177.195 ;
        RECT 84.125 177.175 84.455 177.195 ;
        RECT 84.125 176.995 84.575 177.175 ;
        RECT 84.765 176.995 85.095 177.195 ;
        RECT 83.015 176.580 84.165 176.795 ;
        RECT 82.955 175.635 83.665 176.410 ;
        RECT 83.835 175.805 84.165 176.580 ;
        RECT 84.360 175.880 84.575 176.995 ;
        RECT 84.865 176.655 85.095 176.995 ;
        RECT 85.265 176.895 86.475 177.415 ;
        RECT 86.645 176.725 87.855 177.245 ;
        RECT 88.945 176.895 89.695 177.415 ;
        RECT 84.755 175.635 85.085 176.355 ;
        RECT 85.265 175.635 87.855 176.725 ;
        RECT 88.485 175.635 88.775 176.800 ;
        RECT 89.865 176.725 90.615 177.245 ;
        RECT 88.945 175.635 90.615 176.725 ;
        RECT 91.245 176.775 91.415 177.465 ;
        RECT 91.585 176.945 91.845 177.275 ;
        RECT 91.245 175.805 91.505 176.775 ;
        RECT 91.675 176.395 91.845 176.945 ;
        RECT 92.015 176.575 92.355 177.605 ;
        RECT 92.545 176.825 92.815 177.850 ;
        RECT 92.545 176.655 92.855 176.825 ;
        RECT 92.545 176.575 92.815 176.655 ;
        RECT 93.040 176.575 93.320 177.850 ;
        RECT 93.520 177.685 93.750 178.015 ;
        RECT 93.995 177.805 94.325 178.185 ;
        RECT 93.520 176.395 93.690 177.685 ;
        RECT 94.495 177.615 94.670 178.015 ;
        RECT 94.040 177.445 94.670 177.615 ;
        RECT 94.040 177.275 94.210 177.445 ;
        RECT 94.935 177.375 95.205 178.185 ;
        RECT 95.375 177.375 95.705 178.015 ;
        RECT 95.875 177.375 96.115 178.185 ;
        RECT 96.305 177.415 99.815 178.185 ;
        RECT 99.990 177.680 100.325 178.185 ;
        RECT 100.495 177.615 100.735 177.990 ;
        RECT 101.015 177.855 101.185 178.000 ;
        RECT 101.015 177.660 101.390 177.855 ;
        RECT 101.750 177.690 102.145 178.185 ;
        RECT 93.860 176.945 94.210 177.275 ;
        RECT 91.675 176.225 93.690 176.395 ;
        RECT 94.040 176.425 94.210 176.945 ;
        RECT 94.390 176.595 94.755 177.275 ;
        RECT 94.925 176.945 95.275 177.195 ;
        RECT 95.445 176.775 95.615 177.375 ;
        RECT 95.785 176.945 96.135 177.195 ;
        RECT 96.305 176.895 97.955 177.415 ;
        RECT 94.040 176.255 94.670 176.425 ;
        RECT 91.700 175.635 92.030 176.045 ;
        RECT 92.230 175.805 92.400 176.225 ;
        RECT 92.615 175.635 93.285 176.045 ;
        RECT 93.520 175.805 93.690 176.225 ;
        RECT 93.995 175.635 94.325 176.075 ;
        RECT 94.495 175.805 94.670 176.255 ;
        RECT 94.935 175.635 95.265 176.775 ;
        RECT 95.445 176.605 96.125 176.775 ;
        RECT 98.125 176.725 99.815 177.245 ;
        RECT 95.795 175.820 96.125 176.605 ;
        RECT 96.305 175.635 99.815 176.725 ;
        RECT 100.045 176.655 100.345 177.505 ;
        RECT 100.515 177.465 100.735 177.615 ;
        RECT 100.515 177.135 101.050 177.465 ;
        RECT 101.220 177.325 101.390 177.660 ;
        RECT 102.315 177.495 102.555 178.015 ;
        RECT 100.515 176.485 100.750 177.135 ;
        RECT 101.220 176.965 102.205 177.325 ;
        RECT 100.075 176.255 100.750 176.485 ;
        RECT 100.920 176.945 102.205 176.965 ;
        RECT 100.920 176.795 101.780 176.945 ;
        RECT 100.075 175.825 100.245 176.255 ;
        RECT 100.415 175.635 100.745 176.085 ;
        RECT 100.920 175.850 101.205 176.795 ;
        RECT 102.380 176.690 102.555 177.495 ;
        RECT 101.380 176.315 102.075 176.625 ;
        RECT 101.385 175.635 102.070 176.105 ;
        RECT 102.250 175.905 102.555 176.690 ;
        RECT 102.745 177.710 103.085 177.970 ;
        RECT 102.745 176.105 103.005 177.710 ;
        RECT 103.255 177.705 103.585 178.185 ;
        RECT 103.775 177.535 104.190 177.970 ;
        RECT 104.360 177.670 105.310 177.855 ;
        RECT 103.175 177.460 104.190 177.535 ;
        RECT 103.175 177.365 103.995 177.460 ;
        RECT 103.175 176.445 103.345 177.365 ;
        RECT 103.665 176.635 103.995 177.195 ;
        RECT 104.195 177.165 104.575 177.275 ;
        RECT 104.185 176.995 104.575 177.165 ;
        RECT 104.195 176.945 104.575 176.995 ;
        RECT 104.885 176.945 105.105 177.670 ;
        RECT 105.540 177.275 105.745 177.875 ;
        RECT 105.915 177.460 106.255 178.185 ;
        RECT 106.430 177.710 106.765 177.970 ;
        RECT 106.935 177.785 107.265 178.185 ;
        RECT 107.435 177.785 109.050 177.955 ;
        RECT 104.195 176.650 104.495 176.945 ;
        RECT 105.365 176.645 105.745 177.275 ;
        RECT 105.975 176.645 106.230 177.275 ;
        RECT 103.175 176.275 104.025 176.445 ;
        RECT 102.745 175.845 103.085 176.105 ;
        RECT 103.255 175.635 103.505 176.095 ;
        RECT 103.695 175.845 104.025 176.275 ;
        RECT 104.195 176.305 106.165 176.475 ;
        RECT 104.195 175.805 104.365 176.305 ;
        RECT 104.575 175.635 104.825 176.095 ;
        RECT 105.035 175.805 105.205 176.305 ;
        RECT 105.505 175.635 105.755 176.095 ;
        RECT 105.995 175.805 106.165 176.305 ;
        RECT 106.430 176.355 106.685 177.710 ;
        RECT 107.435 177.615 107.605 177.785 ;
        RECT 107.045 177.445 107.605 177.615 ;
        RECT 107.870 177.505 108.140 177.605 ;
        RECT 107.045 177.275 107.215 177.445 ;
        RECT 107.865 177.335 108.140 177.505 ;
        RECT 106.910 176.945 107.215 177.275 ;
        RECT 107.410 177.165 107.660 177.275 ;
        RECT 107.405 176.995 107.660 177.165 ;
        RECT 107.410 176.945 107.660 176.995 ;
        RECT 107.870 176.945 108.140 177.335 ;
        RECT 108.330 176.945 108.620 177.605 ;
        RECT 108.790 176.945 109.210 177.610 ;
        RECT 109.595 177.465 109.925 178.185 ;
        RECT 110.105 177.415 113.615 178.185 ;
        RECT 114.245 177.460 114.535 178.185 ;
        RECT 114.705 177.415 117.295 178.185 ;
        RECT 109.520 177.165 109.870 177.275 ;
        RECT 109.520 176.995 109.875 177.165 ;
        RECT 109.520 176.945 109.870 176.995 ;
        RECT 107.045 176.775 107.215 176.945 ;
        RECT 107.045 176.605 109.415 176.775 ;
        RECT 109.665 176.655 109.870 176.945 ;
        RECT 110.105 176.895 111.755 177.415 ;
        RECT 111.925 176.725 113.615 177.245 ;
        RECT 114.705 176.895 115.915 177.415 ;
        RECT 117.485 177.375 117.725 178.185 ;
        RECT 117.895 177.375 118.225 178.015 ;
        RECT 118.395 177.375 118.665 178.185 ;
        RECT 118.845 177.415 121.435 178.185 ;
        RECT 106.430 175.845 106.765 176.355 ;
        RECT 107.015 175.635 107.345 176.435 ;
        RECT 107.590 176.225 109.015 176.395 ;
        RECT 107.590 175.805 107.875 176.225 ;
        RECT 108.130 175.635 108.460 176.055 ;
        RECT 108.685 175.975 109.015 176.225 ;
        RECT 109.245 176.145 109.415 176.605 ;
        RECT 109.675 175.975 109.845 176.475 ;
        RECT 108.685 175.805 109.845 175.975 ;
        RECT 110.105 175.635 113.615 176.725 ;
        RECT 114.245 175.635 114.535 176.800 ;
        RECT 116.085 176.725 117.295 177.245 ;
        RECT 117.465 176.945 117.815 177.195 ;
        RECT 117.985 176.775 118.155 177.375 ;
        RECT 118.325 176.945 118.675 177.195 ;
        RECT 118.845 176.895 120.055 177.415 ;
        RECT 114.705 175.635 117.295 176.725 ;
        RECT 117.475 176.605 118.155 176.775 ;
        RECT 117.475 175.820 117.805 176.605 ;
        RECT 118.335 175.635 118.665 176.775 ;
        RECT 120.225 176.725 121.435 177.245 ;
        RECT 118.845 175.635 121.435 176.725 ;
        RECT 122.085 176.605 122.315 177.945 ;
        RECT 122.495 177.105 122.725 178.005 ;
        RECT 122.925 177.405 123.170 178.185 ;
        RECT 123.340 177.645 123.770 178.005 ;
        RECT 124.350 177.815 125.080 178.185 ;
        RECT 123.340 177.455 125.080 177.645 ;
        RECT 123.340 177.225 123.560 177.455 ;
        RECT 122.495 176.425 122.835 177.105 ;
        RECT 122.085 176.225 122.835 176.425 ;
        RECT 123.015 176.925 123.560 177.225 ;
        RECT 122.085 175.835 122.325 176.225 ;
        RECT 122.495 175.635 122.845 176.045 ;
        RECT 123.015 175.815 123.345 176.925 ;
        RECT 123.730 176.655 124.155 177.275 ;
        RECT 124.350 176.655 124.610 177.275 ;
        RECT 124.820 176.945 125.080 177.455 ;
        RECT 123.515 176.285 124.540 176.485 ;
        RECT 123.515 175.815 123.695 176.285 ;
        RECT 123.865 175.635 124.195 176.115 ;
        RECT 124.370 175.815 124.540 176.285 ;
        RECT 124.805 175.635 125.090 176.775 ;
        RECT 125.280 175.815 125.560 178.005 ;
        RECT 125.745 177.640 131.090 178.185 ;
        RECT 131.265 177.640 136.610 178.185 ;
        RECT 127.330 176.810 127.670 177.640 ;
        RECT 129.150 176.070 129.500 177.320 ;
        RECT 132.850 176.810 133.190 177.640 ;
        RECT 136.785 177.415 139.375 178.185 ;
        RECT 140.005 177.460 140.295 178.185 ;
        RECT 140.465 177.640 145.810 178.185 ;
        RECT 134.670 176.070 135.020 177.320 ;
        RECT 136.785 176.895 137.995 177.415 ;
        RECT 138.165 176.725 139.375 177.245 ;
        RECT 142.050 176.810 142.390 177.640 ;
        RECT 145.985 177.415 148.575 178.185 ;
        RECT 149.205 177.435 150.415 178.185 ;
        RECT 125.745 175.635 131.090 176.070 ;
        RECT 131.265 175.635 136.610 176.070 ;
        RECT 136.785 175.635 139.375 176.725 ;
        RECT 140.005 175.635 140.295 176.800 ;
        RECT 143.870 176.070 144.220 177.320 ;
        RECT 145.985 176.895 147.195 177.415 ;
        RECT 147.365 176.725 148.575 177.245 ;
        RECT 140.465 175.635 145.810 176.070 ;
        RECT 145.985 175.635 148.575 176.725 ;
        RECT 149.205 176.725 149.725 177.265 ;
        RECT 149.895 176.895 150.415 177.435 ;
        RECT 149.205 175.635 150.415 176.725 ;
        RECT 11.120 175.465 150.500 175.635 ;
        RECT 11.205 174.375 12.415 175.465 ;
        RECT 12.585 174.375 16.095 175.465 ;
        RECT 11.205 173.665 11.725 174.205 ;
        RECT 11.895 173.835 12.415 174.375 ;
        RECT 12.585 173.685 14.235 174.205 ;
        RECT 14.405 173.855 16.095 174.375 ;
        RECT 16.265 174.390 16.535 175.295 ;
        RECT 16.705 174.705 17.035 175.465 ;
        RECT 17.215 174.535 17.385 175.295 ;
        RECT 17.645 175.030 22.990 175.465 ;
        RECT 11.205 172.915 12.415 173.665 ;
        RECT 12.585 172.915 16.095 173.685 ;
        RECT 16.265 173.590 16.435 174.390 ;
        RECT 16.720 174.365 17.385 174.535 ;
        RECT 16.720 174.220 16.890 174.365 ;
        RECT 16.605 173.890 16.890 174.220 ;
        RECT 16.720 173.635 16.890 173.890 ;
        RECT 17.125 173.815 17.455 174.185 ;
        RECT 16.265 173.085 16.525 173.590 ;
        RECT 16.720 173.465 17.385 173.635 ;
        RECT 16.705 172.915 17.035 173.295 ;
        RECT 17.215 173.085 17.385 173.465 ;
        RECT 19.230 173.460 19.570 174.290 ;
        RECT 21.050 173.780 21.400 175.030 ;
        RECT 24.085 174.300 24.375 175.465 ;
        RECT 24.545 175.030 29.890 175.465 ;
        RECT 30.065 175.030 35.410 175.465 ;
        RECT 17.645 172.915 22.990 173.460 ;
        RECT 24.085 172.915 24.375 173.640 ;
        RECT 26.130 173.460 26.470 174.290 ;
        RECT 27.950 173.780 28.300 175.030 ;
        RECT 31.650 173.460 31.990 174.290 ;
        RECT 33.470 173.780 33.820 175.030 ;
        RECT 35.585 174.375 37.255 175.465 ;
        RECT 35.585 173.685 36.335 174.205 ;
        RECT 36.505 173.855 37.255 174.375 ;
        RECT 37.435 174.495 37.765 175.280 ;
        RECT 37.435 174.325 38.115 174.495 ;
        RECT 38.295 174.325 38.625 175.465 ;
        RECT 38.805 174.375 41.395 175.465 ;
        RECT 42.035 175.085 42.365 175.465 ;
        RECT 37.425 173.905 37.775 174.155 ;
        RECT 37.945 173.725 38.115 174.325 ;
        RECT 38.285 173.905 38.635 174.155 ;
        RECT 24.545 172.915 29.890 173.460 ;
        RECT 30.065 172.915 35.410 173.460 ;
        RECT 35.585 172.915 37.255 173.685 ;
        RECT 37.445 172.915 37.685 173.725 ;
        RECT 37.855 173.085 38.185 173.725 ;
        RECT 38.355 172.915 38.625 173.725 ;
        RECT 38.805 173.685 40.015 174.205 ;
        RECT 40.185 173.855 41.395 174.375 ;
        RECT 38.805 172.915 41.395 173.685 ;
        RECT 42.065 173.585 42.270 174.905 ;
        RECT 42.540 174.495 42.790 175.295 ;
        RECT 43.010 174.745 43.340 175.465 ;
        RECT 43.525 174.495 43.775 175.295 ;
        RECT 44.175 174.665 44.505 175.465 ;
        RECT 42.440 174.325 44.495 174.495 ;
        RECT 44.675 174.325 45.010 175.295 ;
        RECT 45.185 174.665 45.515 175.465 ;
        RECT 45.705 174.375 49.215 175.465 ;
        RECT 42.440 173.415 42.610 174.325 ;
        RECT 42.115 173.085 42.610 173.415 ;
        RECT 42.830 173.250 43.185 174.155 ;
        RECT 43.360 174.135 43.530 174.155 ;
        RECT 43.360 173.245 43.660 174.135 ;
        RECT 43.840 173.245 44.100 174.155 ;
        RECT 44.270 174.145 44.495 174.325 ;
        RECT 44.270 173.905 44.665 174.145 ;
        RECT 44.835 173.765 45.010 174.325 ;
        RECT 44.270 172.915 44.505 173.720 ;
        RECT 44.835 173.635 45.015 173.765 ;
        RECT 45.705 173.685 47.355 174.205 ;
        RECT 47.525 173.855 49.215 174.375 ;
        RECT 49.845 174.300 50.135 175.465 ;
        RECT 50.505 174.795 50.785 175.465 ;
        RECT 50.955 174.575 51.255 175.125 ;
        RECT 51.455 174.745 51.785 175.465 ;
        RECT 51.975 174.745 52.435 175.295 ;
        RECT 50.320 174.155 50.585 174.515 ;
        RECT 50.955 174.405 51.895 174.575 ;
        RECT 51.725 174.155 51.895 174.405 ;
        RECT 50.320 173.905 50.995 174.155 ;
        RECT 51.215 173.905 51.555 174.155 ;
        RECT 51.725 173.825 52.015 174.155 ;
        RECT 51.725 173.735 51.895 173.825 ;
        RECT 44.675 173.595 45.015 173.635 ;
        RECT 44.675 173.170 45.010 173.595 ;
        RECT 44.675 173.125 45.005 173.170 ;
        RECT 45.195 172.915 45.525 173.640 ;
        RECT 45.705 172.915 49.215 173.685 ;
        RECT 49.845 172.915 50.135 173.640 ;
        RECT 50.505 173.545 51.895 173.735 ;
        RECT 50.505 173.185 50.835 173.545 ;
        RECT 52.185 173.375 52.435 174.745 ;
        RECT 52.645 175.125 53.785 175.295 ;
        RECT 52.645 174.665 52.945 175.125 ;
        RECT 53.115 174.495 53.445 174.955 ;
        RECT 52.685 174.275 53.445 174.495 ;
        RECT 53.615 174.495 53.785 175.125 ;
        RECT 53.955 174.665 54.285 175.465 ;
        RECT 54.455 174.495 54.730 175.295 ;
        RECT 53.615 174.285 54.730 174.495 ;
        RECT 54.910 174.325 55.230 175.465 ;
        RECT 52.685 173.735 52.900 174.275 ;
        RECT 55.410 174.155 55.605 175.205 ;
        RECT 55.785 174.615 56.115 175.295 ;
        RECT 56.315 174.665 56.570 175.465 ;
        RECT 56.745 175.030 62.090 175.465 ;
        RECT 55.785 174.335 56.135 174.615 ;
        RECT 54.970 174.105 55.230 174.155 ;
        RECT 53.070 173.905 53.840 174.105 ;
        RECT 54.010 173.905 54.730 174.105 ;
        RECT 54.965 173.935 55.230 174.105 ;
        RECT 54.970 173.825 55.230 173.935 ;
        RECT 55.410 173.825 55.795 174.155 ;
        RECT 55.965 173.955 56.135 174.335 ;
        RECT 56.325 174.125 56.570 174.485 ;
        RECT 55.965 173.785 56.485 173.955 ;
        RECT 52.685 173.565 54.285 173.735 ;
        RECT 53.115 173.555 54.285 173.565 ;
        RECT 51.455 172.915 51.705 173.375 ;
        RECT 51.875 173.085 52.435 173.375 ;
        RECT 52.655 172.915 52.945 173.385 ;
        RECT 53.115 173.085 53.445 173.555 ;
        RECT 53.615 172.915 53.785 173.385 ;
        RECT 53.955 173.085 54.285 173.555 ;
        RECT 54.455 172.915 54.730 173.735 ;
        RECT 54.910 173.445 56.125 173.615 ;
        RECT 54.910 173.095 55.200 173.445 ;
        RECT 55.395 172.915 55.725 173.275 ;
        RECT 55.895 173.140 56.125 173.445 ;
        RECT 56.315 173.220 56.485 173.785 ;
        RECT 58.330 173.460 58.670 174.290 ;
        RECT 60.150 173.780 60.500 175.030 ;
        RECT 62.265 174.375 63.935 175.465 ;
        RECT 62.265 173.685 63.015 174.205 ;
        RECT 63.185 173.855 63.935 174.375 ;
        RECT 64.195 174.535 64.365 175.295 ;
        RECT 64.545 174.705 64.875 175.465 ;
        RECT 64.195 174.365 64.860 174.535 ;
        RECT 65.045 174.390 65.315 175.295 ;
        RECT 64.690 174.220 64.860 174.365 ;
        RECT 64.125 173.815 64.455 174.185 ;
        RECT 64.690 173.890 64.975 174.220 ;
        RECT 56.745 172.915 62.090 173.460 ;
        RECT 62.265 172.915 63.935 173.685 ;
        RECT 64.690 173.635 64.860 173.890 ;
        RECT 64.195 173.465 64.860 173.635 ;
        RECT 65.145 173.590 65.315 174.390 ;
        RECT 65.485 174.375 67.155 175.465 ;
        RECT 64.195 173.085 64.365 173.465 ;
        RECT 64.545 172.915 64.875 173.295 ;
        RECT 65.055 173.085 65.315 173.590 ;
        RECT 65.485 173.685 66.235 174.205 ;
        RECT 66.405 173.855 67.155 174.375 ;
        RECT 67.325 174.615 67.585 175.295 ;
        RECT 67.755 174.685 68.005 175.465 ;
        RECT 68.255 174.915 68.505 175.295 ;
        RECT 68.675 175.085 69.030 175.465 ;
        RECT 70.035 175.075 70.370 175.295 ;
        RECT 69.635 174.915 69.865 174.955 ;
        RECT 68.255 174.715 69.865 174.915 ;
        RECT 68.255 174.705 69.090 174.715 ;
        RECT 69.680 174.625 69.865 174.715 ;
        RECT 65.485 172.915 67.155 173.685 ;
        RECT 67.325 173.415 67.495 174.615 ;
        RECT 69.195 174.515 69.525 174.545 ;
        RECT 67.725 174.455 69.525 174.515 ;
        RECT 70.115 174.455 70.370 175.075 ;
        RECT 67.665 174.345 70.370 174.455 ;
        RECT 70.545 174.375 72.215 175.465 ;
        RECT 67.665 174.310 67.865 174.345 ;
        RECT 67.665 173.735 67.835 174.310 ;
        RECT 69.195 174.285 70.370 174.345 ;
        RECT 68.065 173.870 68.475 174.175 ;
        RECT 68.645 173.905 68.975 174.115 ;
        RECT 67.665 173.615 67.935 173.735 ;
        RECT 67.665 173.570 68.510 173.615 ;
        RECT 67.755 173.445 68.510 173.570 ;
        RECT 68.765 173.505 68.975 173.905 ;
        RECT 69.220 173.905 69.695 174.115 ;
        RECT 69.885 173.905 70.375 174.105 ;
        RECT 69.220 173.505 69.440 173.905 ;
        RECT 70.545 173.685 71.295 174.205 ;
        RECT 71.465 173.855 72.215 174.375 ;
        RECT 72.395 174.515 72.670 175.285 ;
        RECT 72.840 174.855 73.170 175.285 ;
        RECT 73.340 175.025 73.535 175.465 ;
        RECT 73.715 174.855 74.045 175.285 ;
        RECT 72.840 174.685 74.045 174.855 ;
        RECT 72.395 174.325 72.980 174.515 ;
        RECT 73.150 174.355 74.045 174.685 ;
        RECT 74.225 174.375 75.435 175.465 ;
        RECT 67.325 173.085 67.585 173.415 ;
        RECT 68.340 173.295 68.510 173.445 ;
        RECT 67.755 172.915 68.085 173.275 ;
        RECT 68.340 173.085 69.640 173.295 ;
        RECT 69.915 172.915 70.370 173.680 ;
        RECT 70.545 172.915 72.215 173.685 ;
        RECT 72.395 173.505 72.635 174.155 ;
        RECT 72.805 173.655 72.980 174.325 ;
        RECT 73.150 173.825 73.565 174.155 ;
        RECT 73.745 173.825 74.040 174.155 ;
        RECT 72.805 173.475 73.135 173.655 ;
        RECT 72.410 172.915 72.740 173.305 ;
        RECT 72.910 173.095 73.135 173.475 ;
        RECT 73.335 173.205 73.565 173.825 ;
        RECT 74.225 173.665 74.745 174.205 ;
        RECT 74.915 173.835 75.435 174.375 ;
        RECT 75.605 174.300 75.895 175.465 ;
        RECT 76.070 174.325 76.390 175.465 ;
        RECT 76.570 174.155 76.765 175.205 ;
        RECT 76.945 174.615 77.275 175.295 ;
        RECT 77.475 174.665 77.730 175.465 ;
        RECT 76.945 174.335 77.295 174.615 ;
        RECT 76.130 174.105 76.390 174.155 ;
        RECT 76.125 173.935 76.390 174.105 ;
        RECT 76.130 173.825 76.390 173.935 ;
        RECT 76.570 173.825 76.955 174.155 ;
        RECT 77.125 173.955 77.295 174.335 ;
        RECT 77.485 174.125 77.730 174.485 ;
        RECT 77.905 174.375 81.415 175.465 ;
        RECT 77.125 173.785 77.645 173.955 ;
        RECT 77.475 173.765 77.645 173.785 ;
        RECT 73.745 172.915 74.045 173.645 ;
        RECT 74.225 172.915 75.435 173.665 ;
        RECT 75.605 172.915 75.895 173.640 ;
        RECT 76.070 173.445 77.285 173.615 ;
        RECT 76.070 173.095 76.360 173.445 ;
        RECT 76.555 172.915 76.885 173.275 ;
        RECT 77.055 173.140 77.285 173.445 ;
        RECT 77.475 173.595 77.675 173.765 ;
        RECT 77.905 173.685 79.555 174.205 ;
        RECT 79.725 173.855 81.415 174.375 ;
        RECT 82.505 174.325 82.890 175.295 ;
        RECT 83.060 175.005 83.385 175.465 ;
        RECT 83.905 174.835 84.185 175.295 ;
        RECT 83.060 174.615 84.185 174.835 ;
        RECT 77.475 173.220 77.645 173.595 ;
        RECT 77.905 172.915 81.415 173.685 ;
        RECT 82.505 173.655 82.785 174.325 ;
        RECT 83.060 174.155 83.510 174.615 ;
        RECT 84.375 174.445 84.775 175.295 ;
        RECT 85.175 175.005 85.445 175.465 ;
        RECT 85.615 174.835 85.900 175.295 ;
        RECT 82.955 173.825 83.510 174.155 ;
        RECT 83.680 173.885 84.775 174.445 ;
        RECT 83.060 173.715 83.510 173.825 ;
        RECT 82.505 173.085 82.890 173.655 ;
        RECT 83.060 173.545 84.185 173.715 ;
        RECT 83.060 172.915 83.385 173.375 ;
        RECT 83.905 173.085 84.185 173.545 ;
        RECT 84.375 173.085 84.775 173.885 ;
        RECT 84.945 174.615 85.900 174.835 ;
        RECT 84.945 173.715 85.155 174.615 ;
        RECT 85.325 173.885 86.015 174.445 ;
        RECT 86.185 174.375 89.695 175.465 ;
        RECT 84.945 173.545 85.900 173.715 ;
        RECT 85.175 172.915 85.445 173.375 ;
        RECT 85.615 173.085 85.900 173.545 ;
        RECT 86.185 173.685 87.835 174.205 ;
        RECT 88.005 173.855 89.695 174.375 ;
        RECT 89.870 174.325 90.205 175.295 ;
        RECT 90.375 174.325 90.545 175.465 ;
        RECT 90.715 175.125 92.745 175.295 ;
        RECT 86.185 172.915 89.695 173.685 ;
        RECT 89.870 173.655 90.040 174.325 ;
        RECT 90.715 174.155 90.885 175.125 ;
        RECT 90.210 173.825 90.465 174.155 ;
        RECT 90.690 173.825 90.885 174.155 ;
        RECT 91.055 174.785 92.180 174.955 ;
        RECT 90.295 173.655 90.465 173.825 ;
        RECT 91.055 173.655 91.225 174.785 ;
        RECT 89.870 173.085 90.125 173.655 ;
        RECT 90.295 173.485 91.225 173.655 ;
        RECT 91.395 174.445 92.405 174.615 ;
        RECT 91.395 173.645 91.565 174.445 ;
        RECT 91.050 173.450 91.225 173.485 ;
        RECT 90.295 172.915 90.625 173.315 ;
        RECT 91.050 173.085 91.580 173.450 ;
        RECT 91.770 173.425 92.045 174.245 ;
        RECT 91.765 173.255 92.045 173.425 ;
        RECT 91.770 173.085 92.045 173.255 ;
        RECT 92.215 173.085 92.405 174.445 ;
        RECT 92.575 174.460 92.745 175.125 ;
        RECT 92.915 174.705 93.085 175.465 ;
        RECT 93.320 174.705 93.835 175.115 ;
        RECT 92.575 174.270 93.325 174.460 ;
        RECT 93.495 173.895 93.835 174.705 ;
        RECT 94.005 174.375 97.515 175.465 ;
        RECT 98.200 174.595 98.485 175.465 ;
        RECT 98.655 174.835 98.915 175.295 ;
        RECT 99.090 175.005 99.345 175.465 ;
        RECT 99.515 174.835 99.775 175.295 ;
        RECT 98.655 174.665 99.775 174.835 ;
        RECT 99.945 174.665 100.255 175.465 ;
        RECT 98.655 174.415 98.915 174.665 ;
        RECT 100.425 174.495 100.735 175.295 ;
        RECT 92.605 173.725 93.835 173.895 ;
        RECT 92.585 172.915 93.095 173.450 ;
        RECT 93.315 173.120 93.560 173.725 ;
        RECT 94.005 173.685 95.655 174.205 ;
        RECT 95.825 173.855 97.515 174.375 ;
        RECT 98.160 174.245 98.915 174.415 ;
        RECT 99.705 174.325 100.735 174.495 ;
        RECT 98.160 173.735 98.565 174.245 ;
        RECT 99.705 174.075 99.875 174.325 ;
        RECT 98.735 173.905 99.875 174.075 ;
        RECT 94.005 172.915 97.515 173.685 ;
        RECT 98.160 173.565 99.810 173.735 ;
        RECT 100.045 173.585 100.395 174.155 ;
        RECT 98.205 172.915 98.485 173.395 ;
        RECT 98.655 173.175 98.915 173.565 ;
        RECT 99.090 172.915 99.345 173.395 ;
        RECT 99.515 173.175 99.810 173.565 ;
        RECT 100.565 173.415 100.735 174.325 ;
        RECT 101.365 174.300 101.655 175.465 ;
        RECT 101.865 174.325 102.095 175.465 ;
        RECT 102.265 174.315 102.595 175.295 ;
        RECT 102.765 174.325 102.975 175.465 ;
        RECT 103.205 175.030 108.550 175.465 ;
        RECT 101.845 173.905 102.175 174.155 ;
        RECT 99.990 172.915 100.265 173.395 ;
        RECT 100.435 173.085 100.735 173.415 ;
        RECT 101.365 172.915 101.655 173.640 ;
        RECT 101.865 172.915 102.095 173.735 ;
        RECT 102.345 173.715 102.595 174.315 ;
        RECT 102.265 173.085 102.595 173.715 ;
        RECT 102.765 172.915 102.975 173.735 ;
        RECT 104.790 173.460 105.130 174.290 ;
        RECT 106.610 173.780 106.960 175.030 ;
        RECT 109.195 174.405 109.525 175.255 ;
        RECT 109.195 173.640 109.385 174.405 ;
        RECT 109.695 174.325 109.945 175.465 ;
        RECT 110.135 174.825 110.385 175.245 ;
        RECT 110.615 174.995 110.945 175.465 ;
        RECT 111.175 174.825 111.425 175.245 ;
        RECT 110.135 174.655 111.425 174.825 ;
        RECT 111.605 174.825 111.935 175.255 ;
        RECT 111.605 174.655 112.060 174.825 ;
        RECT 112.410 174.665 112.665 175.465 ;
        RECT 110.125 174.155 110.340 174.485 ;
        RECT 109.555 173.825 109.865 174.155 ;
        RECT 110.035 173.825 110.340 174.155 ;
        RECT 110.515 173.825 110.800 174.485 ;
        RECT 110.995 173.825 111.260 174.485 ;
        RECT 111.475 173.825 111.720 174.485 ;
        RECT 109.695 173.655 109.865 173.825 ;
        RECT 111.890 173.655 112.060 174.655 ;
        RECT 112.865 174.615 113.195 175.295 ;
        RECT 112.410 174.125 112.655 174.485 ;
        RECT 112.845 174.335 113.195 174.615 ;
        RECT 112.845 173.955 113.015 174.335 ;
        RECT 113.375 174.155 113.570 175.205 ;
        RECT 113.750 174.325 114.070 175.465 ;
        RECT 114.245 174.375 115.455 175.465 ;
        RECT 103.205 172.915 108.550 173.460 ;
        RECT 109.195 173.130 109.525 173.640 ;
        RECT 109.695 173.485 112.060 173.655 ;
        RECT 112.495 173.785 113.015 173.955 ;
        RECT 113.185 173.825 113.570 174.155 ;
        RECT 113.750 174.105 114.010 174.155 ;
        RECT 113.750 173.935 114.015 174.105 ;
        RECT 113.750 173.825 114.010 173.935 ;
        RECT 109.695 172.915 110.025 173.315 ;
        RECT 111.075 173.145 111.405 173.485 ;
        RECT 111.575 172.915 111.905 173.315 ;
        RECT 112.495 173.220 112.665 173.785 ;
        RECT 114.245 173.665 114.765 174.205 ;
        RECT 114.935 173.835 115.455 174.375 ;
        RECT 115.625 174.745 116.085 175.295 ;
        RECT 116.275 174.745 116.605 175.465 ;
        RECT 112.855 173.445 114.070 173.615 ;
        RECT 112.855 173.140 113.085 173.445 ;
        RECT 113.255 172.915 113.585 173.275 ;
        RECT 113.780 173.095 114.070 173.445 ;
        RECT 114.245 172.915 115.455 173.665 ;
        RECT 115.625 173.375 115.875 174.745 ;
        RECT 116.805 174.575 117.105 175.125 ;
        RECT 117.275 174.795 117.555 175.465 ;
        RECT 116.165 174.405 117.105 174.575 ;
        RECT 116.165 174.155 116.335 174.405 ;
        RECT 117.475 174.155 117.740 174.515 ;
        RECT 118.850 174.325 119.170 175.465 ;
        RECT 119.350 174.155 119.545 175.205 ;
        RECT 119.725 174.615 120.055 175.295 ;
        RECT 120.255 174.665 120.510 175.465 ;
        RECT 120.690 175.075 121.025 175.295 ;
        RECT 122.030 175.085 122.385 175.465 ;
        RECT 119.725 174.335 120.075 174.615 ;
        RECT 116.045 173.825 116.335 174.155 ;
        RECT 116.505 173.905 116.845 174.155 ;
        RECT 117.065 173.905 117.740 174.155 ;
        RECT 118.910 174.105 119.170 174.155 ;
        RECT 118.905 173.935 119.170 174.105 ;
        RECT 118.910 173.825 119.170 173.935 ;
        RECT 119.350 173.825 119.735 174.155 ;
        RECT 119.905 173.955 120.075 174.335 ;
        RECT 120.265 174.125 120.510 174.485 ;
        RECT 120.690 174.455 120.945 175.075 ;
        RECT 121.195 174.915 121.425 174.955 ;
        RECT 122.555 174.915 122.805 175.295 ;
        RECT 121.195 174.715 122.805 174.915 ;
        RECT 121.195 174.625 121.380 174.715 ;
        RECT 121.970 174.705 122.805 174.715 ;
        RECT 123.055 174.685 123.305 175.465 ;
        RECT 123.475 174.615 123.735 175.295 ;
        RECT 121.535 174.515 121.865 174.545 ;
        RECT 121.535 174.455 123.335 174.515 ;
        RECT 120.690 174.345 123.395 174.455 ;
        RECT 120.690 174.285 121.865 174.345 ;
        RECT 123.195 174.310 123.395 174.345 ;
        RECT 116.165 173.735 116.335 173.825 ;
        RECT 119.905 173.785 120.425 173.955 ;
        RECT 120.685 173.905 121.175 174.105 ;
        RECT 121.365 173.905 121.840 174.115 ;
        RECT 120.255 173.765 120.425 173.785 ;
        RECT 116.165 173.545 117.555 173.735 ;
        RECT 115.625 173.085 116.185 173.375 ;
        RECT 116.355 172.915 116.605 173.375 ;
        RECT 117.225 173.185 117.555 173.545 ;
        RECT 118.850 173.445 120.065 173.615 ;
        RECT 118.850 173.095 119.140 173.445 ;
        RECT 119.335 172.915 119.665 173.275 ;
        RECT 119.835 173.140 120.065 173.445 ;
        RECT 120.255 173.595 120.455 173.765 ;
        RECT 120.255 173.220 120.425 173.595 ;
        RECT 120.690 172.915 121.145 173.680 ;
        RECT 121.620 173.505 121.840 173.905 ;
        RECT 122.085 173.905 122.415 174.115 ;
        RECT 122.085 173.505 122.295 173.905 ;
        RECT 122.585 173.870 122.995 174.175 ;
        RECT 123.225 173.735 123.395 174.310 ;
        RECT 123.125 173.615 123.395 173.735 ;
        RECT 122.550 173.570 123.395 173.615 ;
        RECT 122.550 173.445 123.305 173.570 ;
        RECT 122.550 173.295 122.720 173.445 ;
        RECT 123.565 173.425 123.735 174.615 ;
        RECT 123.905 174.375 126.495 175.465 ;
        RECT 123.505 173.415 123.735 173.425 ;
        RECT 121.420 173.085 122.720 173.295 ;
        RECT 122.975 172.915 123.305 173.275 ;
        RECT 123.475 173.085 123.735 173.415 ;
        RECT 123.905 173.685 125.115 174.205 ;
        RECT 125.285 173.855 126.495 174.375 ;
        RECT 127.125 174.300 127.415 175.465 ;
        RECT 127.585 175.030 132.930 175.465 ;
        RECT 133.105 175.030 138.450 175.465 ;
        RECT 138.625 175.030 143.970 175.465 ;
        RECT 123.905 172.915 126.495 173.685 ;
        RECT 127.125 172.915 127.415 173.640 ;
        RECT 129.170 173.460 129.510 174.290 ;
        RECT 130.990 173.780 131.340 175.030 ;
        RECT 134.690 173.460 135.030 174.290 ;
        RECT 136.510 173.780 136.860 175.030 ;
        RECT 140.210 173.460 140.550 174.290 ;
        RECT 142.030 173.780 142.380 175.030 ;
        RECT 144.145 174.375 147.655 175.465 ;
        RECT 147.825 174.375 149.035 175.465 ;
        RECT 144.145 173.685 145.795 174.205 ;
        RECT 145.965 173.855 147.655 174.375 ;
        RECT 127.585 172.915 132.930 173.460 ;
        RECT 133.105 172.915 138.450 173.460 ;
        RECT 138.625 172.915 143.970 173.460 ;
        RECT 144.145 172.915 147.655 173.685 ;
        RECT 147.825 173.665 148.345 174.205 ;
        RECT 148.515 173.835 149.035 174.375 ;
        RECT 149.205 174.375 150.415 175.465 ;
        RECT 149.205 173.835 149.725 174.375 ;
        RECT 149.895 173.665 150.415 174.205 ;
        RECT 147.825 172.915 149.035 173.665 ;
        RECT 149.205 172.915 150.415 173.665 ;
        RECT 11.120 172.745 150.500 172.915 ;
        RECT 11.205 171.995 12.415 172.745 ;
        RECT 11.205 171.455 11.725 171.995 ;
        RECT 12.585 171.975 14.255 172.745 ;
        RECT 14.975 172.195 15.145 172.485 ;
        RECT 15.315 172.365 15.645 172.745 ;
        RECT 14.975 172.025 15.640 172.195 ;
        RECT 11.895 171.285 12.415 171.825 ;
        RECT 12.585 171.455 13.335 171.975 ;
        RECT 13.505 171.285 14.255 171.805 ;
        RECT 11.205 170.195 12.415 171.285 ;
        RECT 12.585 170.195 14.255 171.285 ;
        RECT 14.890 171.205 15.240 171.855 ;
        RECT 15.410 171.035 15.640 172.025 ;
        RECT 14.975 170.865 15.640 171.035 ;
        RECT 14.975 170.365 15.145 170.865 ;
        RECT 15.315 170.195 15.645 170.695 ;
        RECT 15.815 170.365 16.000 172.485 ;
        RECT 16.255 172.285 16.505 172.745 ;
        RECT 16.675 172.295 17.010 172.465 ;
        RECT 17.205 172.295 17.880 172.465 ;
        RECT 16.675 172.155 16.845 172.295 ;
        RECT 16.170 171.165 16.450 172.115 ;
        RECT 16.620 172.025 16.845 172.155 ;
        RECT 16.620 170.920 16.790 172.025 ;
        RECT 17.015 171.875 17.540 172.095 ;
        RECT 16.960 171.110 17.200 171.705 ;
        RECT 17.370 171.175 17.540 171.875 ;
        RECT 17.710 171.515 17.880 172.295 ;
        RECT 18.200 172.245 18.570 172.745 ;
        RECT 18.750 172.295 19.155 172.465 ;
        RECT 19.325 172.295 20.110 172.465 ;
        RECT 18.750 172.065 18.920 172.295 ;
        RECT 18.090 171.765 18.920 172.065 ;
        RECT 19.305 171.795 19.770 172.125 ;
        RECT 18.090 171.735 18.290 171.765 ;
        RECT 18.410 171.515 18.580 171.585 ;
        RECT 17.710 171.345 18.580 171.515 ;
        RECT 18.070 171.255 18.580 171.345 ;
        RECT 16.620 170.790 16.925 170.920 ;
        RECT 17.370 170.810 17.900 171.175 ;
        RECT 16.240 170.195 16.505 170.655 ;
        RECT 16.675 170.365 16.925 170.790 ;
        RECT 18.070 170.640 18.240 171.255 ;
        RECT 17.135 170.470 18.240 170.640 ;
        RECT 18.410 170.195 18.580 170.995 ;
        RECT 18.750 170.695 18.920 171.765 ;
        RECT 19.090 170.865 19.280 171.585 ;
        RECT 19.450 170.835 19.770 171.795 ;
        RECT 19.940 171.835 20.110 172.295 ;
        RECT 20.385 172.215 20.595 172.745 ;
        RECT 20.855 172.005 21.185 172.530 ;
        RECT 21.355 172.135 21.525 172.745 ;
        RECT 21.695 172.090 22.025 172.525 ;
        RECT 23.165 172.095 23.425 172.575 ;
        RECT 23.595 172.205 23.845 172.745 ;
        RECT 21.695 172.005 22.075 172.090 ;
        RECT 20.985 171.835 21.185 172.005 ;
        RECT 21.850 171.965 22.075 172.005 ;
        RECT 19.940 171.505 20.815 171.835 ;
        RECT 20.985 171.505 21.735 171.835 ;
        RECT 18.750 170.365 19.000 170.695 ;
        RECT 19.940 170.665 20.110 171.505 ;
        RECT 20.985 171.300 21.175 171.505 ;
        RECT 21.905 171.385 22.075 171.965 ;
        RECT 21.860 171.335 22.075 171.385 ;
        RECT 20.280 170.925 21.175 171.300 ;
        RECT 21.685 171.255 22.075 171.335 ;
        RECT 19.225 170.495 20.110 170.665 ;
        RECT 20.290 170.195 20.605 170.695 ;
        RECT 20.835 170.365 21.175 170.925 ;
        RECT 21.345 170.195 21.515 171.205 ;
        RECT 21.685 170.410 22.015 171.255 ;
        RECT 23.165 171.065 23.335 172.095 ;
        RECT 24.015 172.040 24.235 172.525 ;
        RECT 23.505 171.445 23.735 171.840 ;
        RECT 23.905 171.615 24.235 172.040 ;
        RECT 24.405 172.365 25.295 172.535 ;
        RECT 24.405 171.640 24.575 172.365 ;
        RECT 24.745 171.810 25.295 172.195 ;
        RECT 25.465 171.975 28.055 172.745 ;
        RECT 24.405 171.570 25.295 171.640 ;
        RECT 24.400 171.545 25.295 171.570 ;
        RECT 24.390 171.530 25.295 171.545 ;
        RECT 24.385 171.515 25.295 171.530 ;
        RECT 24.375 171.510 25.295 171.515 ;
        RECT 24.370 171.500 25.295 171.510 ;
        RECT 24.365 171.490 25.295 171.500 ;
        RECT 24.355 171.485 25.295 171.490 ;
        RECT 24.345 171.475 25.295 171.485 ;
        RECT 24.335 171.470 25.295 171.475 ;
        RECT 24.335 171.465 24.670 171.470 ;
        RECT 24.320 171.460 24.670 171.465 ;
        RECT 24.305 171.450 24.670 171.460 ;
        RECT 24.280 171.445 24.670 171.450 ;
        RECT 23.505 171.440 24.670 171.445 ;
        RECT 23.505 171.405 24.640 171.440 ;
        RECT 23.505 171.380 24.605 171.405 ;
        RECT 23.505 171.350 24.575 171.380 ;
        RECT 23.505 171.320 24.555 171.350 ;
        RECT 23.505 171.290 24.535 171.320 ;
        RECT 23.505 171.280 24.465 171.290 ;
        RECT 23.505 171.270 24.440 171.280 ;
        RECT 23.505 171.255 24.420 171.270 ;
        RECT 23.505 171.240 24.400 171.255 ;
        RECT 23.610 171.230 24.395 171.240 ;
        RECT 23.610 171.195 24.380 171.230 ;
        RECT 23.165 170.365 23.440 171.065 ;
        RECT 23.610 170.945 24.365 171.195 ;
        RECT 24.535 170.875 24.865 171.120 ;
        RECT 25.035 171.020 25.295 171.470 ;
        RECT 25.465 171.455 26.675 171.975 ;
        RECT 28.225 171.925 28.485 172.745 ;
        RECT 28.655 171.925 28.985 172.345 ;
        RECT 29.165 172.260 29.955 172.525 ;
        RECT 28.735 171.835 28.985 171.925 ;
        RECT 26.845 171.285 28.055 171.805 ;
        RECT 24.680 170.850 24.865 170.875 ;
        RECT 24.680 170.750 25.295 170.850 ;
        RECT 23.610 170.195 23.865 170.740 ;
        RECT 24.035 170.365 24.515 170.705 ;
        RECT 24.690 170.195 25.295 170.750 ;
        RECT 25.465 170.195 28.055 171.285 ;
        RECT 28.225 170.875 28.565 171.755 ;
        RECT 28.735 171.585 29.530 171.835 ;
        RECT 28.225 170.195 28.485 170.705 ;
        RECT 28.735 170.365 28.905 171.585 ;
        RECT 29.700 171.405 29.955 172.260 ;
        RECT 30.125 172.105 30.325 172.525 ;
        RECT 30.515 172.285 30.845 172.745 ;
        RECT 30.125 171.585 30.535 172.105 ;
        RECT 31.015 172.095 31.275 172.575 ;
        RECT 30.705 171.405 30.935 171.835 ;
        RECT 29.145 171.235 30.935 171.405 ;
        RECT 29.145 170.870 29.395 171.235 ;
        RECT 29.565 170.875 29.895 171.065 ;
        RECT 30.115 170.940 30.830 171.235 ;
        RECT 31.105 171.065 31.275 172.095 ;
        RECT 29.565 170.700 29.760 170.875 ;
        RECT 29.145 170.195 29.760 170.700 ;
        RECT 29.930 170.365 30.405 170.705 ;
        RECT 30.575 170.195 30.790 170.740 ;
        RECT 31.000 170.365 31.275 171.065 ;
        RECT 32.375 172.020 32.705 172.530 ;
        RECT 32.875 172.345 33.205 172.745 ;
        RECT 34.255 172.175 34.585 172.515 ;
        RECT 34.755 172.345 35.085 172.745 ;
        RECT 32.375 171.255 32.565 172.020 ;
        RECT 32.875 172.005 35.240 172.175 ;
        RECT 32.875 171.835 33.045 172.005 ;
        RECT 32.735 171.505 33.045 171.835 ;
        RECT 33.215 171.505 33.520 171.835 ;
        RECT 32.375 170.405 32.705 171.255 ;
        RECT 32.875 170.195 33.125 171.335 ;
        RECT 33.305 171.175 33.520 171.505 ;
        RECT 33.695 171.175 33.980 171.835 ;
        RECT 34.175 171.175 34.440 171.835 ;
        RECT 34.655 171.175 34.900 171.835 ;
        RECT 35.070 171.005 35.240 172.005 ;
        RECT 35.585 171.995 36.795 172.745 ;
        RECT 36.965 172.020 37.255 172.745 ;
        RECT 37.425 171.995 38.635 172.745 ;
        RECT 35.585 171.455 36.105 171.995 ;
        RECT 36.275 171.285 36.795 171.825 ;
        RECT 37.425 171.455 37.945 171.995 ;
        RECT 38.805 171.925 39.065 172.745 ;
        RECT 39.235 171.925 39.565 172.345 ;
        RECT 39.745 172.260 40.535 172.525 ;
        RECT 39.315 171.835 39.565 171.925 ;
        RECT 33.315 170.835 34.605 171.005 ;
        RECT 33.315 170.415 33.565 170.835 ;
        RECT 33.795 170.195 34.125 170.665 ;
        RECT 34.355 170.415 34.605 170.835 ;
        RECT 34.785 170.835 35.240 171.005 ;
        RECT 34.785 170.405 35.115 170.835 ;
        RECT 35.585 170.195 36.795 171.285 ;
        RECT 36.965 170.195 37.255 171.360 ;
        RECT 38.115 171.285 38.635 171.825 ;
        RECT 37.425 170.195 38.635 171.285 ;
        RECT 38.805 170.875 39.145 171.755 ;
        RECT 39.315 171.585 40.110 171.835 ;
        RECT 38.805 170.195 39.065 170.705 ;
        RECT 39.315 170.365 39.485 171.585 ;
        RECT 40.280 171.405 40.535 172.260 ;
        RECT 40.705 172.105 40.905 172.525 ;
        RECT 41.095 172.285 41.425 172.745 ;
        RECT 40.705 171.585 41.115 172.105 ;
        RECT 41.595 172.095 41.855 172.575 ;
        RECT 41.285 171.405 41.515 171.835 ;
        RECT 39.725 171.235 41.515 171.405 ;
        RECT 39.725 170.870 39.975 171.235 ;
        RECT 40.145 170.875 40.475 171.065 ;
        RECT 40.695 170.940 41.410 171.235 ;
        RECT 41.685 171.065 41.855 172.095 ;
        RECT 42.040 172.175 42.295 172.525 ;
        RECT 42.465 172.345 42.795 172.745 ;
        RECT 42.965 172.175 43.135 172.525 ;
        RECT 43.305 172.345 43.685 172.745 ;
        RECT 42.040 172.005 43.705 172.175 ;
        RECT 43.875 172.070 44.150 172.415 ;
        RECT 43.535 171.835 43.705 172.005 ;
        RECT 42.025 171.505 42.370 171.835 ;
        RECT 42.540 171.505 43.365 171.835 ;
        RECT 43.535 171.505 43.810 171.835 ;
        RECT 40.145 170.700 40.340 170.875 ;
        RECT 39.725 170.195 40.340 170.700 ;
        RECT 40.510 170.365 40.985 170.705 ;
        RECT 41.155 170.195 41.370 170.740 ;
        RECT 41.580 170.365 41.855 171.065 ;
        RECT 42.045 171.045 42.370 171.335 ;
        RECT 42.540 171.215 42.735 171.505 ;
        RECT 43.535 171.335 43.705 171.505 ;
        RECT 43.980 171.335 44.150 172.070 ;
        RECT 44.330 172.005 44.665 172.745 ;
        RECT 44.835 171.835 45.050 172.530 ;
        RECT 45.240 172.005 45.590 172.530 ;
        RECT 45.760 172.005 46.455 172.575 ;
        RECT 45.385 171.835 45.590 172.005 ;
        RECT 44.350 171.505 44.635 171.835 ;
        RECT 44.835 171.505 45.215 171.835 ;
        RECT 45.385 171.505 45.695 171.835 ;
        RECT 45.865 171.335 46.035 172.005 ;
        RECT 46.625 171.975 48.295 172.745 ;
        RECT 48.630 172.235 48.870 172.745 ;
        RECT 49.050 172.235 49.330 172.565 ;
        RECT 49.560 172.235 49.775 172.745 ;
        RECT 43.045 171.165 43.705 171.335 ;
        RECT 43.045 171.045 43.215 171.165 ;
        RECT 42.045 170.875 43.215 171.045 ;
        RECT 42.025 170.415 43.215 170.705 ;
        RECT 43.385 170.195 43.665 170.995 ;
        RECT 43.875 170.365 44.150 171.335 ;
        RECT 44.325 170.195 44.585 171.335 ;
        RECT 44.755 171.165 46.035 171.335 ;
        RECT 46.215 171.165 46.455 171.835 ;
        RECT 46.625 171.455 47.375 171.975 ;
        RECT 47.545 171.285 48.295 171.805 ;
        RECT 48.525 171.505 48.880 172.065 ;
        RECT 49.050 171.335 49.220 172.235 ;
        RECT 49.390 171.505 49.655 172.065 ;
        RECT 49.945 172.005 50.560 172.575 ;
        RECT 50.765 172.200 56.110 172.745 ;
        RECT 49.905 171.335 50.075 171.835 ;
        RECT 44.755 170.365 45.085 171.165 ;
        RECT 45.255 170.195 45.425 170.995 ;
        RECT 45.625 170.365 45.955 171.165 ;
        RECT 46.155 170.195 46.435 170.995 ;
        RECT 46.625 170.195 48.295 171.285 ;
        RECT 48.650 171.165 50.075 171.335 ;
        RECT 48.650 170.990 49.040 171.165 ;
        RECT 49.525 170.195 49.855 170.995 ;
        RECT 50.245 170.985 50.560 172.005 ;
        RECT 52.350 171.370 52.690 172.200 ;
        RECT 56.285 171.975 57.955 172.745 ;
        RECT 58.140 172.175 58.395 172.525 ;
        RECT 58.565 172.345 58.895 172.745 ;
        RECT 59.065 172.175 59.235 172.525 ;
        RECT 59.405 172.345 59.785 172.745 ;
        RECT 58.140 172.005 59.805 172.175 ;
        RECT 59.975 172.070 60.250 172.415 ;
        RECT 50.025 170.365 50.560 170.985 ;
        RECT 54.170 170.630 54.520 171.880 ;
        RECT 56.285 171.455 57.035 171.975 ;
        RECT 59.635 171.835 59.805 172.005 ;
        RECT 57.205 171.285 57.955 171.805 ;
        RECT 58.125 171.505 58.470 171.835 ;
        RECT 58.640 171.505 59.465 171.835 ;
        RECT 59.635 171.505 59.910 171.835 ;
        RECT 50.765 170.195 56.110 170.630 ;
        RECT 56.285 170.195 57.955 171.285 ;
        RECT 58.145 171.045 58.470 171.335 ;
        RECT 58.640 171.215 58.835 171.505 ;
        RECT 59.635 171.335 59.805 171.505 ;
        RECT 60.080 171.335 60.250 172.070 ;
        RECT 60.425 171.975 62.095 172.745 ;
        RECT 62.725 172.020 63.015 172.745 ;
        RECT 63.275 172.195 63.445 172.485 ;
        RECT 63.615 172.365 63.945 172.745 ;
        RECT 63.275 172.025 63.940 172.195 ;
        RECT 60.425 171.455 61.175 171.975 ;
        RECT 59.145 171.165 59.805 171.335 ;
        RECT 59.145 171.045 59.315 171.165 ;
        RECT 58.145 170.875 59.315 171.045 ;
        RECT 58.125 170.415 59.315 170.705 ;
        RECT 59.485 170.195 59.765 170.995 ;
        RECT 59.975 170.365 60.250 171.335 ;
        RECT 61.345 171.285 62.095 171.805 ;
        RECT 60.425 170.195 62.095 171.285 ;
        RECT 62.725 170.195 63.015 171.360 ;
        RECT 63.190 171.205 63.540 171.855 ;
        RECT 63.710 171.035 63.940 172.025 ;
        RECT 63.275 170.865 63.940 171.035 ;
        RECT 63.275 170.365 63.445 170.865 ;
        RECT 63.615 170.195 63.945 170.695 ;
        RECT 64.115 170.365 64.300 172.485 ;
        RECT 64.555 172.285 64.805 172.745 ;
        RECT 64.975 172.295 65.310 172.465 ;
        RECT 65.505 172.295 66.180 172.465 ;
        RECT 64.975 172.155 65.145 172.295 ;
        RECT 64.470 171.165 64.750 172.115 ;
        RECT 64.920 172.025 65.145 172.155 ;
        RECT 64.920 170.920 65.090 172.025 ;
        RECT 65.315 171.875 65.840 172.095 ;
        RECT 65.260 171.110 65.500 171.705 ;
        RECT 65.670 171.175 65.840 171.875 ;
        RECT 66.010 171.515 66.180 172.295 ;
        RECT 66.500 172.245 66.870 172.745 ;
        RECT 67.050 172.295 67.455 172.465 ;
        RECT 67.625 172.295 68.410 172.465 ;
        RECT 67.050 172.065 67.220 172.295 ;
        RECT 66.390 171.765 67.220 172.065 ;
        RECT 67.605 171.795 68.070 172.125 ;
        RECT 66.390 171.735 66.590 171.765 ;
        RECT 66.710 171.515 66.880 171.585 ;
        RECT 66.010 171.345 66.880 171.515 ;
        RECT 66.370 171.255 66.880 171.345 ;
        RECT 64.920 170.790 65.225 170.920 ;
        RECT 65.670 170.810 66.200 171.175 ;
        RECT 64.540 170.195 64.805 170.655 ;
        RECT 64.975 170.365 65.225 170.790 ;
        RECT 66.370 170.640 66.540 171.255 ;
        RECT 65.435 170.470 66.540 170.640 ;
        RECT 66.710 170.195 66.880 170.995 ;
        RECT 67.050 170.695 67.220 171.765 ;
        RECT 67.390 170.865 67.580 171.585 ;
        RECT 67.750 170.835 68.070 171.795 ;
        RECT 68.240 171.835 68.410 172.295 ;
        RECT 68.685 172.215 68.895 172.745 ;
        RECT 69.155 172.005 69.485 172.530 ;
        RECT 69.655 172.135 69.825 172.745 ;
        RECT 69.995 172.090 70.325 172.525 ;
        RECT 69.995 172.005 70.375 172.090 ;
        RECT 69.285 171.835 69.485 172.005 ;
        RECT 70.150 171.965 70.375 172.005 ;
        RECT 68.240 171.505 69.115 171.835 ;
        RECT 69.285 171.505 70.035 171.835 ;
        RECT 67.050 170.365 67.300 170.695 ;
        RECT 68.240 170.665 68.410 171.505 ;
        RECT 69.285 171.300 69.475 171.505 ;
        RECT 70.205 171.385 70.375 171.965 ;
        RECT 70.545 171.975 72.215 172.745 ;
        RECT 70.545 171.455 71.295 171.975 ;
        RECT 72.905 171.925 73.115 172.745 ;
        RECT 73.285 171.945 73.615 172.575 ;
        RECT 70.160 171.335 70.375 171.385 ;
        RECT 68.580 170.925 69.475 171.300 ;
        RECT 69.985 171.255 70.375 171.335 ;
        RECT 71.465 171.285 72.215 171.805 ;
        RECT 73.285 171.345 73.535 171.945 ;
        RECT 73.785 171.925 74.015 172.745 ;
        RECT 74.240 172.175 74.495 172.525 ;
        RECT 74.665 172.345 74.995 172.745 ;
        RECT 75.165 172.175 75.335 172.525 ;
        RECT 75.505 172.345 75.885 172.745 ;
        RECT 74.240 172.005 75.905 172.175 ;
        RECT 76.075 172.070 76.350 172.415 ;
        RECT 75.735 171.835 75.905 172.005 ;
        RECT 73.705 171.505 74.035 171.755 ;
        RECT 74.225 171.505 74.570 171.835 ;
        RECT 74.740 171.505 75.565 171.835 ;
        RECT 75.735 171.505 76.010 171.835 ;
        RECT 67.525 170.495 68.410 170.665 ;
        RECT 68.590 170.195 68.905 170.695 ;
        RECT 69.135 170.365 69.475 170.925 ;
        RECT 69.645 170.195 69.815 171.205 ;
        RECT 69.985 170.410 70.315 171.255 ;
        RECT 70.545 170.195 72.215 171.285 ;
        RECT 72.905 170.195 73.115 171.335 ;
        RECT 73.285 170.365 73.615 171.345 ;
        RECT 73.785 170.195 74.015 171.335 ;
        RECT 74.245 171.045 74.570 171.335 ;
        RECT 74.740 171.215 74.935 171.505 ;
        RECT 75.735 171.335 75.905 171.505 ;
        RECT 76.180 171.335 76.350 172.070 ;
        RECT 75.245 171.165 75.905 171.335 ;
        RECT 75.245 171.045 75.415 171.165 ;
        RECT 74.245 170.875 75.415 171.045 ;
        RECT 74.225 170.415 75.415 170.705 ;
        RECT 75.585 170.195 75.865 170.995 ;
        RECT 76.075 170.365 76.350 171.335 ;
        RECT 76.525 172.095 76.785 172.575 ;
        RECT 76.955 172.205 77.205 172.745 ;
        RECT 76.525 171.065 76.695 172.095 ;
        RECT 77.375 172.040 77.595 172.525 ;
        RECT 76.865 171.445 77.095 171.840 ;
        RECT 77.265 171.615 77.595 172.040 ;
        RECT 77.765 172.365 78.655 172.535 ;
        RECT 77.765 171.640 77.935 172.365 ;
        RECT 78.915 172.195 79.085 172.485 ;
        RECT 79.255 172.365 79.585 172.745 ;
        RECT 78.105 171.810 78.655 172.195 ;
        RECT 78.915 172.025 79.580 172.195 ;
        RECT 77.765 171.570 78.655 171.640 ;
        RECT 77.760 171.545 78.655 171.570 ;
        RECT 77.750 171.530 78.655 171.545 ;
        RECT 77.745 171.515 78.655 171.530 ;
        RECT 77.735 171.510 78.655 171.515 ;
        RECT 77.730 171.500 78.655 171.510 ;
        RECT 77.725 171.490 78.655 171.500 ;
        RECT 77.715 171.485 78.655 171.490 ;
        RECT 77.705 171.475 78.655 171.485 ;
        RECT 77.695 171.470 78.655 171.475 ;
        RECT 77.695 171.465 78.030 171.470 ;
        RECT 77.680 171.460 78.030 171.465 ;
        RECT 77.665 171.450 78.030 171.460 ;
        RECT 77.640 171.445 78.030 171.450 ;
        RECT 76.865 171.440 78.030 171.445 ;
        RECT 76.865 171.405 78.000 171.440 ;
        RECT 76.865 171.380 77.965 171.405 ;
        RECT 76.865 171.350 77.935 171.380 ;
        RECT 76.865 171.320 77.915 171.350 ;
        RECT 76.865 171.290 77.895 171.320 ;
        RECT 76.865 171.280 77.825 171.290 ;
        RECT 76.865 171.270 77.800 171.280 ;
        RECT 76.865 171.255 77.780 171.270 ;
        RECT 76.865 171.240 77.760 171.255 ;
        RECT 76.970 171.230 77.755 171.240 ;
        RECT 76.970 171.195 77.740 171.230 ;
        RECT 76.525 170.365 76.800 171.065 ;
        RECT 76.970 170.945 77.725 171.195 ;
        RECT 77.895 170.875 78.225 171.120 ;
        RECT 78.395 171.020 78.655 171.470 ;
        RECT 78.830 171.205 79.180 171.855 ;
        RECT 79.350 171.035 79.580 172.025 ;
        RECT 78.040 170.850 78.225 170.875 ;
        RECT 78.915 170.865 79.580 171.035 ;
        RECT 78.040 170.750 78.655 170.850 ;
        RECT 76.970 170.195 77.225 170.740 ;
        RECT 77.395 170.365 77.875 170.705 ;
        RECT 78.050 170.195 78.655 170.750 ;
        RECT 78.915 170.365 79.085 170.865 ;
        RECT 79.255 170.195 79.585 170.695 ;
        RECT 79.755 170.365 79.940 172.485 ;
        RECT 80.195 172.285 80.445 172.745 ;
        RECT 80.615 172.295 80.950 172.465 ;
        RECT 81.145 172.295 81.820 172.465 ;
        RECT 80.615 172.155 80.785 172.295 ;
        RECT 80.110 171.165 80.390 172.115 ;
        RECT 80.560 172.025 80.785 172.155 ;
        RECT 80.560 170.920 80.730 172.025 ;
        RECT 80.955 171.875 81.480 172.095 ;
        RECT 80.900 171.110 81.140 171.705 ;
        RECT 81.310 171.175 81.480 171.875 ;
        RECT 81.650 171.515 81.820 172.295 ;
        RECT 82.140 172.245 82.510 172.745 ;
        RECT 82.690 172.295 83.095 172.465 ;
        RECT 83.265 172.295 84.050 172.465 ;
        RECT 82.690 172.065 82.860 172.295 ;
        RECT 82.030 171.765 82.860 172.065 ;
        RECT 83.245 171.795 83.710 172.125 ;
        RECT 82.030 171.735 82.230 171.765 ;
        RECT 82.350 171.515 82.520 171.585 ;
        RECT 81.650 171.345 82.520 171.515 ;
        RECT 82.010 171.255 82.520 171.345 ;
        RECT 80.560 170.790 80.865 170.920 ;
        RECT 81.310 170.810 81.840 171.175 ;
        RECT 80.180 170.195 80.445 170.655 ;
        RECT 80.615 170.365 80.865 170.790 ;
        RECT 82.010 170.640 82.180 171.255 ;
        RECT 81.075 170.470 82.180 170.640 ;
        RECT 82.350 170.195 82.520 170.995 ;
        RECT 82.690 170.695 82.860 171.765 ;
        RECT 83.030 170.865 83.220 171.585 ;
        RECT 83.390 170.835 83.710 171.795 ;
        RECT 83.880 171.835 84.050 172.295 ;
        RECT 84.325 172.215 84.535 172.745 ;
        RECT 84.795 172.005 85.125 172.530 ;
        RECT 85.295 172.135 85.465 172.745 ;
        RECT 85.635 172.090 85.965 172.525 ;
        RECT 86.135 172.230 86.305 172.745 ;
        RECT 85.635 172.005 86.015 172.090 ;
        RECT 84.925 171.835 85.125 172.005 ;
        RECT 85.790 171.965 86.015 172.005 ;
        RECT 83.880 171.505 84.755 171.835 ;
        RECT 84.925 171.505 85.675 171.835 ;
        RECT 82.690 170.365 82.940 170.695 ;
        RECT 83.880 170.665 84.050 171.505 ;
        RECT 84.925 171.300 85.115 171.505 ;
        RECT 85.845 171.385 86.015 171.965 ;
        RECT 86.645 171.975 88.315 172.745 ;
        RECT 88.485 172.020 88.775 172.745 ;
        RECT 89.430 172.095 89.740 172.565 ;
        RECT 89.910 172.265 90.645 172.745 ;
        RECT 90.815 172.175 90.985 172.525 ;
        RECT 91.155 172.345 91.535 172.745 ;
        RECT 86.645 171.455 87.395 171.975 ;
        RECT 89.430 171.925 90.165 172.095 ;
        RECT 90.815 172.005 91.555 172.175 ;
        RECT 91.725 172.070 91.995 172.415 ;
        RECT 89.915 171.835 90.165 171.925 ;
        RECT 91.385 171.835 91.555 172.005 ;
        RECT 85.800 171.335 86.015 171.385 ;
        RECT 84.220 170.925 85.115 171.300 ;
        RECT 85.625 171.255 86.015 171.335 ;
        RECT 87.565 171.285 88.315 171.805 ;
        RECT 89.410 171.505 89.745 171.755 ;
        RECT 89.915 171.505 90.655 171.835 ;
        RECT 91.385 171.505 91.615 171.835 ;
        RECT 83.165 170.495 84.050 170.665 ;
        RECT 84.230 170.195 84.545 170.695 ;
        RECT 84.775 170.365 85.115 170.925 ;
        RECT 85.285 170.195 85.455 171.205 ;
        RECT 85.625 170.410 85.955 171.255 ;
        RECT 86.125 170.195 86.295 171.110 ;
        RECT 86.645 170.195 88.315 171.285 ;
        RECT 88.485 170.195 88.775 171.360 ;
        RECT 89.410 170.195 89.665 171.335 ;
        RECT 89.915 170.945 90.085 171.505 ;
        RECT 91.385 171.335 91.555 171.505 ;
        RECT 91.825 171.335 91.995 172.070 ;
        RECT 92.190 172.095 92.500 172.565 ;
        RECT 92.670 172.265 93.405 172.745 ;
        RECT 93.575 172.175 93.745 172.525 ;
        RECT 93.915 172.345 94.295 172.745 ;
        RECT 92.190 171.925 92.925 172.095 ;
        RECT 93.575 172.005 94.315 172.175 ;
        RECT 94.485 172.070 94.755 172.415 ;
        RECT 94.925 172.200 100.270 172.745 ;
        RECT 92.675 171.835 92.925 171.925 ;
        RECT 94.145 171.835 94.315 172.005 ;
        RECT 92.170 171.505 92.505 171.755 ;
        RECT 92.675 171.505 93.415 171.835 ;
        RECT 94.145 171.505 94.375 171.835 ;
        RECT 90.310 171.165 91.555 171.335 ;
        RECT 90.310 170.915 90.730 171.165 ;
        RECT 89.860 170.415 91.055 170.745 ;
        RECT 91.235 170.195 91.515 170.995 ;
        RECT 91.725 170.365 91.995 171.335 ;
        RECT 92.170 170.195 92.425 171.335 ;
        RECT 92.675 170.945 92.845 171.505 ;
        RECT 94.145 171.335 94.315 171.505 ;
        RECT 94.585 171.335 94.755 172.070 ;
        RECT 96.510 171.370 96.850 172.200 ;
        RECT 100.445 171.995 101.655 172.745 ;
        RECT 93.070 171.165 94.315 171.335 ;
        RECT 93.070 170.915 93.490 171.165 ;
        RECT 92.620 170.415 93.815 170.745 ;
        RECT 93.995 170.195 94.275 170.995 ;
        RECT 94.485 170.365 94.755 171.335 ;
        RECT 98.330 170.630 98.680 171.880 ;
        RECT 100.445 171.455 100.965 171.995 ;
        RECT 101.885 171.925 102.095 172.745 ;
        RECT 102.265 171.945 102.595 172.575 ;
        RECT 101.135 171.285 101.655 171.825 ;
        RECT 102.265 171.345 102.515 171.945 ;
        RECT 102.765 171.925 102.995 172.745 ;
        RECT 103.205 171.975 105.795 172.745 ;
        RECT 105.965 172.005 106.350 172.575 ;
        RECT 106.520 172.285 106.845 172.745 ;
        RECT 107.365 172.115 107.645 172.575 ;
        RECT 102.685 171.505 103.015 171.755 ;
        RECT 103.205 171.455 104.415 171.975 ;
        RECT 94.925 170.195 100.270 170.630 ;
        RECT 100.445 170.195 101.655 171.285 ;
        RECT 101.885 170.195 102.095 171.335 ;
        RECT 102.265 170.365 102.595 171.345 ;
        RECT 102.765 170.195 102.995 171.335 ;
        RECT 104.585 171.285 105.795 171.805 ;
        RECT 103.205 170.195 105.795 171.285 ;
        RECT 105.965 171.335 106.245 172.005 ;
        RECT 106.520 171.945 107.645 172.115 ;
        RECT 106.520 171.835 106.970 171.945 ;
        RECT 106.415 171.505 106.970 171.835 ;
        RECT 107.835 171.775 108.235 172.575 ;
        RECT 108.635 172.285 108.905 172.745 ;
        RECT 109.075 172.115 109.360 172.575 ;
        RECT 105.965 170.365 106.350 171.335 ;
        RECT 106.520 171.045 106.970 171.505 ;
        RECT 107.140 171.215 108.235 171.775 ;
        RECT 106.520 170.825 107.645 171.045 ;
        RECT 106.520 170.195 106.845 170.655 ;
        RECT 107.365 170.365 107.645 170.825 ;
        RECT 107.835 170.365 108.235 171.215 ;
        RECT 108.405 171.945 109.360 172.115 ;
        RECT 109.645 171.975 111.315 172.745 ;
        RECT 111.980 172.005 112.595 172.575 ;
        RECT 112.765 172.235 112.980 172.745 ;
        RECT 113.210 172.235 113.490 172.565 ;
        RECT 113.670 172.235 113.910 172.745 ;
        RECT 108.405 171.045 108.615 171.945 ;
        RECT 108.785 171.215 109.475 171.775 ;
        RECT 109.645 171.455 110.395 171.975 ;
        RECT 110.565 171.285 111.315 171.805 ;
        RECT 108.405 170.825 109.360 171.045 ;
        RECT 108.635 170.195 108.905 170.655 ;
        RECT 109.075 170.365 109.360 170.825 ;
        RECT 109.645 170.195 111.315 171.285 ;
        RECT 111.980 170.985 112.295 172.005 ;
        RECT 112.465 171.335 112.635 171.835 ;
        RECT 112.885 171.505 113.150 172.065 ;
        RECT 113.320 171.335 113.490 172.235 ;
        RECT 113.660 171.505 114.015 172.065 ;
        RECT 114.245 172.020 114.535 172.745 ;
        RECT 114.730 172.355 115.060 172.745 ;
        RECT 115.230 172.185 115.455 172.565 ;
        RECT 114.715 171.505 114.955 172.155 ;
        RECT 115.125 172.005 115.455 172.185 ;
        RECT 112.465 171.165 113.890 171.335 ;
        RECT 111.980 170.365 112.515 170.985 ;
        RECT 112.685 170.195 113.015 170.995 ;
        RECT 113.500 170.990 113.890 171.165 ;
        RECT 114.245 170.195 114.535 171.360 ;
        RECT 115.125 171.335 115.300 172.005 ;
        RECT 115.655 171.835 115.885 172.455 ;
        RECT 116.065 172.015 116.365 172.745 ;
        RECT 117.170 172.235 117.410 172.745 ;
        RECT 117.590 172.235 117.870 172.565 ;
        RECT 118.100 172.235 118.315 172.745 ;
        RECT 115.470 171.505 115.885 171.835 ;
        RECT 116.065 171.505 116.360 171.835 ;
        RECT 117.065 171.505 117.420 172.065 ;
        RECT 117.590 171.335 117.760 172.235 ;
        RECT 117.930 171.505 118.195 172.065 ;
        RECT 118.485 172.005 119.100 172.575 ;
        RECT 118.445 171.335 118.615 171.835 ;
        RECT 114.715 171.145 115.300 171.335 ;
        RECT 114.715 170.375 114.990 171.145 ;
        RECT 115.470 170.975 116.365 171.305 ;
        RECT 117.190 171.165 118.615 171.335 ;
        RECT 117.190 170.990 117.580 171.165 ;
        RECT 115.160 170.805 116.365 170.975 ;
        RECT 115.160 170.375 115.490 170.805 ;
        RECT 115.660 170.195 115.855 170.635 ;
        RECT 116.035 170.375 116.365 170.805 ;
        RECT 118.065 170.195 118.395 170.995 ;
        RECT 118.785 170.985 119.100 172.005 ;
        RECT 119.305 171.975 122.815 172.745 ;
        RECT 123.075 172.195 123.245 172.485 ;
        RECT 123.415 172.365 123.745 172.745 ;
        RECT 123.075 172.025 123.740 172.195 ;
        RECT 119.305 171.455 120.955 171.975 ;
        RECT 121.125 171.285 122.815 171.805 ;
        RECT 118.565 170.365 119.100 170.985 ;
        RECT 119.305 170.195 122.815 171.285 ;
        RECT 122.990 171.205 123.340 171.855 ;
        RECT 123.510 171.035 123.740 172.025 ;
        RECT 123.075 170.865 123.740 171.035 ;
        RECT 123.075 170.365 123.245 170.865 ;
        RECT 123.415 170.195 123.745 170.695 ;
        RECT 123.915 170.365 124.100 172.485 ;
        RECT 124.355 172.285 124.605 172.745 ;
        RECT 124.775 172.295 125.110 172.465 ;
        RECT 125.305 172.295 125.980 172.465 ;
        RECT 124.775 172.155 124.945 172.295 ;
        RECT 124.270 171.165 124.550 172.115 ;
        RECT 124.720 172.025 124.945 172.155 ;
        RECT 124.720 170.920 124.890 172.025 ;
        RECT 125.115 171.875 125.640 172.095 ;
        RECT 125.060 171.110 125.300 171.705 ;
        RECT 125.470 171.175 125.640 171.875 ;
        RECT 125.810 171.515 125.980 172.295 ;
        RECT 126.300 172.245 126.670 172.745 ;
        RECT 126.850 172.295 127.255 172.465 ;
        RECT 127.425 172.295 128.210 172.465 ;
        RECT 126.850 172.065 127.020 172.295 ;
        RECT 126.190 171.765 127.020 172.065 ;
        RECT 127.405 171.795 127.870 172.125 ;
        RECT 126.190 171.735 126.390 171.765 ;
        RECT 126.510 171.515 126.680 171.585 ;
        RECT 125.810 171.345 126.680 171.515 ;
        RECT 126.170 171.255 126.680 171.345 ;
        RECT 124.720 170.790 125.025 170.920 ;
        RECT 125.470 170.810 126.000 171.175 ;
        RECT 124.340 170.195 124.605 170.655 ;
        RECT 124.775 170.365 125.025 170.790 ;
        RECT 126.170 170.640 126.340 171.255 ;
        RECT 125.235 170.470 126.340 170.640 ;
        RECT 126.510 170.195 126.680 170.995 ;
        RECT 126.850 170.695 127.020 171.765 ;
        RECT 127.190 170.865 127.380 171.585 ;
        RECT 127.550 170.835 127.870 171.795 ;
        RECT 128.040 171.835 128.210 172.295 ;
        RECT 128.485 172.215 128.695 172.745 ;
        RECT 128.955 172.005 129.285 172.530 ;
        RECT 129.455 172.135 129.625 172.745 ;
        RECT 129.795 172.090 130.125 172.525 ;
        RECT 130.295 172.230 130.465 172.745 ;
        RECT 130.805 172.200 136.150 172.745 ;
        RECT 129.795 172.005 130.175 172.090 ;
        RECT 129.085 171.835 129.285 172.005 ;
        RECT 129.950 171.965 130.175 172.005 ;
        RECT 128.040 171.505 128.915 171.835 ;
        RECT 129.085 171.505 129.835 171.835 ;
        RECT 126.850 170.365 127.100 170.695 ;
        RECT 128.040 170.665 128.210 171.505 ;
        RECT 129.085 171.300 129.275 171.505 ;
        RECT 130.005 171.385 130.175 171.965 ;
        RECT 129.960 171.335 130.175 171.385 ;
        RECT 132.390 171.370 132.730 172.200 ;
        RECT 136.325 171.975 139.835 172.745 ;
        RECT 140.005 172.020 140.295 172.745 ;
        RECT 140.465 172.200 145.810 172.745 ;
        RECT 128.380 170.925 129.275 171.300 ;
        RECT 129.785 171.255 130.175 171.335 ;
        RECT 127.325 170.495 128.210 170.665 ;
        RECT 128.390 170.195 128.705 170.695 ;
        RECT 128.935 170.365 129.275 170.925 ;
        RECT 129.445 170.195 129.615 171.205 ;
        RECT 129.785 170.410 130.115 171.255 ;
        RECT 130.285 170.195 130.455 171.110 ;
        RECT 134.210 170.630 134.560 171.880 ;
        RECT 136.325 171.455 137.975 171.975 ;
        RECT 138.145 171.285 139.835 171.805 ;
        RECT 142.050 171.370 142.390 172.200 ;
        RECT 145.985 171.975 148.575 172.745 ;
        RECT 149.205 171.995 150.415 172.745 ;
        RECT 130.805 170.195 136.150 170.630 ;
        RECT 136.325 170.195 139.835 171.285 ;
        RECT 140.005 170.195 140.295 171.360 ;
        RECT 143.870 170.630 144.220 171.880 ;
        RECT 145.985 171.455 147.195 171.975 ;
        RECT 147.365 171.285 148.575 171.805 ;
        RECT 140.465 170.195 145.810 170.630 ;
        RECT 145.985 170.195 148.575 171.285 ;
        RECT 149.205 171.285 149.725 171.825 ;
        RECT 149.895 171.455 150.415 171.995 ;
        RECT 149.205 170.195 150.415 171.285 ;
        RECT 11.120 170.025 150.500 170.195 ;
        RECT 11.205 168.935 12.415 170.025 ;
        RECT 12.585 168.935 15.175 170.025 ;
        RECT 15.345 169.515 15.605 170.025 ;
        RECT 11.205 168.225 11.725 168.765 ;
        RECT 11.895 168.395 12.415 168.935 ;
        RECT 12.585 168.245 13.795 168.765 ;
        RECT 13.965 168.415 15.175 168.935 ;
        RECT 15.345 168.465 15.685 169.345 ;
        RECT 15.855 168.635 16.025 169.855 ;
        RECT 16.265 169.520 16.880 170.025 ;
        RECT 16.265 168.985 16.515 169.350 ;
        RECT 16.685 169.345 16.880 169.520 ;
        RECT 17.050 169.515 17.525 169.855 ;
        RECT 17.695 169.480 17.910 170.025 ;
        RECT 16.685 169.155 17.015 169.345 ;
        RECT 17.235 168.985 17.950 169.280 ;
        RECT 18.120 169.155 18.395 169.855 ;
        RECT 16.265 168.815 18.055 168.985 ;
        RECT 15.855 168.385 16.650 168.635 ;
        RECT 15.855 168.295 16.105 168.385 ;
        RECT 11.205 167.475 12.415 168.225 ;
        RECT 12.585 167.475 15.175 168.245 ;
        RECT 15.345 167.475 15.605 168.295 ;
        RECT 15.775 167.875 16.105 168.295 ;
        RECT 16.820 167.960 17.075 168.815 ;
        RECT 16.285 167.695 17.075 167.960 ;
        RECT 17.245 168.115 17.655 168.635 ;
        RECT 17.825 168.385 18.055 168.815 ;
        RECT 18.225 168.125 18.395 169.155 ;
        RECT 18.565 168.935 20.235 170.025 ;
        RECT 17.245 167.695 17.445 168.115 ;
        RECT 17.635 167.475 17.965 167.935 ;
        RECT 18.135 167.645 18.395 168.125 ;
        RECT 18.565 168.245 19.315 168.765 ;
        RECT 19.485 168.415 20.235 168.935 ;
        RECT 20.415 169.055 20.745 169.840 ;
        RECT 20.415 168.885 21.095 169.055 ;
        RECT 21.275 168.885 21.605 170.025 ;
        RECT 21.820 169.235 22.355 169.855 ;
        RECT 20.405 168.465 20.755 168.715 ;
        RECT 20.925 168.285 21.095 168.885 ;
        RECT 21.265 168.465 21.615 168.715 ;
        RECT 18.565 167.475 20.235 168.245 ;
        RECT 20.425 167.475 20.665 168.285 ;
        RECT 20.835 167.645 21.165 168.285 ;
        RECT 21.335 167.475 21.605 168.285 ;
        RECT 21.820 168.215 22.135 169.235 ;
        RECT 22.525 169.225 22.855 170.025 ;
        RECT 23.340 169.055 23.730 169.230 ;
        RECT 22.305 168.885 23.730 169.055 ;
        RECT 22.305 168.385 22.475 168.885 ;
        RECT 21.820 167.645 22.435 168.215 ;
        RECT 22.725 168.155 22.990 168.715 ;
        RECT 23.160 167.985 23.330 168.885 ;
        RECT 24.085 168.860 24.375 170.025 ;
        RECT 24.545 169.305 25.005 169.855 ;
        RECT 25.195 169.305 25.525 170.025 ;
        RECT 23.500 168.155 23.855 168.715 ;
        RECT 22.605 167.475 22.820 167.985 ;
        RECT 23.050 167.655 23.330 167.985 ;
        RECT 23.510 167.475 23.750 167.985 ;
        RECT 24.085 167.475 24.375 168.200 ;
        RECT 24.545 167.935 24.795 169.305 ;
        RECT 25.725 169.135 26.025 169.685 ;
        RECT 26.195 169.355 26.475 170.025 ;
        RECT 26.850 169.225 27.105 170.025 ;
        RECT 27.305 169.175 27.635 169.855 ;
        RECT 25.085 168.965 26.025 169.135 ;
        RECT 25.085 168.715 25.255 168.965 ;
        RECT 26.395 168.715 26.660 169.075 ;
        RECT 24.965 168.385 25.255 168.715 ;
        RECT 25.425 168.465 25.765 168.715 ;
        RECT 25.985 168.465 26.660 168.715 ;
        RECT 26.850 168.685 27.095 169.045 ;
        RECT 27.285 168.895 27.635 169.175 ;
        RECT 27.285 168.515 27.455 168.895 ;
        RECT 27.815 168.715 28.010 169.765 ;
        RECT 28.190 168.885 28.510 170.025 ;
        RECT 29.235 169.355 29.405 169.855 ;
        RECT 29.575 169.525 29.905 170.025 ;
        RECT 29.235 169.185 29.900 169.355 ;
        RECT 25.085 168.295 25.255 168.385 ;
        RECT 26.935 168.345 27.455 168.515 ;
        RECT 27.625 168.385 28.010 168.715 ;
        RECT 28.190 168.665 28.450 168.715 ;
        RECT 28.190 168.495 28.455 168.665 ;
        RECT 28.190 168.385 28.450 168.495 ;
        RECT 29.150 168.365 29.500 169.015 ;
        RECT 26.935 168.325 27.105 168.345 ;
        RECT 25.085 168.105 26.475 168.295 ;
        RECT 26.905 168.155 27.105 168.325 ;
        RECT 29.670 168.195 29.900 169.185 ;
        RECT 24.545 167.645 25.105 167.935 ;
        RECT 25.275 167.475 25.525 167.935 ;
        RECT 26.145 167.745 26.475 168.105 ;
        RECT 26.935 167.780 27.105 168.155 ;
        RECT 27.295 168.005 28.510 168.175 ;
        RECT 27.295 167.700 27.525 168.005 ;
        RECT 27.695 167.475 28.025 167.835 ;
        RECT 28.220 167.655 28.510 168.005 ;
        RECT 29.235 168.025 29.900 168.195 ;
        RECT 29.235 167.735 29.405 168.025 ;
        RECT 29.575 167.475 29.905 167.855 ;
        RECT 30.075 167.735 30.260 169.855 ;
        RECT 30.500 169.565 30.765 170.025 ;
        RECT 30.935 169.430 31.185 169.855 ;
        RECT 31.395 169.580 32.500 169.750 ;
        RECT 30.880 169.300 31.185 169.430 ;
        RECT 30.430 168.105 30.710 169.055 ;
        RECT 30.880 168.195 31.050 169.300 ;
        RECT 31.220 168.515 31.460 169.110 ;
        RECT 31.630 169.045 32.160 169.410 ;
        RECT 31.630 168.345 31.800 169.045 ;
        RECT 32.330 168.965 32.500 169.580 ;
        RECT 32.670 169.225 32.840 170.025 ;
        RECT 33.010 169.525 33.260 169.855 ;
        RECT 33.485 169.555 34.370 169.725 ;
        RECT 32.330 168.875 32.840 168.965 ;
        RECT 30.880 168.065 31.105 168.195 ;
        RECT 31.275 168.125 31.800 168.345 ;
        RECT 31.970 168.705 32.840 168.875 ;
        RECT 30.515 167.475 30.765 167.935 ;
        RECT 30.935 167.925 31.105 168.065 ;
        RECT 31.970 167.925 32.140 168.705 ;
        RECT 32.670 168.635 32.840 168.705 ;
        RECT 32.350 168.455 32.550 168.485 ;
        RECT 33.010 168.455 33.180 169.525 ;
        RECT 33.350 168.635 33.540 169.355 ;
        RECT 32.350 168.155 33.180 168.455 ;
        RECT 33.710 168.425 34.030 169.385 ;
        RECT 30.935 167.755 31.270 167.925 ;
        RECT 31.465 167.755 32.140 167.925 ;
        RECT 32.460 167.475 32.830 167.975 ;
        RECT 33.010 167.925 33.180 168.155 ;
        RECT 33.565 168.095 34.030 168.425 ;
        RECT 34.200 168.715 34.370 169.555 ;
        RECT 34.550 169.525 34.865 170.025 ;
        RECT 35.095 169.295 35.435 169.855 ;
        RECT 34.540 168.920 35.435 169.295 ;
        RECT 35.605 169.015 35.775 170.025 ;
        RECT 35.245 168.715 35.435 168.920 ;
        RECT 35.945 168.965 36.275 169.810 ;
        RECT 35.945 168.885 36.335 168.965 ;
        RECT 36.505 168.935 37.715 170.025 ;
        RECT 36.120 168.835 36.335 168.885 ;
        RECT 34.200 168.385 35.075 168.715 ;
        RECT 35.245 168.385 35.995 168.715 ;
        RECT 34.200 167.925 34.370 168.385 ;
        RECT 35.245 168.215 35.445 168.385 ;
        RECT 36.165 168.255 36.335 168.835 ;
        RECT 36.110 168.215 36.335 168.255 ;
        RECT 33.010 167.755 33.415 167.925 ;
        RECT 33.585 167.755 34.370 167.925 ;
        RECT 34.645 167.475 34.855 168.005 ;
        RECT 35.115 167.690 35.445 168.215 ;
        RECT 35.955 168.130 36.335 168.215 ;
        RECT 36.505 168.225 37.025 168.765 ;
        RECT 37.195 168.395 37.715 168.935 ;
        RECT 37.885 169.155 38.160 169.855 ;
        RECT 38.330 169.480 38.585 170.025 ;
        RECT 38.755 169.515 39.235 169.855 ;
        RECT 39.410 169.470 40.015 170.025 ;
        RECT 39.400 169.370 40.015 169.470 ;
        RECT 39.400 169.345 39.585 169.370 ;
        RECT 35.615 167.475 35.785 168.085 ;
        RECT 35.955 167.695 36.285 168.130 ;
        RECT 36.505 167.475 37.715 168.225 ;
        RECT 37.885 168.125 38.055 169.155 ;
        RECT 38.330 169.025 39.085 169.275 ;
        RECT 39.255 169.100 39.585 169.345 ;
        RECT 38.330 168.990 39.100 169.025 ;
        RECT 38.330 168.980 39.115 168.990 ;
        RECT 38.225 168.965 39.120 168.980 ;
        RECT 38.225 168.950 39.140 168.965 ;
        RECT 38.225 168.940 39.160 168.950 ;
        RECT 38.225 168.930 39.185 168.940 ;
        RECT 38.225 168.900 39.255 168.930 ;
        RECT 38.225 168.870 39.275 168.900 ;
        RECT 38.225 168.840 39.295 168.870 ;
        RECT 38.225 168.815 39.325 168.840 ;
        RECT 38.225 168.780 39.360 168.815 ;
        RECT 38.225 168.775 39.390 168.780 ;
        RECT 38.225 168.380 38.455 168.775 ;
        RECT 39.000 168.770 39.390 168.775 ;
        RECT 39.025 168.760 39.390 168.770 ;
        RECT 39.040 168.755 39.390 168.760 ;
        RECT 39.055 168.750 39.390 168.755 ;
        RECT 39.755 168.750 40.015 169.200 ;
        RECT 40.185 168.935 41.395 170.025 ;
        RECT 39.055 168.745 40.015 168.750 ;
        RECT 39.065 168.735 40.015 168.745 ;
        RECT 39.075 168.730 40.015 168.735 ;
        RECT 39.085 168.720 40.015 168.730 ;
        RECT 39.090 168.710 40.015 168.720 ;
        RECT 39.095 168.705 40.015 168.710 ;
        RECT 39.105 168.690 40.015 168.705 ;
        RECT 39.110 168.675 40.015 168.690 ;
        RECT 39.120 168.650 40.015 168.675 ;
        RECT 38.625 168.180 38.955 168.605 ;
        RECT 37.885 167.645 38.145 168.125 ;
        RECT 38.315 167.475 38.565 168.015 ;
        RECT 38.735 167.695 38.955 168.180 ;
        RECT 39.125 168.580 40.015 168.650 ;
        RECT 39.125 167.855 39.295 168.580 ;
        RECT 39.465 168.025 40.015 168.410 ;
        RECT 40.185 168.225 40.705 168.765 ;
        RECT 40.875 168.395 41.395 168.935 ;
        RECT 41.575 169.415 41.905 169.845 ;
        RECT 42.085 169.585 42.280 170.025 ;
        RECT 42.450 169.415 42.780 169.845 ;
        RECT 41.575 169.245 42.780 169.415 ;
        RECT 41.575 168.915 42.470 169.245 ;
        RECT 42.950 169.075 43.225 169.845 ;
        RECT 43.405 169.590 48.750 170.025 ;
        RECT 42.640 168.885 43.225 169.075 ;
        RECT 41.580 168.385 41.875 168.715 ;
        RECT 42.055 168.385 42.470 168.715 ;
        RECT 39.125 167.685 40.015 167.855 ;
        RECT 40.185 167.475 41.395 168.225 ;
        RECT 41.575 167.475 41.875 168.205 ;
        RECT 42.055 167.765 42.285 168.385 ;
        RECT 42.640 168.215 42.815 168.885 ;
        RECT 42.485 168.035 42.815 168.215 ;
        RECT 42.985 168.065 43.225 168.715 ;
        RECT 42.485 167.655 42.710 168.035 ;
        RECT 44.990 168.020 45.330 168.850 ;
        RECT 46.810 168.340 47.160 169.590 ;
        RECT 49.845 168.860 50.135 170.025 ;
        RECT 50.325 169.515 50.625 170.025 ;
        RECT 50.795 169.515 51.175 169.685 ;
        RECT 51.755 169.515 52.385 170.025 ;
        RECT 50.795 169.345 50.965 169.515 ;
        RECT 52.555 169.345 52.885 169.855 ;
        RECT 53.055 169.515 53.355 170.025 ;
        RECT 53.545 169.515 53.845 170.025 ;
        RECT 54.015 169.515 54.395 169.685 ;
        RECT 54.975 169.515 55.605 170.025 ;
        RECT 54.015 169.345 54.185 169.515 ;
        RECT 55.775 169.345 56.105 169.855 ;
        RECT 56.275 169.515 56.575 170.025 ;
        RECT 50.305 169.145 50.965 169.345 ;
        RECT 51.135 169.175 53.355 169.345 ;
        RECT 50.305 168.215 50.475 169.145 ;
        RECT 51.135 168.975 51.305 169.175 ;
        RECT 50.645 168.805 51.305 168.975 ;
        RECT 51.475 168.835 53.015 169.005 ;
        RECT 50.645 168.385 50.815 168.805 ;
        RECT 51.475 168.635 51.645 168.835 ;
        RECT 51.045 168.465 51.645 168.635 ;
        RECT 51.815 168.465 52.510 168.665 ;
        RECT 52.770 168.385 53.015 168.835 ;
        RECT 51.135 168.215 52.045 168.295 ;
        RECT 42.880 167.475 43.210 167.865 ;
        RECT 43.405 167.475 48.750 168.020 ;
        RECT 49.845 167.475 50.135 168.200 ;
        RECT 50.305 167.735 50.625 168.215 ;
        RECT 50.795 168.125 52.045 168.215 ;
        RECT 50.795 168.045 51.305 168.125 ;
        RECT 50.795 167.645 51.025 168.045 ;
        RECT 51.195 167.475 51.545 167.865 ;
        RECT 51.715 167.645 52.045 168.125 ;
        RECT 52.215 167.475 52.385 168.295 ;
        RECT 53.185 168.215 53.355 169.175 ;
        RECT 52.890 167.670 53.355 168.215 ;
        RECT 53.525 169.145 54.185 169.345 ;
        RECT 54.355 169.175 56.575 169.345 ;
        RECT 53.525 168.215 53.695 169.145 ;
        RECT 54.355 168.975 54.525 169.175 ;
        RECT 53.865 168.805 54.525 168.975 ;
        RECT 54.695 168.835 56.235 169.005 ;
        RECT 53.865 168.385 54.035 168.805 ;
        RECT 54.695 168.635 54.865 168.835 ;
        RECT 54.265 168.465 54.865 168.635 ;
        RECT 55.035 168.465 55.730 168.665 ;
        RECT 55.990 168.385 56.235 168.835 ;
        RECT 54.355 168.215 55.265 168.295 ;
        RECT 53.525 167.735 53.845 168.215 ;
        RECT 54.015 168.125 55.265 168.215 ;
        RECT 54.015 168.045 54.525 168.125 ;
        RECT 54.015 167.645 54.245 168.045 ;
        RECT 54.415 167.475 54.765 167.865 ;
        RECT 54.935 167.645 55.265 168.125 ;
        RECT 55.435 167.475 55.605 168.295 ;
        RECT 56.405 168.215 56.575 169.175 ;
        RECT 56.110 167.670 56.575 168.215 ;
        RECT 56.745 168.420 57.025 169.855 ;
        RECT 57.195 169.250 57.905 170.025 ;
        RECT 58.075 169.080 58.405 169.855 ;
        RECT 57.255 168.865 58.405 169.080 ;
        RECT 56.745 167.645 57.085 168.420 ;
        RECT 57.255 168.295 57.540 168.865 ;
        RECT 57.725 168.465 58.195 168.695 ;
        RECT 58.600 168.665 58.815 169.780 ;
        RECT 58.995 169.305 59.325 170.025 ;
        RECT 59.105 168.665 59.335 169.005 ;
        RECT 59.565 168.885 59.775 170.025 ;
        RECT 58.365 168.485 58.815 168.665 ;
        RECT 58.365 168.465 58.695 168.485 ;
        RECT 59.005 168.465 59.335 168.665 ;
        RECT 59.945 168.875 60.275 169.855 ;
        RECT 60.445 168.885 60.675 170.025 ;
        RECT 60.885 169.590 66.230 170.025 ;
        RECT 57.255 168.105 57.965 168.295 ;
        RECT 57.665 167.965 57.965 168.105 ;
        RECT 58.155 168.105 59.335 168.295 ;
        RECT 58.155 168.025 58.485 168.105 ;
        RECT 57.665 167.955 57.980 167.965 ;
        RECT 57.665 167.945 57.990 167.955 ;
        RECT 57.665 167.940 58.000 167.945 ;
        RECT 57.255 167.475 57.425 167.935 ;
        RECT 57.665 167.930 58.005 167.940 ;
        RECT 57.665 167.925 58.010 167.930 ;
        RECT 57.665 167.915 58.015 167.925 ;
        RECT 57.665 167.910 58.020 167.915 ;
        RECT 57.665 167.645 58.025 167.910 ;
        RECT 58.655 167.475 58.825 167.935 ;
        RECT 58.995 167.645 59.335 168.105 ;
        RECT 59.565 167.475 59.775 168.295 ;
        RECT 59.945 168.275 60.195 168.875 ;
        RECT 60.365 168.465 60.695 168.715 ;
        RECT 59.945 167.645 60.275 168.275 ;
        RECT 60.445 167.475 60.675 168.295 ;
        RECT 62.470 168.020 62.810 168.850 ;
        RECT 64.290 168.340 64.640 169.590 ;
        RECT 66.955 169.355 67.125 169.855 ;
        RECT 67.295 169.525 67.625 170.025 ;
        RECT 66.955 169.185 67.620 169.355 ;
        RECT 66.870 168.365 67.220 169.015 ;
        RECT 67.390 168.195 67.620 169.185 ;
        RECT 66.955 168.025 67.620 168.195 ;
        RECT 60.885 167.475 66.230 168.020 ;
        RECT 66.955 167.735 67.125 168.025 ;
        RECT 67.295 167.475 67.625 167.855 ;
        RECT 67.795 167.735 67.980 169.855 ;
        RECT 68.220 169.565 68.485 170.025 ;
        RECT 68.655 169.430 68.905 169.855 ;
        RECT 69.115 169.580 70.220 169.750 ;
        RECT 68.600 169.300 68.905 169.430 ;
        RECT 68.150 168.105 68.430 169.055 ;
        RECT 68.600 168.195 68.770 169.300 ;
        RECT 68.940 168.515 69.180 169.110 ;
        RECT 69.350 169.045 69.880 169.410 ;
        RECT 69.350 168.345 69.520 169.045 ;
        RECT 70.050 168.965 70.220 169.580 ;
        RECT 70.390 169.225 70.560 170.025 ;
        RECT 70.730 169.525 70.980 169.855 ;
        RECT 71.205 169.555 72.090 169.725 ;
        RECT 70.050 168.875 70.560 168.965 ;
        RECT 68.600 168.065 68.825 168.195 ;
        RECT 68.995 168.125 69.520 168.345 ;
        RECT 69.690 168.705 70.560 168.875 ;
        RECT 68.235 167.475 68.485 167.935 ;
        RECT 68.655 167.925 68.825 168.065 ;
        RECT 69.690 167.925 69.860 168.705 ;
        RECT 70.390 168.635 70.560 168.705 ;
        RECT 70.070 168.455 70.270 168.485 ;
        RECT 70.730 168.455 70.900 169.525 ;
        RECT 71.070 168.635 71.260 169.355 ;
        RECT 70.070 168.155 70.900 168.455 ;
        RECT 71.430 168.425 71.750 169.385 ;
        RECT 68.655 167.755 68.990 167.925 ;
        RECT 69.185 167.755 69.860 167.925 ;
        RECT 70.180 167.475 70.550 167.975 ;
        RECT 70.730 167.925 70.900 168.155 ;
        RECT 71.285 168.095 71.750 168.425 ;
        RECT 71.920 168.715 72.090 169.555 ;
        RECT 72.270 169.525 72.585 170.025 ;
        RECT 72.815 169.295 73.155 169.855 ;
        RECT 72.260 168.920 73.155 169.295 ;
        RECT 73.325 169.015 73.495 170.025 ;
        RECT 72.965 168.715 73.155 168.920 ;
        RECT 73.665 168.965 73.995 169.810 ;
        RECT 73.665 168.885 74.055 168.965 ;
        RECT 74.225 168.935 75.435 170.025 ;
        RECT 73.840 168.835 74.055 168.885 ;
        RECT 71.920 168.385 72.795 168.715 ;
        RECT 72.965 168.385 73.715 168.715 ;
        RECT 71.920 167.925 72.090 168.385 ;
        RECT 72.965 168.215 73.165 168.385 ;
        RECT 73.885 168.255 74.055 168.835 ;
        RECT 73.830 168.215 74.055 168.255 ;
        RECT 70.730 167.755 71.135 167.925 ;
        RECT 71.305 167.755 72.090 167.925 ;
        RECT 72.365 167.475 72.575 168.005 ;
        RECT 72.835 167.690 73.165 168.215 ;
        RECT 73.675 168.130 74.055 168.215 ;
        RECT 74.225 168.225 74.745 168.765 ;
        RECT 74.915 168.395 75.435 168.935 ;
        RECT 75.605 168.860 75.895 170.025 ;
        RECT 76.155 169.280 76.425 170.025 ;
        RECT 77.055 170.020 83.330 170.025 ;
        RECT 76.595 169.110 76.885 169.850 ;
        RECT 77.055 169.295 77.310 170.020 ;
        RECT 77.495 169.125 77.755 169.850 ;
        RECT 77.925 169.295 78.170 170.020 ;
        RECT 78.355 169.125 78.615 169.850 ;
        RECT 78.785 169.295 79.030 170.020 ;
        RECT 79.215 169.125 79.475 169.850 ;
        RECT 79.645 169.295 79.890 170.020 ;
        RECT 80.060 169.125 80.320 169.850 ;
        RECT 80.490 169.295 80.750 170.020 ;
        RECT 80.920 169.125 81.180 169.850 ;
        RECT 81.350 169.295 81.610 170.020 ;
        RECT 81.780 169.125 82.040 169.850 ;
        RECT 82.210 169.295 82.470 170.020 ;
        RECT 82.640 169.125 82.900 169.850 ;
        RECT 83.070 169.225 83.330 170.020 ;
        RECT 77.495 169.110 82.900 169.125 ;
        RECT 76.155 168.885 82.900 169.110 ;
        RECT 76.155 168.295 77.320 168.885 ;
        RECT 83.500 168.715 83.750 169.850 ;
        RECT 83.930 169.215 84.190 170.025 ;
        RECT 84.365 168.715 84.610 169.855 ;
        RECT 84.790 169.215 85.085 170.025 ;
        RECT 85.725 169.175 86.105 169.855 ;
        RECT 86.695 169.175 86.865 170.025 ;
        RECT 87.035 169.345 87.365 169.855 ;
        RECT 87.535 169.515 87.705 170.025 ;
        RECT 87.875 169.345 88.275 169.855 ;
        RECT 87.035 169.175 88.275 169.345 ;
        RECT 77.490 168.465 84.610 168.715 ;
        RECT 73.335 167.475 73.505 168.085 ;
        RECT 73.675 167.695 74.005 168.130 ;
        RECT 74.225 167.475 75.435 168.225 ;
        RECT 75.605 167.475 75.895 168.200 ;
        RECT 76.155 168.125 82.900 168.295 ;
        RECT 76.155 167.475 76.455 167.955 ;
        RECT 76.625 167.670 76.885 168.125 ;
        RECT 77.055 167.475 77.315 167.955 ;
        RECT 77.495 167.670 77.755 168.125 ;
        RECT 77.925 167.475 78.175 167.955 ;
        RECT 78.355 167.670 78.615 168.125 ;
        RECT 78.785 167.475 79.035 167.955 ;
        RECT 79.215 167.670 79.475 168.125 ;
        RECT 79.645 167.475 79.890 167.955 ;
        RECT 80.060 167.670 80.335 168.125 ;
        RECT 80.505 167.475 80.750 167.955 ;
        RECT 80.920 167.670 81.180 168.125 ;
        RECT 81.350 167.475 81.610 167.955 ;
        RECT 81.780 167.670 82.040 168.125 ;
        RECT 82.210 167.475 82.470 167.955 ;
        RECT 82.640 167.670 82.900 168.125 ;
        RECT 83.070 167.475 83.330 168.035 ;
        RECT 83.500 167.655 83.750 168.465 ;
        RECT 83.930 167.475 84.190 168.000 ;
        RECT 84.360 167.655 84.610 168.465 ;
        RECT 84.780 168.155 85.095 168.715 ;
        RECT 85.725 168.215 85.895 169.175 ;
        RECT 86.065 168.835 87.370 169.005 ;
        RECT 88.455 168.925 88.775 169.855 ;
        RECT 88.945 169.590 94.290 170.025 ;
        RECT 86.065 168.385 86.310 168.835 ;
        RECT 86.480 168.465 87.030 168.665 ;
        RECT 87.200 168.635 87.370 168.835 ;
        RECT 88.145 168.755 88.775 168.925 ;
        RECT 87.200 168.465 87.575 168.635 ;
        RECT 87.745 168.215 87.975 168.715 ;
        RECT 85.725 168.045 87.975 168.215 ;
        RECT 84.790 167.475 85.095 167.985 ;
        RECT 85.775 167.475 86.105 167.865 ;
        RECT 86.275 167.725 86.445 168.045 ;
        RECT 88.145 167.875 88.315 168.755 ;
        RECT 86.615 167.475 86.945 167.865 ;
        RECT 87.360 167.705 88.315 167.875 ;
        RECT 88.485 167.475 88.775 168.310 ;
        RECT 90.530 168.020 90.870 168.850 ;
        RECT 92.350 168.340 92.700 169.590 ;
        RECT 94.465 168.935 97.975 170.025 ;
        RECT 94.465 168.245 96.115 168.765 ;
        RECT 96.285 168.415 97.975 168.935 ;
        RECT 98.185 169.075 98.475 169.845 ;
        RECT 99.045 169.485 99.305 169.845 ;
        RECT 99.475 169.655 99.805 170.025 ;
        RECT 99.975 169.485 100.235 169.845 ;
        RECT 99.045 169.255 100.235 169.485 ;
        RECT 100.425 169.305 100.755 170.025 ;
        RECT 100.925 169.075 101.190 169.845 ;
        RECT 98.185 168.895 100.680 169.075 ;
        RECT 98.155 168.385 98.425 168.715 ;
        RECT 98.605 168.385 99.040 168.715 ;
        RECT 99.220 168.385 99.795 168.715 ;
        RECT 99.975 168.385 100.255 168.715 ;
        RECT 88.945 167.475 94.290 168.020 ;
        RECT 94.465 167.475 97.975 168.245 ;
        RECT 100.455 168.205 100.680 168.895 ;
        RECT 98.195 168.015 100.680 168.205 ;
        RECT 98.195 167.655 98.420 168.015 ;
        RECT 98.600 167.475 98.930 167.845 ;
        RECT 99.110 167.655 99.365 168.015 ;
        RECT 99.930 167.475 100.675 167.845 ;
        RECT 100.855 167.655 101.190 169.075 ;
        RECT 101.365 168.860 101.655 170.025 ;
        RECT 101.915 169.355 102.085 169.855 ;
        RECT 102.255 169.525 102.585 170.025 ;
        RECT 101.915 169.185 102.580 169.355 ;
        RECT 101.830 168.365 102.180 169.015 ;
        RECT 101.365 167.475 101.655 168.200 ;
        RECT 102.350 168.195 102.580 169.185 ;
        RECT 101.915 168.025 102.580 168.195 ;
        RECT 101.915 167.735 102.085 168.025 ;
        RECT 102.255 167.475 102.585 167.855 ;
        RECT 102.755 167.735 102.940 169.855 ;
        RECT 103.180 169.565 103.445 170.025 ;
        RECT 103.615 169.430 103.865 169.855 ;
        RECT 104.075 169.580 105.180 169.750 ;
        RECT 103.560 169.300 103.865 169.430 ;
        RECT 103.110 168.105 103.390 169.055 ;
        RECT 103.560 168.195 103.730 169.300 ;
        RECT 103.900 168.515 104.140 169.110 ;
        RECT 104.310 169.045 104.840 169.410 ;
        RECT 104.310 168.345 104.480 169.045 ;
        RECT 105.010 168.965 105.180 169.580 ;
        RECT 105.350 169.225 105.520 170.025 ;
        RECT 105.690 169.525 105.940 169.855 ;
        RECT 106.165 169.555 107.050 169.725 ;
        RECT 105.010 168.875 105.520 168.965 ;
        RECT 103.560 168.065 103.785 168.195 ;
        RECT 103.955 168.125 104.480 168.345 ;
        RECT 104.650 168.705 105.520 168.875 ;
        RECT 103.195 167.475 103.445 167.935 ;
        RECT 103.615 167.925 103.785 168.065 ;
        RECT 104.650 167.925 104.820 168.705 ;
        RECT 105.350 168.635 105.520 168.705 ;
        RECT 105.030 168.455 105.230 168.485 ;
        RECT 105.690 168.455 105.860 169.525 ;
        RECT 106.030 168.635 106.220 169.355 ;
        RECT 105.030 168.155 105.860 168.455 ;
        RECT 106.390 168.425 106.710 169.385 ;
        RECT 103.615 167.755 103.950 167.925 ;
        RECT 104.145 167.755 104.820 167.925 ;
        RECT 105.140 167.475 105.510 167.975 ;
        RECT 105.690 167.925 105.860 168.155 ;
        RECT 106.245 168.095 106.710 168.425 ;
        RECT 106.880 168.715 107.050 169.555 ;
        RECT 107.230 169.525 107.545 170.025 ;
        RECT 107.775 169.295 108.115 169.855 ;
        RECT 107.220 168.920 108.115 169.295 ;
        RECT 108.285 169.015 108.455 170.025 ;
        RECT 107.925 168.715 108.115 168.920 ;
        RECT 108.625 168.965 108.955 169.810 ;
        RECT 109.125 169.110 109.295 170.025 ;
        RECT 109.695 169.010 109.950 169.850 ;
        RECT 110.125 169.205 110.455 170.025 ;
        RECT 110.695 169.035 110.905 169.850 ;
        RECT 108.625 168.885 109.015 168.965 ;
        RECT 108.800 168.835 109.015 168.885 ;
        RECT 106.880 168.385 107.755 168.715 ;
        RECT 107.925 168.385 108.675 168.715 ;
        RECT 106.880 167.925 107.050 168.385 ;
        RECT 107.925 168.215 108.125 168.385 ;
        RECT 108.845 168.255 109.015 168.835 ;
        RECT 108.790 168.215 109.015 168.255 ;
        RECT 105.690 167.755 106.095 167.925 ;
        RECT 106.265 167.755 107.050 167.925 ;
        RECT 107.325 167.475 107.535 168.005 ;
        RECT 107.795 167.690 108.125 168.215 ;
        RECT 108.635 168.130 109.015 168.215 ;
        RECT 108.295 167.475 108.465 168.085 ;
        RECT 108.635 167.695 108.965 168.130 ;
        RECT 109.135 167.475 109.305 167.990 ;
        RECT 109.695 167.645 110.025 169.010 ;
        RECT 110.255 168.855 110.905 169.035 ;
        RECT 110.255 168.215 110.475 168.855 ;
        RECT 111.075 168.680 111.280 169.855 ;
        RECT 110.850 168.440 111.280 168.680 ;
        RECT 111.450 168.440 111.780 169.855 ;
        RECT 111.960 168.385 112.240 169.855 ;
        RECT 112.420 169.055 112.705 169.850 ;
        RECT 112.885 169.225 113.100 170.025 ;
        RECT 113.280 169.055 113.550 169.850 ;
        RECT 112.420 168.885 113.550 169.055 ;
        RECT 113.785 168.935 116.375 170.025 ;
        RECT 112.465 168.385 112.850 168.715 ;
        RECT 113.070 168.415 113.570 168.680 ;
        RECT 112.545 168.235 112.850 168.385 ;
        RECT 113.785 168.245 114.995 168.765 ;
        RECT 115.165 168.415 116.375 168.935 ;
        RECT 116.545 169.155 116.820 169.855 ;
        RECT 116.990 169.480 117.245 170.025 ;
        RECT 117.415 169.515 117.895 169.855 ;
        RECT 118.070 169.470 118.675 170.025 ;
        RECT 118.060 169.370 118.675 169.470 ;
        RECT 118.060 169.345 118.245 169.370 ;
        RECT 110.255 168.045 112.365 168.215 ;
        RECT 110.255 168.040 111.475 168.045 ;
        RECT 110.195 167.475 110.870 167.860 ;
        RECT 111.145 167.650 111.475 168.040 ;
        RECT 111.645 167.475 111.990 167.875 ;
        RECT 112.160 167.650 112.365 168.045 ;
        RECT 112.545 167.675 113.100 168.235 ;
        RECT 113.275 167.475 113.515 168.150 ;
        RECT 113.785 167.475 116.375 168.245 ;
        RECT 116.545 168.125 116.715 169.155 ;
        RECT 116.990 169.025 117.745 169.275 ;
        RECT 117.915 169.100 118.245 169.345 ;
        RECT 116.990 168.990 117.760 169.025 ;
        RECT 116.990 168.980 117.775 168.990 ;
        RECT 116.885 168.965 117.780 168.980 ;
        RECT 116.885 168.950 117.800 168.965 ;
        RECT 116.885 168.940 117.820 168.950 ;
        RECT 116.885 168.930 117.845 168.940 ;
        RECT 116.885 168.900 117.915 168.930 ;
        RECT 116.885 168.870 117.935 168.900 ;
        RECT 116.885 168.840 117.955 168.870 ;
        RECT 116.885 168.815 117.985 168.840 ;
        RECT 116.885 168.780 118.020 168.815 ;
        RECT 116.885 168.775 118.050 168.780 ;
        RECT 116.885 168.380 117.115 168.775 ;
        RECT 117.660 168.770 118.050 168.775 ;
        RECT 117.685 168.760 118.050 168.770 ;
        RECT 117.700 168.755 118.050 168.760 ;
        RECT 117.715 168.750 118.050 168.755 ;
        RECT 118.415 168.750 118.675 169.200 ;
        RECT 118.845 168.885 119.105 170.025 ;
        RECT 119.275 168.875 119.605 169.855 ;
        RECT 119.775 168.885 120.055 170.025 ;
        RECT 121.345 169.355 121.625 170.025 ;
        RECT 121.795 169.135 122.095 169.685 ;
        RECT 122.295 169.305 122.625 170.025 ;
        RECT 122.815 169.305 123.275 169.855 ;
        RECT 119.365 168.835 119.540 168.875 ;
        RECT 117.715 168.745 118.675 168.750 ;
        RECT 117.725 168.735 118.675 168.745 ;
        RECT 117.735 168.730 118.675 168.735 ;
        RECT 117.745 168.720 118.675 168.730 ;
        RECT 117.750 168.710 118.675 168.720 ;
        RECT 117.755 168.705 118.675 168.710 ;
        RECT 117.765 168.690 118.675 168.705 ;
        RECT 117.770 168.675 118.675 168.690 ;
        RECT 117.780 168.650 118.675 168.675 ;
        RECT 117.285 168.180 117.615 168.605 ;
        RECT 116.545 167.645 116.805 168.125 ;
        RECT 116.975 167.475 117.225 168.015 ;
        RECT 117.395 167.695 117.615 168.180 ;
        RECT 117.785 168.580 118.675 168.650 ;
        RECT 117.785 167.855 117.955 168.580 ;
        RECT 118.865 168.465 119.200 168.715 ;
        RECT 118.125 168.025 118.675 168.410 ;
        RECT 119.370 168.275 119.540 168.835 ;
        RECT 121.160 168.715 121.425 169.075 ;
        RECT 121.795 168.965 122.735 169.135 ;
        RECT 122.565 168.715 122.735 168.965 ;
        RECT 119.710 168.445 120.045 168.715 ;
        RECT 121.160 168.465 121.835 168.715 ;
        RECT 122.055 168.465 122.395 168.715 ;
        RECT 122.565 168.385 122.855 168.715 ;
        RECT 122.565 168.295 122.735 168.385 ;
        RECT 117.785 167.685 118.675 167.855 ;
        RECT 118.845 167.645 119.540 168.275 ;
        RECT 119.745 167.475 120.055 168.275 ;
        RECT 121.345 168.105 122.735 168.295 ;
        RECT 121.345 167.745 121.675 168.105 ;
        RECT 123.025 167.935 123.275 169.305 ;
        RECT 122.295 167.475 122.545 167.935 ;
        RECT 122.715 167.645 123.275 167.935 ;
        RECT 124.365 168.950 124.635 169.855 ;
        RECT 124.805 169.265 125.135 170.025 ;
        RECT 125.315 169.095 125.485 169.855 ;
        RECT 124.365 168.150 124.535 168.950 ;
        RECT 124.820 168.925 125.485 169.095 ;
        RECT 125.745 168.935 126.955 170.025 ;
        RECT 124.820 168.780 124.990 168.925 ;
        RECT 124.705 168.450 124.990 168.780 ;
        RECT 124.820 168.195 124.990 168.450 ;
        RECT 125.225 168.375 125.555 168.745 ;
        RECT 125.745 168.225 126.265 168.765 ;
        RECT 126.435 168.395 126.955 168.935 ;
        RECT 127.125 168.860 127.415 170.025 ;
        RECT 127.585 169.590 132.930 170.025 ;
        RECT 133.105 169.590 138.450 170.025 ;
        RECT 138.625 169.590 143.970 170.025 ;
        RECT 124.365 167.645 124.625 168.150 ;
        RECT 124.820 168.025 125.485 168.195 ;
        RECT 124.805 167.475 125.135 167.855 ;
        RECT 125.315 167.645 125.485 168.025 ;
        RECT 125.745 167.475 126.955 168.225 ;
        RECT 127.125 167.475 127.415 168.200 ;
        RECT 129.170 168.020 129.510 168.850 ;
        RECT 130.990 168.340 131.340 169.590 ;
        RECT 134.690 168.020 135.030 168.850 ;
        RECT 136.510 168.340 136.860 169.590 ;
        RECT 140.210 168.020 140.550 168.850 ;
        RECT 142.030 168.340 142.380 169.590 ;
        RECT 144.145 168.935 147.655 170.025 ;
        RECT 147.825 168.935 149.035 170.025 ;
        RECT 144.145 168.245 145.795 168.765 ;
        RECT 145.965 168.415 147.655 168.935 ;
        RECT 127.585 167.475 132.930 168.020 ;
        RECT 133.105 167.475 138.450 168.020 ;
        RECT 138.625 167.475 143.970 168.020 ;
        RECT 144.145 167.475 147.655 168.245 ;
        RECT 147.825 168.225 148.345 168.765 ;
        RECT 148.515 168.395 149.035 168.935 ;
        RECT 149.205 168.935 150.415 170.025 ;
        RECT 149.205 168.395 149.725 168.935 ;
        RECT 149.895 168.225 150.415 168.765 ;
        RECT 147.825 167.475 149.035 168.225 ;
        RECT 149.205 167.475 150.415 168.225 ;
        RECT 11.120 167.305 150.500 167.475 ;
        RECT 11.205 166.555 12.415 167.305 ;
        RECT 12.585 166.760 17.930 167.305 ;
        RECT 18.105 166.760 23.450 167.305 ;
        RECT 11.205 166.015 11.725 166.555 ;
        RECT 11.895 165.845 12.415 166.385 ;
        RECT 14.170 165.930 14.510 166.760 ;
        RECT 11.205 164.755 12.415 165.845 ;
        RECT 15.990 165.190 16.340 166.440 ;
        RECT 19.690 165.930 20.030 166.760 ;
        RECT 23.625 166.535 25.295 167.305 ;
        RECT 26.040 166.675 26.325 167.135 ;
        RECT 26.495 166.845 26.765 167.305 ;
        RECT 21.510 165.190 21.860 166.440 ;
        RECT 23.625 166.015 24.375 166.535 ;
        RECT 26.040 166.505 26.995 166.675 ;
        RECT 24.545 165.845 25.295 166.365 ;
        RECT 12.585 164.755 17.930 165.190 ;
        RECT 18.105 164.755 23.450 165.190 ;
        RECT 23.625 164.755 25.295 165.845 ;
        RECT 25.925 165.775 26.615 166.335 ;
        RECT 26.785 165.605 26.995 166.505 ;
        RECT 26.040 165.385 26.995 165.605 ;
        RECT 27.165 166.335 27.565 167.135 ;
        RECT 27.755 166.675 28.035 167.135 ;
        RECT 28.555 166.845 28.880 167.305 ;
        RECT 27.755 166.505 28.880 166.675 ;
        RECT 29.050 166.565 29.435 167.135 ;
        RECT 28.430 166.395 28.880 166.505 ;
        RECT 27.165 165.775 28.260 166.335 ;
        RECT 28.430 166.065 28.985 166.395 ;
        RECT 26.040 164.925 26.325 165.385 ;
        RECT 26.495 164.755 26.765 165.215 ;
        RECT 27.165 164.925 27.565 165.775 ;
        RECT 28.430 165.605 28.880 166.065 ;
        RECT 29.155 165.895 29.435 166.565 ;
        RECT 27.755 165.385 28.880 165.605 ;
        RECT 27.755 164.925 28.035 165.385 ;
        RECT 28.555 164.755 28.880 165.215 ;
        RECT 29.050 164.925 29.435 165.895 ;
        RECT 30.065 166.805 30.365 167.135 ;
        RECT 30.535 166.825 30.810 167.305 ;
        RECT 30.065 165.895 30.235 166.805 ;
        RECT 30.990 166.655 31.285 167.045 ;
        RECT 31.455 166.825 31.710 167.305 ;
        RECT 31.885 166.655 32.145 167.045 ;
        RECT 32.315 166.825 32.595 167.305 ;
        RECT 30.405 166.065 30.755 166.635 ;
        RECT 30.990 166.485 32.640 166.655 ;
        RECT 30.925 166.145 32.065 166.315 ;
        RECT 30.925 165.895 31.095 166.145 ;
        RECT 32.235 165.975 32.640 166.485 ;
        RECT 30.065 165.725 31.095 165.895 ;
        RECT 31.885 165.805 32.640 165.975 ;
        RECT 32.825 166.630 33.085 167.135 ;
        RECT 33.265 166.925 33.595 167.305 ;
        RECT 33.775 166.755 33.945 167.135 ;
        RECT 32.825 165.830 32.995 166.630 ;
        RECT 33.280 166.585 33.945 166.755 ;
        RECT 33.280 166.330 33.450 166.585 ;
        RECT 34.205 166.535 36.795 167.305 ;
        RECT 36.965 166.580 37.255 167.305 ;
        RECT 37.425 166.535 40.935 167.305 ;
        RECT 41.105 166.565 41.570 167.110 ;
        RECT 33.165 166.000 33.450 166.330 ;
        RECT 33.685 166.035 34.015 166.405 ;
        RECT 34.205 166.015 35.415 166.535 ;
        RECT 33.280 165.855 33.450 166.000 ;
        RECT 30.065 164.925 30.375 165.725 ;
        RECT 31.885 165.555 32.145 165.805 ;
        RECT 30.545 164.755 30.855 165.555 ;
        RECT 31.025 165.385 32.145 165.555 ;
        RECT 31.025 164.925 31.285 165.385 ;
        RECT 31.455 164.755 31.710 165.215 ;
        RECT 31.885 164.925 32.145 165.385 ;
        RECT 32.315 164.755 32.600 165.625 ;
        RECT 32.825 164.925 33.095 165.830 ;
        RECT 33.280 165.685 33.945 165.855 ;
        RECT 35.585 165.845 36.795 166.365 ;
        RECT 37.425 166.015 39.075 166.535 ;
        RECT 33.265 164.755 33.595 165.515 ;
        RECT 33.775 164.925 33.945 165.685 ;
        RECT 34.205 164.755 36.795 165.845 ;
        RECT 36.965 164.755 37.255 165.920 ;
        RECT 39.245 165.845 40.935 166.365 ;
        RECT 37.425 164.755 40.935 165.845 ;
        RECT 41.105 165.605 41.275 166.565 ;
        RECT 42.075 166.485 42.245 167.305 ;
        RECT 42.415 166.655 42.745 167.135 ;
        RECT 42.915 166.915 43.265 167.305 ;
        RECT 43.435 166.735 43.665 167.135 ;
        RECT 43.155 166.655 43.665 166.735 ;
        RECT 42.415 166.565 43.665 166.655 ;
        RECT 43.835 166.565 44.155 167.045 ;
        RECT 44.325 166.760 49.670 167.305 ;
        RECT 42.415 166.485 43.325 166.565 ;
        RECT 41.445 165.945 41.690 166.395 ;
        RECT 41.950 166.115 42.645 166.315 ;
        RECT 42.815 166.145 43.415 166.315 ;
        RECT 42.815 165.945 42.985 166.145 ;
        RECT 43.645 165.975 43.815 166.395 ;
        RECT 41.445 165.775 42.985 165.945 ;
        RECT 43.155 165.805 43.815 165.975 ;
        RECT 43.155 165.605 43.325 165.805 ;
        RECT 43.985 165.635 44.155 166.565 ;
        RECT 45.910 165.930 46.250 166.760 ;
        RECT 49.845 166.535 51.515 167.305 ;
        RECT 52.155 166.575 52.455 167.305 ;
        RECT 41.105 165.435 43.325 165.605 ;
        RECT 43.495 165.435 44.155 165.635 ;
        RECT 41.105 164.755 41.405 165.265 ;
        RECT 41.575 164.925 41.905 165.435 ;
        RECT 43.495 165.265 43.665 165.435 ;
        RECT 42.075 164.755 42.705 165.265 ;
        RECT 43.285 165.095 43.665 165.265 ;
        RECT 43.835 164.755 44.135 165.265 ;
        RECT 47.730 165.190 48.080 166.440 ;
        RECT 49.845 166.015 50.595 166.535 ;
        RECT 52.635 166.395 52.865 167.015 ;
        RECT 53.065 166.745 53.290 167.125 ;
        RECT 53.460 166.915 53.790 167.305 ;
        RECT 53.985 166.760 59.330 167.305 ;
        RECT 53.065 166.565 53.395 166.745 ;
        RECT 50.765 165.845 51.515 166.365 ;
        RECT 52.160 166.065 52.455 166.395 ;
        RECT 52.635 166.065 53.050 166.395 ;
        RECT 53.220 165.895 53.395 166.565 ;
        RECT 53.565 166.065 53.805 166.715 ;
        RECT 55.570 165.930 55.910 166.760 ;
        RECT 59.505 166.535 62.095 167.305 ;
        RECT 62.725 166.580 63.015 167.305 ;
        RECT 63.300 166.675 63.585 167.135 ;
        RECT 63.755 166.845 64.025 167.305 ;
        RECT 44.325 164.755 49.670 165.190 ;
        RECT 49.845 164.755 51.515 165.845 ;
        RECT 52.155 165.535 53.050 165.865 ;
        RECT 53.220 165.705 53.805 165.895 ;
        RECT 52.155 165.365 53.360 165.535 ;
        RECT 52.155 164.935 52.485 165.365 ;
        RECT 52.665 164.755 52.860 165.195 ;
        RECT 53.030 164.935 53.360 165.365 ;
        RECT 53.530 164.935 53.805 165.705 ;
        RECT 57.390 165.190 57.740 166.440 ;
        RECT 59.505 166.015 60.715 166.535 ;
        RECT 63.300 166.505 64.255 166.675 ;
        RECT 60.885 165.845 62.095 166.365 ;
        RECT 53.985 164.755 59.330 165.190 ;
        RECT 59.505 164.755 62.095 165.845 ;
        RECT 62.725 164.755 63.015 165.920 ;
        RECT 63.185 165.775 63.875 166.335 ;
        RECT 64.045 165.605 64.255 166.505 ;
        RECT 63.300 165.385 64.255 165.605 ;
        RECT 64.425 166.335 64.825 167.135 ;
        RECT 65.015 166.675 65.295 167.135 ;
        RECT 65.815 166.845 66.140 167.305 ;
        RECT 65.015 166.505 66.140 166.675 ;
        RECT 66.310 166.565 66.695 167.135 ;
        RECT 65.690 166.395 66.140 166.505 ;
        RECT 64.425 165.775 65.520 166.335 ;
        RECT 65.690 166.065 66.245 166.395 ;
        RECT 63.300 164.925 63.585 165.385 ;
        RECT 63.755 164.755 64.025 165.215 ;
        RECT 64.425 164.925 64.825 165.775 ;
        RECT 65.690 165.605 66.140 166.065 ;
        RECT 66.415 165.895 66.695 166.565 ;
        RECT 66.865 166.505 67.175 167.305 ;
        RECT 67.380 166.505 68.075 167.135 ;
        RECT 68.245 166.630 68.505 167.135 ;
        RECT 68.685 166.925 69.015 167.305 ;
        RECT 69.195 166.755 69.365 167.135 ;
        RECT 66.875 166.065 67.210 166.335 ;
        RECT 67.380 165.905 67.550 166.505 ;
        RECT 67.720 166.065 68.055 166.315 ;
        RECT 65.015 165.385 66.140 165.605 ;
        RECT 65.015 164.925 65.295 165.385 ;
        RECT 65.815 164.755 66.140 165.215 ;
        RECT 66.310 164.925 66.695 165.895 ;
        RECT 66.865 164.755 67.145 165.895 ;
        RECT 67.315 164.925 67.645 165.905 ;
        RECT 67.815 164.755 68.075 165.895 ;
        RECT 68.245 165.830 68.415 166.630 ;
        RECT 68.700 166.585 69.365 166.755 ;
        RECT 68.700 166.330 68.870 166.585 ;
        RECT 69.625 166.535 73.135 167.305 ;
        RECT 73.765 166.805 74.065 167.135 ;
        RECT 74.235 166.825 74.510 167.305 ;
        RECT 68.585 166.000 68.870 166.330 ;
        RECT 69.105 166.035 69.435 166.405 ;
        RECT 69.625 166.015 71.275 166.535 ;
        RECT 68.700 165.855 68.870 166.000 ;
        RECT 68.245 164.925 68.515 165.830 ;
        RECT 68.700 165.685 69.365 165.855 ;
        RECT 71.445 165.845 73.135 166.365 ;
        RECT 68.685 164.755 69.015 165.515 ;
        RECT 69.195 164.925 69.365 165.685 ;
        RECT 69.625 164.755 73.135 165.845 ;
        RECT 73.765 165.895 73.935 166.805 ;
        RECT 74.690 166.655 74.985 167.045 ;
        RECT 75.155 166.825 75.410 167.305 ;
        RECT 75.585 166.655 75.845 167.045 ;
        RECT 76.015 166.825 76.295 167.305 ;
        RECT 74.105 166.065 74.455 166.635 ;
        RECT 74.690 166.485 76.340 166.655 ;
        RECT 76.730 166.525 77.230 167.135 ;
        RECT 74.625 166.145 75.765 166.315 ;
        RECT 74.625 165.895 74.795 166.145 ;
        RECT 75.935 165.975 76.340 166.485 ;
        RECT 76.525 166.065 76.875 166.315 ;
        RECT 73.765 165.725 74.795 165.895 ;
        RECT 75.585 165.805 76.340 165.975 ;
        RECT 77.060 165.895 77.230 166.525 ;
        RECT 77.860 166.655 78.190 167.135 ;
        RECT 78.360 166.845 78.585 167.305 ;
        RECT 78.755 166.655 79.085 167.135 ;
        RECT 77.860 166.485 79.085 166.655 ;
        RECT 79.275 166.505 79.525 167.305 ;
        RECT 79.695 166.505 80.035 167.135 ;
        RECT 80.205 166.760 85.550 167.305 ;
        RECT 77.400 166.115 77.730 166.315 ;
        RECT 77.900 166.115 78.230 166.315 ;
        RECT 78.400 166.115 78.820 166.315 ;
        RECT 78.995 166.145 79.690 166.315 ;
        RECT 78.995 165.895 79.165 166.145 ;
        RECT 79.860 165.895 80.035 166.505 ;
        RECT 81.790 165.930 82.130 166.760 ;
        RECT 85.725 166.535 88.315 167.305 ;
        RECT 88.485 166.580 88.775 167.305 ;
        RECT 88.945 166.535 91.535 167.305 ;
        RECT 91.755 166.915 92.085 167.305 ;
        RECT 92.255 166.735 92.425 167.055 ;
        RECT 92.595 166.915 92.925 167.305 ;
        RECT 93.340 166.905 94.295 167.075 ;
        RECT 91.705 166.565 93.955 166.735 ;
        RECT 73.765 164.925 74.075 165.725 ;
        RECT 75.585 165.555 75.845 165.805 ;
        RECT 76.730 165.725 79.165 165.895 ;
        RECT 74.245 164.755 74.555 165.555 ;
        RECT 74.725 165.385 75.845 165.555 ;
        RECT 74.725 164.925 74.985 165.385 ;
        RECT 75.155 164.755 75.410 165.215 ;
        RECT 75.585 164.925 75.845 165.385 ;
        RECT 76.015 164.755 76.300 165.625 ;
        RECT 76.730 164.925 77.060 165.725 ;
        RECT 77.230 164.755 77.560 165.555 ;
        RECT 77.860 164.925 78.190 165.725 ;
        RECT 78.835 164.755 79.085 165.555 ;
        RECT 79.355 164.755 79.525 165.895 ;
        RECT 79.695 164.925 80.035 165.895 ;
        RECT 83.610 165.190 83.960 166.440 ;
        RECT 85.725 166.015 86.935 166.535 ;
        RECT 87.105 165.845 88.315 166.365 ;
        RECT 88.945 166.015 90.155 166.535 ;
        RECT 80.205 164.755 85.550 165.190 ;
        RECT 85.725 164.755 88.315 165.845 ;
        RECT 88.485 164.755 88.775 165.920 ;
        RECT 90.325 165.845 91.535 166.365 ;
        RECT 88.945 164.755 91.535 165.845 ;
        RECT 91.705 165.605 91.875 166.565 ;
        RECT 92.045 165.945 92.290 166.395 ;
        RECT 92.460 166.115 93.010 166.315 ;
        RECT 93.180 166.145 93.555 166.315 ;
        RECT 93.180 165.945 93.350 166.145 ;
        RECT 93.725 166.065 93.955 166.565 ;
        RECT 92.045 165.775 93.350 165.945 ;
        RECT 94.125 166.025 94.295 166.905 ;
        RECT 94.465 166.470 94.755 167.305 ;
        RECT 94.950 166.915 95.280 167.305 ;
        RECT 95.450 166.745 95.675 167.125 ;
        RECT 94.935 166.065 95.175 166.715 ;
        RECT 95.345 166.565 95.675 166.745 ;
        RECT 94.125 165.855 94.755 166.025 ;
        RECT 95.345 165.895 95.520 166.565 ;
        RECT 95.875 166.395 96.105 167.015 ;
        RECT 96.285 166.575 96.585 167.305 ;
        RECT 96.765 166.535 100.275 167.305 ;
        RECT 101.390 166.915 101.720 167.305 ;
        RECT 101.890 166.745 102.115 167.125 ;
        RECT 95.690 166.065 96.105 166.395 ;
        RECT 96.285 166.065 96.580 166.395 ;
        RECT 96.765 166.015 98.415 166.535 ;
        RECT 91.705 164.925 92.085 165.605 ;
        RECT 92.675 164.755 92.845 165.605 ;
        RECT 93.015 165.435 94.255 165.605 ;
        RECT 93.015 164.925 93.345 165.435 ;
        RECT 93.515 164.755 93.685 165.265 ;
        RECT 93.855 164.925 94.255 165.435 ;
        RECT 94.435 164.925 94.755 165.855 ;
        RECT 94.935 165.705 95.520 165.895 ;
        RECT 94.935 164.935 95.210 165.705 ;
        RECT 95.690 165.535 96.585 165.865 ;
        RECT 98.585 165.845 100.275 166.365 ;
        RECT 101.375 166.065 101.615 166.715 ;
        RECT 101.785 166.565 102.115 166.745 ;
        RECT 101.785 165.895 101.960 166.565 ;
        RECT 102.315 166.395 102.545 167.015 ;
        RECT 102.725 166.575 103.025 167.305 ;
        RECT 103.205 166.535 106.715 167.305 ;
        RECT 107.810 166.565 108.065 167.135 ;
        RECT 108.235 166.905 108.565 167.305 ;
        RECT 108.990 166.770 109.520 167.135 ;
        RECT 108.990 166.735 109.165 166.770 ;
        RECT 108.235 166.565 109.165 166.735 ;
        RECT 102.130 166.065 102.545 166.395 ;
        RECT 102.725 166.065 103.020 166.395 ;
        RECT 103.205 166.015 104.855 166.535 ;
        RECT 95.380 165.365 96.585 165.535 ;
        RECT 95.380 164.935 95.710 165.365 ;
        RECT 95.880 164.755 96.075 165.195 ;
        RECT 96.255 164.935 96.585 165.365 ;
        RECT 96.765 164.755 100.275 165.845 ;
        RECT 101.375 165.705 101.960 165.895 ;
        RECT 101.375 164.935 101.650 165.705 ;
        RECT 102.130 165.535 103.025 165.865 ;
        RECT 105.025 165.845 106.715 166.365 ;
        RECT 101.820 165.365 103.025 165.535 ;
        RECT 101.820 164.935 102.150 165.365 ;
        RECT 102.320 164.755 102.515 165.195 ;
        RECT 102.695 164.935 103.025 165.365 ;
        RECT 103.205 164.755 106.715 165.845 ;
        RECT 107.810 165.895 107.980 166.565 ;
        RECT 108.235 166.395 108.405 166.565 ;
        RECT 108.150 166.065 108.405 166.395 ;
        RECT 108.630 166.065 108.825 166.395 ;
        RECT 107.810 164.925 108.145 165.895 ;
        RECT 108.315 164.755 108.485 165.895 ;
        RECT 108.655 165.095 108.825 166.065 ;
        RECT 108.995 165.435 109.165 166.565 ;
        RECT 109.335 165.775 109.505 166.575 ;
        RECT 109.710 166.285 109.985 167.135 ;
        RECT 109.705 166.115 109.985 166.285 ;
        RECT 109.710 165.975 109.985 166.115 ;
        RECT 110.155 165.775 110.345 167.135 ;
        RECT 110.525 166.770 111.035 167.305 ;
        RECT 111.255 166.495 111.500 167.100 ;
        RECT 112.035 166.625 112.205 167.000 ;
        RECT 110.545 166.325 111.775 166.495 ;
        RECT 112.005 166.455 112.205 166.625 ;
        RECT 112.395 166.775 112.625 167.080 ;
        RECT 112.795 166.945 113.125 167.305 ;
        RECT 113.320 166.775 113.610 167.125 ;
        RECT 112.395 166.605 113.610 166.775 ;
        RECT 114.245 166.580 114.535 167.305 ;
        RECT 109.335 165.605 110.345 165.775 ;
        RECT 110.515 165.760 111.265 165.950 ;
        RECT 108.995 165.265 110.120 165.435 ;
        RECT 110.515 165.095 110.685 165.760 ;
        RECT 111.435 165.515 111.775 166.325 ;
        RECT 112.035 166.435 112.205 166.455 ;
        RECT 114.705 166.535 118.215 167.305 ;
        RECT 118.475 166.755 118.645 167.135 ;
        RECT 118.860 166.925 119.190 167.305 ;
        RECT 118.475 166.585 119.190 166.755 ;
        RECT 112.035 166.265 112.555 166.435 ;
        RECT 111.950 165.735 112.195 166.095 ;
        RECT 112.385 165.885 112.555 166.265 ;
        RECT 112.725 166.065 113.110 166.395 ;
        RECT 113.290 166.285 113.550 166.395 ;
        RECT 113.290 166.115 113.555 166.285 ;
        RECT 113.290 166.065 113.550 166.115 ;
        RECT 112.385 165.605 112.735 165.885 ;
        RECT 108.655 164.925 110.685 165.095 ;
        RECT 110.855 164.755 111.025 165.515 ;
        RECT 111.260 165.105 111.775 165.515 ;
        RECT 111.950 164.755 112.205 165.555 ;
        RECT 112.405 164.925 112.735 165.605 ;
        RECT 112.915 165.015 113.110 166.065 ;
        RECT 114.705 166.015 116.355 166.535 ;
        RECT 113.290 164.755 113.610 165.895 ;
        RECT 114.245 164.755 114.535 165.920 ;
        RECT 116.525 165.845 118.215 166.365 ;
        RECT 118.385 166.035 118.740 166.405 ;
        RECT 119.020 166.395 119.190 166.585 ;
        RECT 119.360 166.560 119.615 167.135 ;
        RECT 119.020 166.065 119.275 166.395 ;
        RECT 119.020 165.855 119.190 166.065 ;
        RECT 114.705 164.755 118.215 165.845 ;
        RECT 118.475 165.685 119.190 165.855 ;
        RECT 119.445 165.830 119.615 166.560 ;
        RECT 119.790 166.465 120.050 167.305 ;
        RECT 120.225 166.535 123.735 167.305 ;
        RECT 123.905 166.555 125.115 167.305 ;
        RECT 120.225 166.015 121.875 166.535 ;
        RECT 118.475 164.925 118.645 165.685 ;
        RECT 118.860 164.755 119.190 165.515 ;
        RECT 119.360 164.925 119.615 165.830 ;
        RECT 119.790 164.755 120.050 165.905 ;
        RECT 122.045 165.845 123.735 166.365 ;
        RECT 123.905 166.015 124.425 166.555 ;
        RECT 125.435 166.505 125.765 167.305 ;
        RECT 125.935 166.655 126.105 167.135 ;
        RECT 126.275 166.825 126.605 167.305 ;
        RECT 126.775 166.655 126.945 167.135 ;
        RECT 127.195 166.825 127.435 167.305 ;
        RECT 127.615 166.655 127.785 167.135 ;
        RECT 128.045 166.760 133.390 167.305 ;
        RECT 133.565 166.760 138.910 167.305 ;
        RECT 125.935 166.485 126.945 166.655 ;
        RECT 127.150 166.485 127.785 166.655 ;
        RECT 125.935 166.455 126.435 166.485 ;
        RECT 124.595 165.845 125.115 166.385 ;
        RECT 125.935 165.945 126.430 166.455 ;
        RECT 127.150 166.315 127.320 166.485 ;
        RECT 126.820 166.145 127.320 166.315 ;
        RECT 120.225 164.755 123.735 165.845 ;
        RECT 123.905 164.755 125.115 165.845 ;
        RECT 125.435 164.755 125.765 165.905 ;
        RECT 125.935 165.775 126.945 165.945 ;
        RECT 125.935 164.925 126.105 165.775 ;
        RECT 126.275 164.755 126.605 165.555 ;
        RECT 126.775 164.925 126.945 165.775 ;
        RECT 127.150 165.905 127.320 166.145 ;
        RECT 127.490 166.075 127.870 166.315 ;
        RECT 129.630 165.930 129.970 166.760 ;
        RECT 127.150 165.735 127.865 165.905 ;
        RECT 127.125 164.755 127.365 165.555 ;
        RECT 127.535 164.925 127.865 165.735 ;
        RECT 131.450 165.190 131.800 166.440 ;
        RECT 135.150 165.930 135.490 166.760 ;
        RECT 140.005 166.580 140.295 167.305 ;
        RECT 140.465 166.760 145.810 167.305 ;
        RECT 136.970 165.190 137.320 166.440 ;
        RECT 142.050 165.930 142.390 166.760 ;
        RECT 145.985 166.535 148.575 167.305 ;
        RECT 149.205 166.555 150.415 167.305 ;
        RECT 128.045 164.755 133.390 165.190 ;
        RECT 133.565 164.755 138.910 165.190 ;
        RECT 140.005 164.755 140.295 165.920 ;
        RECT 143.870 165.190 144.220 166.440 ;
        RECT 145.985 166.015 147.195 166.535 ;
        RECT 147.365 165.845 148.575 166.365 ;
        RECT 140.465 164.755 145.810 165.190 ;
        RECT 145.985 164.755 148.575 165.845 ;
        RECT 149.205 165.845 149.725 166.385 ;
        RECT 149.895 166.015 150.415 166.555 ;
        RECT 149.205 164.755 150.415 165.845 ;
        RECT 11.120 164.585 150.500 164.755 ;
        RECT 11.205 163.495 12.415 164.585 ;
        RECT 12.585 163.495 16.095 164.585 ;
        RECT 16.355 163.915 16.525 164.415 ;
        RECT 16.695 164.085 17.025 164.585 ;
        RECT 16.355 163.745 17.020 163.915 ;
        RECT 11.205 162.785 11.725 163.325 ;
        RECT 11.895 162.955 12.415 163.495 ;
        RECT 12.585 162.805 14.235 163.325 ;
        RECT 14.405 162.975 16.095 163.495 ;
        RECT 16.270 162.925 16.620 163.575 ;
        RECT 11.205 162.035 12.415 162.785 ;
        RECT 12.585 162.035 16.095 162.805 ;
        RECT 16.790 162.755 17.020 163.745 ;
        RECT 16.355 162.585 17.020 162.755 ;
        RECT 16.355 162.295 16.525 162.585 ;
        RECT 16.695 162.035 17.025 162.415 ;
        RECT 17.195 162.295 17.380 164.415 ;
        RECT 17.620 164.125 17.885 164.585 ;
        RECT 18.055 163.990 18.305 164.415 ;
        RECT 18.515 164.140 19.620 164.310 ;
        RECT 18.000 163.860 18.305 163.990 ;
        RECT 17.550 162.665 17.830 163.615 ;
        RECT 18.000 162.755 18.170 163.860 ;
        RECT 18.340 163.075 18.580 163.670 ;
        RECT 18.750 163.605 19.280 163.970 ;
        RECT 18.750 162.905 18.920 163.605 ;
        RECT 19.450 163.525 19.620 164.140 ;
        RECT 19.790 163.785 19.960 164.585 ;
        RECT 20.130 164.085 20.380 164.415 ;
        RECT 20.605 164.115 21.490 164.285 ;
        RECT 19.450 163.435 19.960 163.525 ;
        RECT 18.000 162.625 18.225 162.755 ;
        RECT 18.395 162.685 18.920 162.905 ;
        RECT 19.090 163.265 19.960 163.435 ;
        RECT 17.635 162.035 17.885 162.495 ;
        RECT 18.055 162.485 18.225 162.625 ;
        RECT 19.090 162.485 19.260 163.265 ;
        RECT 19.790 163.195 19.960 163.265 ;
        RECT 19.470 163.015 19.670 163.045 ;
        RECT 20.130 163.015 20.300 164.085 ;
        RECT 20.470 163.195 20.660 163.915 ;
        RECT 19.470 162.715 20.300 163.015 ;
        RECT 20.830 162.985 21.150 163.945 ;
        RECT 18.055 162.315 18.390 162.485 ;
        RECT 18.585 162.315 19.260 162.485 ;
        RECT 19.580 162.035 19.950 162.535 ;
        RECT 20.130 162.485 20.300 162.715 ;
        RECT 20.685 162.655 21.150 162.985 ;
        RECT 21.320 163.275 21.490 164.115 ;
        RECT 21.670 164.085 21.985 164.585 ;
        RECT 22.215 163.855 22.555 164.415 ;
        RECT 21.660 163.480 22.555 163.855 ;
        RECT 22.725 163.575 22.895 164.585 ;
        RECT 22.365 163.275 22.555 163.480 ;
        RECT 23.065 163.525 23.395 164.370 ;
        RECT 23.565 163.670 23.735 164.585 ;
        RECT 23.065 163.445 23.455 163.525 ;
        RECT 23.240 163.395 23.455 163.445 ;
        RECT 24.085 163.420 24.375 164.585 ;
        RECT 24.545 163.495 28.055 164.585 ;
        RECT 29.145 164.075 29.445 164.585 ;
        RECT 29.615 163.905 29.945 164.415 ;
        RECT 30.115 164.075 30.745 164.585 ;
        RECT 31.325 164.075 31.705 164.245 ;
        RECT 31.875 164.075 32.175 164.585 ;
        RECT 32.365 164.075 32.665 164.585 ;
        RECT 31.535 163.905 31.705 164.075 ;
        RECT 32.835 163.905 33.165 164.415 ;
        RECT 33.335 164.075 33.965 164.585 ;
        RECT 34.545 164.075 34.925 164.245 ;
        RECT 35.095 164.075 35.395 164.585 ;
        RECT 34.755 163.905 34.925 164.075 ;
        RECT 21.320 162.945 22.195 163.275 ;
        RECT 22.365 162.945 23.115 163.275 ;
        RECT 21.320 162.485 21.490 162.945 ;
        RECT 22.365 162.775 22.565 162.945 ;
        RECT 23.285 162.815 23.455 163.395 ;
        RECT 23.230 162.775 23.455 162.815 ;
        RECT 20.130 162.315 20.535 162.485 ;
        RECT 20.705 162.315 21.490 162.485 ;
        RECT 21.765 162.035 21.975 162.565 ;
        RECT 22.235 162.250 22.565 162.775 ;
        RECT 23.075 162.690 23.455 162.775 ;
        RECT 24.545 162.805 26.195 163.325 ;
        RECT 26.365 162.975 28.055 163.495 ;
        RECT 29.145 163.735 31.365 163.905 ;
        RECT 22.735 162.035 22.905 162.645 ;
        RECT 23.075 162.255 23.405 162.690 ;
        RECT 23.575 162.035 23.745 162.550 ;
        RECT 24.085 162.035 24.375 162.760 ;
        RECT 24.545 162.035 28.055 162.805 ;
        RECT 29.145 162.775 29.315 163.735 ;
        RECT 29.485 163.395 31.025 163.565 ;
        RECT 29.485 162.945 29.730 163.395 ;
        RECT 29.990 163.025 30.685 163.225 ;
        RECT 30.855 163.195 31.025 163.395 ;
        RECT 31.195 163.535 31.365 163.735 ;
        RECT 31.535 163.705 32.195 163.905 ;
        RECT 31.195 163.365 31.855 163.535 ;
        RECT 30.855 163.025 31.455 163.195 ;
        RECT 31.685 162.945 31.855 163.365 ;
        RECT 29.145 162.230 29.610 162.775 ;
        RECT 30.115 162.035 30.285 162.855 ;
        RECT 30.455 162.775 31.365 162.855 ;
        RECT 32.025 162.775 32.195 163.705 ;
        RECT 30.455 162.685 31.705 162.775 ;
        RECT 30.455 162.205 30.785 162.685 ;
        RECT 31.195 162.605 31.705 162.685 ;
        RECT 30.955 162.035 31.305 162.425 ;
        RECT 31.475 162.205 31.705 162.605 ;
        RECT 31.875 162.295 32.195 162.775 ;
        RECT 32.365 163.735 34.585 163.905 ;
        RECT 32.365 162.775 32.535 163.735 ;
        RECT 32.705 163.395 34.245 163.565 ;
        RECT 32.705 162.945 32.950 163.395 ;
        RECT 33.210 163.025 33.905 163.225 ;
        RECT 34.075 163.195 34.245 163.395 ;
        RECT 34.415 163.535 34.585 163.735 ;
        RECT 34.755 163.705 35.415 163.905 ;
        RECT 34.415 163.365 35.075 163.535 ;
        RECT 34.075 163.025 34.675 163.195 ;
        RECT 34.905 162.945 35.075 163.365 ;
        RECT 32.365 162.230 32.830 162.775 ;
        RECT 33.335 162.035 33.505 162.855 ;
        RECT 33.675 162.775 34.585 162.855 ;
        RECT 35.245 162.775 35.415 163.705 ;
        RECT 35.585 163.495 37.255 164.585 ;
        RECT 33.675 162.685 34.925 162.775 ;
        RECT 33.675 162.205 34.005 162.685 ;
        RECT 34.415 162.605 34.925 162.685 ;
        RECT 34.175 162.035 34.525 162.425 ;
        RECT 34.695 162.205 34.925 162.605 ;
        RECT 35.095 162.295 35.415 162.775 ;
        RECT 35.585 162.805 36.335 163.325 ;
        RECT 36.505 162.975 37.255 163.495 ;
        RECT 37.885 164.155 38.225 164.415 ;
        RECT 35.585 162.035 37.255 162.805 ;
        RECT 37.885 162.755 38.145 164.155 ;
        RECT 38.395 163.785 38.725 164.585 ;
        RECT 39.190 163.615 39.440 164.415 ;
        RECT 39.625 163.865 39.955 164.585 ;
        RECT 40.175 163.615 40.425 164.415 ;
        RECT 40.595 164.205 40.930 164.585 ;
        RECT 38.335 163.445 40.525 163.615 ;
        RECT 38.335 163.275 38.650 163.445 ;
        RECT 38.320 163.025 38.650 163.275 ;
        RECT 37.885 162.245 38.225 162.755 ;
        RECT 38.395 162.035 38.665 162.835 ;
        RECT 38.845 162.305 39.125 163.275 ;
        RECT 39.305 162.305 39.605 163.275 ;
        RECT 39.785 162.310 40.135 163.275 ;
        RECT 40.355 162.535 40.525 163.445 ;
        RECT 40.695 162.715 40.935 164.025 ;
        RECT 41.650 163.965 41.825 164.415 ;
        RECT 41.995 164.145 42.325 164.585 ;
        RECT 42.630 163.995 42.800 164.415 ;
        RECT 43.035 164.175 43.705 164.585 ;
        RECT 43.920 163.995 44.090 164.415 ;
        RECT 44.290 164.175 44.620 164.585 ;
        RECT 41.650 163.795 42.280 163.965 ;
        RECT 41.565 162.945 41.930 163.625 ;
        RECT 42.110 163.275 42.280 163.795 ;
        RECT 42.630 163.825 44.645 163.995 ;
        RECT 42.110 162.945 42.460 163.275 ;
        RECT 42.110 162.775 42.280 162.945 ;
        RECT 41.650 162.605 42.280 162.775 ;
        RECT 40.355 162.205 40.850 162.535 ;
        RECT 41.650 162.205 41.825 162.605 ;
        RECT 42.630 162.535 42.800 163.825 ;
        RECT 41.995 162.035 42.325 162.415 ;
        RECT 42.570 162.205 42.800 162.535 ;
        RECT 43.000 162.370 43.280 163.645 ;
        RECT 43.505 162.545 43.775 163.645 ;
        RECT 43.965 162.615 44.305 163.645 ;
        RECT 44.475 163.275 44.645 163.825 ;
        RECT 44.815 163.445 45.075 164.415 ;
        RECT 45.245 163.495 46.455 164.585 ;
        RECT 46.625 164.075 46.925 164.585 ;
        RECT 47.095 163.905 47.425 164.415 ;
        RECT 47.595 164.075 48.225 164.585 ;
        RECT 48.805 164.075 49.185 164.245 ;
        RECT 49.355 164.075 49.655 164.585 ;
        RECT 49.015 163.905 49.185 164.075 ;
        RECT 44.475 162.945 44.735 163.275 ;
        RECT 44.905 162.755 45.075 163.445 ;
        RECT 43.465 162.375 43.775 162.545 ;
        RECT 43.505 162.370 43.775 162.375 ;
        RECT 44.235 162.035 44.565 162.415 ;
        RECT 44.735 162.290 45.075 162.755 ;
        RECT 45.245 162.785 45.765 163.325 ;
        RECT 45.935 162.955 46.455 163.495 ;
        RECT 46.625 163.735 48.845 163.905 ;
        RECT 44.735 162.245 45.070 162.290 ;
        RECT 45.245 162.035 46.455 162.785 ;
        RECT 46.625 162.775 46.795 163.735 ;
        RECT 46.965 163.395 48.505 163.565 ;
        RECT 46.965 162.945 47.210 163.395 ;
        RECT 47.470 163.025 48.165 163.225 ;
        RECT 48.335 163.195 48.505 163.395 ;
        RECT 48.675 163.535 48.845 163.735 ;
        RECT 49.015 163.705 49.675 163.905 ;
        RECT 48.675 163.365 49.335 163.535 ;
        RECT 48.335 163.025 48.935 163.195 ;
        RECT 49.165 162.945 49.335 163.365 ;
        RECT 46.625 162.230 47.090 162.775 ;
        RECT 47.595 162.035 47.765 162.855 ;
        RECT 47.935 162.775 48.845 162.855 ;
        RECT 49.505 162.775 49.675 163.705 ;
        RECT 49.845 163.420 50.135 164.585 ;
        RECT 50.305 163.495 51.515 164.585 ;
        RECT 51.985 163.945 52.315 164.375 ;
        RECT 47.935 162.685 49.185 162.775 ;
        RECT 47.935 162.205 48.265 162.685 ;
        RECT 48.675 162.605 49.185 162.685 ;
        RECT 48.435 162.035 48.785 162.425 ;
        RECT 48.955 162.205 49.185 162.605 ;
        RECT 49.355 162.295 49.675 162.775 ;
        RECT 50.305 162.785 50.825 163.325 ;
        RECT 50.995 162.955 51.515 163.495 ;
        RECT 51.860 163.775 52.315 163.945 ;
        RECT 52.495 163.945 52.745 164.365 ;
        RECT 52.975 164.115 53.305 164.585 ;
        RECT 53.535 163.945 53.785 164.365 ;
        RECT 52.495 163.775 53.785 163.945 ;
        RECT 49.845 162.035 50.135 162.760 ;
        RECT 50.305 162.035 51.515 162.785 ;
        RECT 51.860 162.775 52.030 163.775 ;
        RECT 52.200 162.945 52.445 163.605 ;
        RECT 52.660 162.945 52.925 163.605 ;
        RECT 53.120 162.945 53.405 163.605 ;
        RECT 53.580 163.275 53.795 163.605 ;
        RECT 53.975 163.445 54.225 164.585 ;
        RECT 54.395 163.525 54.725 164.375 ;
        RECT 53.580 162.945 53.885 163.275 ;
        RECT 54.055 162.945 54.365 163.275 ;
        RECT 54.055 162.775 54.225 162.945 ;
        RECT 51.860 162.605 54.225 162.775 ;
        RECT 54.535 162.760 54.725 163.525 ;
        RECT 54.910 164.195 55.245 164.415 ;
        RECT 56.250 164.205 56.605 164.585 ;
        RECT 54.910 163.575 55.165 164.195 ;
        RECT 55.415 164.035 55.645 164.075 ;
        RECT 56.775 164.035 57.025 164.415 ;
        RECT 55.415 163.835 57.025 164.035 ;
        RECT 55.415 163.745 55.600 163.835 ;
        RECT 56.190 163.825 57.025 163.835 ;
        RECT 57.275 163.805 57.525 164.585 ;
        RECT 57.695 163.735 57.955 164.415 ;
        RECT 58.125 164.150 63.470 164.585 ;
        RECT 55.755 163.635 56.085 163.665 ;
        RECT 55.755 163.575 57.555 163.635 ;
        RECT 54.910 163.465 57.615 163.575 ;
        RECT 54.910 163.405 56.085 163.465 ;
        RECT 57.415 163.430 57.615 163.465 ;
        RECT 54.905 163.025 55.395 163.225 ;
        RECT 55.585 163.025 56.060 163.235 ;
        RECT 52.015 162.035 52.345 162.435 ;
        RECT 52.515 162.265 52.845 162.605 ;
        RECT 53.895 162.035 54.225 162.435 ;
        RECT 54.395 162.250 54.725 162.760 ;
        RECT 54.910 162.035 55.365 162.800 ;
        RECT 55.840 162.625 56.060 163.025 ;
        RECT 56.305 163.025 56.635 163.235 ;
        RECT 56.305 162.625 56.515 163.025 ;
        RECT 56.805 162.990 57.215 163.295 ;
        RECT 57.445 162.855 57.615 163.430 ;
        RECT 57.345 162.735 57.615 162.855 ;
        RECT 56.770 162.690 57.615 162.735 ;
        RECT 56.770 162.565 57.525 162.690 ;
        RECT 56.770 162.415 56.940 162.565 ;
        RECT 57.785 162.545 57.955 163.735 ;
        RECT 59.710 162.580 60.050 163.410 ;
        RECT 61.530 162.900 61.880 164.150 ;
        RECT 63.645 163.495 66.235 164.585 ;
        RECT 66.865 164.075 67.125 164.585 ;
        RECT 63.645 162.805 64.855 163.325 ;
        RECT 65.025 162.975 66.235 163.495 ;
        RECT 66.865 163.025 67.205 163.905 ;
        RECT 67.375 163.195 67.545 164.415 ;
        RECT 67.785 164.080 68.400 164.585 ;
        RECT 67.785 163.545 68.035 163.910 ;
        RECT 68.205 163.905 68.400 164.080 ;
        RECT 68.570 164.075 69.045 164.415 ;
        RECT 69.215 164.040 69.430 164.585 ;
        RECT 68.205 163.715 68.535 163.905 ;
        RECT 68.755 163.545 69.470 163.840 ;
        RECT 69.640 163.715 69.915 164.415 ;
        RECT 67.785 163.375 69.575 163.545 ;
        RECT 67.375 162.945 68.170 163.195 ;
        RECT 67.375 162.855 67.625 162.945 ;
        RECT 57.725 162.535 57.955 162.545 ;
        RECT 55.640 162.205 56.940 162.415 ;
        RECT 57.195 162.035 57.525 162.395 ;
        RECT 57.695 162.205 57.955 162.535 ;
        RECT 58.125 162.035 63.470 162.580 ;
        RECT 63.645 162.035 66.235 162.805 ;
        RECT 66.865 162.035 67.125 162.855 ;
        RECT 67.295 162.435 67.625 162.855 ;
        RECT 68.340 162.520 68.595 163.375 ;
        RECT 67.805 162.255 68.595 162.520 ;
        RECT 68.765 162.675 69.175 163.195 ;
        RECT 69.345 162.945 69.575 163.375 ;
        RECT 69.745 162.685 69.915 163.715 ;
        RECT 68.765 162.255 68.965 162.675 ;
        RECT 69.155 162.035 69.485 162.495 ;
        RECT 69.655 162.205 69.915 162.685 ;
        RECT 70.120 163.795 70.655 164.415 ;
        RECT 70.120 162.775 70.435 163.795 ;
        RECT 70.825 163.785 71.155 164.585 ;
        RECT 73.305 164.030 73.910 164.585 ;
        RECT 74.085 164.075 74.565 164.415 ;
        RECT 74.735 164.040 74.990 164.585 ;
        RECT 73.305 163.930 73.920 164.030 ;
        RECT 73.735 163.905 73.920 163.930 ;
        RECT 71.640 163.615 72.030 163.790 ;
        RECT 70.605 163.445 72.030 163.615 ;
        RECT 70.605 162.945 70.775 163.445 ;
        RECT 70.120 162.205 70.735 162.775 ;
        RECT 71.025 162.715 71.290 163.275 ;
        RECT 71.460 162.545 71.630 163.445 ;
        RECT 73.305 163.310 73.565 163.760 ;
        RECT 73.735 163.660 74.065 163.905 ;
        RECT 74.235 163.585 74.990 163.835 ;
        RECT 75.160 163.715 75.435 164.415 ;
        RECT 74.220 163.550 74.990 163.585 ;
        RECT 74.205 163.540 74.990 163.550 ;
        RECT 74.200 163.525 75.095 163.540 ;
        RECT 74.180 163.510 75.095 163.525 ;
        RECT 74.160 163.500 75.095 163.510 ;
        RECT 74.135 163.490 75.095 163.500 ;
        RECT 74.065 163.460 75.095 163.490 ;
        RECT 74.045 163.430 75.095 163.460 ;
        RECT 74.025 163.400 75.095 163.430 ;
        RECT 73.995 163.375 75.095 163.400 ;
        RECT 73.960 163.340 75.095 163.375 ;
        RECT 73.930 163.335 75.095 163.340 ;
        RECT 73.930 163.330 74.320 163.335 ;
        RECT 73.930 163.320 74.295 163.330 ;
        RECT 73.930 163.315 74.280 163.320 ;
        RECT 73.930 163.310 74.265 163.315 ;
        RECT 73.305 163.305 74.265 163.310 ;
        RECT 73.305 163.295 74.255 163.305 ;
        RECT 73.305 163.290 74.245 163.295 ;
        RECT 73.305 163.280 74.235 163.290 ;
        RECT 71.800 162.715 72.155 163.275 ;
        RECT 73.305 163.270 74.230 163.280 ;
        RECT 73.305 163.265 74.225 163.270 ;
        RECT 73.305 163.250 74.215 163.265 ;
        RECT 73.305 163.235 74.210 163.250 ;
        RECT 73.305 163.210 74.200 163.235 ;
        RECT 73.305 163.140 74.195 163.210 ;
        RECT 73.305 162.585 73.855 162.970 ;
        RECT 70.905 162.035 71.120 162.545 ;
        RECT 71.350 162.215 71.630 162.545 ;
        RECT 71.810 162.035 72.050 162.545 ;
        RECT 74.025 162.415 74.195 163.140 ;
        RECT 73.305 162.245 74.195 162.415 ;
        RECT 74.365 162.740 74.695 163.165 ;
        RECT 74.865 162.940 75.095 163.335 ;
        RECT 74.365 162.255 74.585 162.740 ;
        RECT 75.265 162.685 75.435 163.715 ;
        RECT 75.605 163.420 75.895 164.585 ;
        RECT 76.075 163.775 76.370 164.585 ;
        RECT 76.550 163.275 76.795 164.415 ;
        RECT 76.970 163.775 77.230 164.585 ;
        RECT 77.830 164.580 84.105 164.585 ;
        RECT 77.410 163.275 77.660 164.410 ;
        RECT 77.830 163.785 78.090 164.580 ;
        RECT 78.260 163.685 78.520 164.410 ;
        RECT 78.690 163.855 78.950 164.580 ;
        RECT 79.120 163.685 79.380 164.410 ;
        RECT 79.550 163.855 79.810 164.580 ;
        RECT 79.980 163.685 80.240 164.410 ;
        RECT 80.410 163.855 80.670 164.580 ;
        RECT 80.840 163.685 81.100 164.410 ;
        RECT 81.270 163.855 81.515 164.580 ;
        RECT 81.685 163.685 81.945 164.410 ;
        RECT 82.130 163.855 82.375 164.580 ;
        RECT 82.545 163.685 82.805 164.410 ;
        RECT 82.990 163.855 83.235 164.580 ;
        RECT 83.405 163.685 83.665 164.410 ;
        RECT 83.850 163.855 84.105 164.580 ;
        RECT 78.260 163.670 83.665 163.685 ;
        RECT 84.275 163.670 84.565 164.410 ;
        RECT 84.735 163.840 85.005 164.585 ;
        RECT 78.260 163.445 85.005 163.670 ;
        RECT 85.325 163.525 85.655 164.370 ;
        RECT 85.825 163.575 85.995 164.585 ;
        RECT 86.165 163.855 86.505 164.415 ;
        RECT 86.735 164.085 87.050 164.585 ;
        RECT 87.230 164.115 88.115 164.285 ;
        RECT 74.755 162.035 75.005 162.575 ;
        RECT 75.175 162.205 75.435 162.685 ;
        RECT 75.605 162.035 75.895 162.760 ;
        RECT 76.065 162.715 76.380 163.275 ;
        RECT 76.550 163.025 83.670 163.275 ;
        RECT 76.065 162.035 76.370 162.545 ;
        RECT 76.550 162.215 76.800 163.025 ;
        RECT 76.970 162.035 77.230 162.560 ;
        RECT 77.410 162.215 77.660 163.025 ;
        RECT 83.840 162.855 85.005 163.445 ;
        RECT 78.260 162.685 85.005 162.855 ;
        RECT 85.265 163.445 85.655 163.525 ;
        RECT 86.165 163.480 87.060 163.855 ;
        RECT 85.265 163.395 85.480 163.445 ;
        RECT 85.265 162.815 85.435 163.395 ;
        RECT 86.165 163.275 86.355 163.480 ;
        RECT 87.230 163.275 87.400 164.115 ;
        RECT 88.340 164.085 88.590 164.415 ;
        RECT 85.605 162.945 86.355 163.275 ;
        RECT 86.525 162.945 87.400 163.275 ;
        RECT 85.265 162.775 85.490 162.815 ;
        RECT 86.155 162.775 86.355 162.945 ;
        RECT 85.265 162.690 85.645 162.775 ;
        RECT 77.830 162.035 78.090 162.595 ;
        RECT 78.260 162.230 78.520 162.685 ;
        RECT 78.690 162.035 78.950 162.515 ;
        RECT 79.120 162.230 79.380 162.685 ;
        RECT 79.550 162.035 79.810 162.515 ;
        RECT 79.980 162.230 80.240 162.685 ;
        RECT 80.410 162.035 80.655 162.515 ;
        RECT 80.825 162.230 81.100 162.685 ;
        RECT 81.270 162.035 81.515 162.515 ;
        RECT 81.685 162.230 81.945 162.685 ;
        RECT 82.125 162.035 82.375 162.515 ;
        RECT 82.545 162.230 82.805 162.685 ;
        RECT 82.985 162.035 83.235 162.515 ;
        RECT 83.405 162.230 83.665 162.685 ;
        RECT 83.845 162.035 84.105 162.515 ;
        RECT 84.275 162.230 84.535 162.685 ;
        RECT 84.705 162.035 85.005 162.515 ;
        RECT 85.315 162.255 85.645 162.690 ;
        RECT 85.815 162.035 85.985 162.645 ;
        RECT 86.155 162.250 86.485 162.775 ;
        RECT 86.745 162.035 86.955 162.565 ;
        RECT 87.230 162.485 87.400 162.945 ;
        RECT 87.570 162.985 87.890 163.945 ;
        RECT 88.060 163.195 88.250 163.915 ;
        RECT 88.420 163.015 88.590 164.085 ;
        RECT 88.760 163.785 88.930 164.585 ;
        RECT 89.100 164.140 90.205 164.310 ;
        RECT 89.100 163.525 89.270 164.140 ;
        RECT 90.415 163.990 90.665 164.415 ;
        RECT 90.835 164.125 91.100 164.585 ;
        RECT 89.440 163.605 89.970 163.970 ;
        RECT 90.415 163.860 90.720 163.990 ;
        RECT 88.760 163.435 89.270 163.525 ;
        RECT 88.760 163.265 89.630 163.435 ;
        RECT 88.760 163.195 88.930 163.265 ;
        RECT 89.050 163.015 89.250 163.045 ;
        RECT 87.570 162.655 88.035 162.985 ;
        RECT 88.420 162.715 89.250 163.015 ;
        RECT 88.420 162.485 88.590 162.715 ;
        RECT 87.230 162.315 88.015 162.485 ;
        RECT 88.185 162.315 88.590 162.485 ;
        RECT 88.770 162.035 89.140 162.535 ;
        RECT 89.460 162.485 89.630 163.265 ;
        RECT 89.800 162.905 89.970 163.605 ;
        RECT 90.140 163.075 90.380 163.670 ;
        RECT 89.800 162.685 90.325 162.905 ;
        RECT 90.550 162.755 90.720 163.860 ;
        RECT 90.495 162.625 90.720 162.755 ;
        RECT 90.890 162.665 91.170 163.615 ;
        RECT 90.495 162.485 90.665 162.625 ;
        RECT 89.460 162.315 90.135 162.485 ;
        RECT 90.330 162.315 90.665 162.485 ;
        RECT 90.835 162.035 91.085 162.495 ;
        RECT 91.340 162.295 91.525 164.415 ;
        RECT 91.695 164.085 92.025 164.585 ;
        RECT 92.195 163.915 92.365 164.415 ;
        RECT 91.700 163.745 92.365 163.915 ;
        RECT 92.660 163.795 93.195 164.415 ;
        RECT 91.700 162.755 91.930 163.745 ;
        RECT 92.100 162.925 92.450 163.575 ;
        RECT 92.660 162.775 92.975 163.795 ;
        RECT 93.365 163.785 93.695 164.585 ;
        RECT 94.180 163.615 94.570 163.790 ;
        RECT 93.145 163.445 94.570 163.615 ;
        RECT 94.925 163.445 95.205 164.585 ;
        RECT 93.145 162.945 93.315 163.445 ;
        RECT 91.700 162.585 92.365 162.755 ;
        RECT 91.695 162.035 92.025 162.415 ;
        RECT 92.195 162.295 92.365 162.585 ;
        RECT 92.660 162.205 93.275 162.775 ;
        RECT 93.565 162.715 93.830 163.275 ;
        RECT 94.000 162.545 94.170 163.445 ;
        RECT 95.375 163.435 95.705 164.415 ;
        RECT 95.875 163.445 96.135 164.585 ;
        RECT 96.305 163.495 99.815 164.585 ;
        RECT 99.985 163.495 101.195 164.585 ;
        RECT 94.340 162.715 94.695 163.275 ;
        RECT 94.935 163.005 95.270 163.275 ;
        RECT 95.440 162.835 95.610 163.435 ;
        RECT 95.780 163.025 96.115 163.275 ;
        RECT 93.445 162.035 93.660 162.545 ;
        RECT 93.890 162.215 94.170 162.545 ;
        RECT 94.350 162.035 94.590 162.545 ;
        RECT 94.925 162.035 95.235 162.835 ;
        RECT 95.440 162.205 96.135 162.835 ;
        RECT 96.305 162.805 97.955 163.325 ;
        RECT 98.125 162.975 99.815 163.495 ;
        RECT 96.305 162.035 99.815 162.805 ;
        RECT 99.985 162.785 100.505 163.325 ;
        RECT 100.675 162.955 101.195 163.495 ;
        RECT 101.365 163.420 101.655 164.585 ;
        RECT 101.825 163.495 105.335 164.585 ;
        RECT 101.825 162.805 103.475 163.325 ;
        RECT 103.645 162.975 105.335 163.495 ;
        RECT 105.975 163.445 106.305 164.585 ;
        RECT 106.835 163.615 107.165 164.400 ;
        RECT 107.345 164.150 112.690 164.585 ;
        RECT 112.865 164.150 118.210 164.585 ;
        RECT 118.385 164.150 123.730 164.585 ;
        RECT 106.485 163.445 107.165 163.615 ;
        RECT 105.965 163.025 106.315 163.275 ;
        RECT 106.485 162.845 106.655 163.445 ;
        RECT 106.825 163.025 107.175 163.275 ;
        RECT 99.985 162.035 101.195 162.785 ;
        RECT 101.365 162.035 101.655 162.760 ;
        RECT 101.825 162.035 105.335 162.805 ;
        RECT 105.975 162.035 106.245 162.845 ;
        RECT 106.415 162.205 106.745 162.845 ;
        RECT 106.915 162.035 107.155 162.845 ;
        RECT 108.930 162.580 109.270 163.410 ;
        RECT 110.750 162.900 111.100 164.150 ;
        RECT 114.450 162.580 114.790 163.410 ;
        RECT 116.270 162.900 116.620 164.150 ;
        RECT 119.970 162.580 120.310 163.410 ;
        RECT 121.790 162.900 122.140 164.150 ;
        RECT 123.905 163.495 126.495 164.585 ;
        RECT 123.905 162.805 125.115 163.325 ;
        RECT 125.285 162.975 126.495 163.495 ;
        RECT 127.125 163.420 127.415 164.585 ;
        RECT 127.585 164.150 132.930 164.585 ;
        RECT 133.105 164.150 138.450 164.585 ;
        RECT 138.625 164.150 143.970 164.585 ;
        RECT 107.345 162.035 112.690 162.580 ;
        RECT 112.865 162.035 118.210 162.580 ;
        RECT 118.385 162.035 123.730 162.580 ;
        RECT 123.905 162.035 126.495 162.805 ;
        RECT 127.125 162.035 127.415 162.760 ;
        RECT 129.170 162.580 129.510 163.410 ;
        RECT 130.990 162.900 131.340 164.150 ;
        RECT 134.690 162.580 135.030 163.410 ;
        RECT 136.510 162.900 136.860 164.150 ;
        RECT 140.210 162.580 140.550 163.410 ;
        RECT 142.030 162.900 142.380 164.150 ;
        RECT 144.145 163.495 147.655 164.585 ;
        RECT 147.825 163.495 149.035 164.585 ;
        RECT 144.145 162.805 145.795 163.325 ;
        RECT 145.965 162.975 147.655 163.495 ;
        RECT 127.585 162.035 132.930 162.580 ;
        RECT 133.105 162.035 138.450 162.580 ;
        RECT 138.625 162.035 143.970 162.580 ;
        RECT 144.145 162.035 147.655 162.805 ;
        RECT 147.825 162.785 148.345 163.325 ;
        RECT 148.515 162.955 149.035 163.495 ;
        RECT 149.205 163.495 150.415 164.585 ;
        RECT 149.205 162.955 149.725 163.495 ;
        RECT 149.895 162.785 150.415 163.325 ;
        RECT 147.825 162.035 149.035 162.785 ;
        RECT 149.205 162.035 150.415 162.785 ;
        RECT 11.120 161.865 150.500 162.035 ;
        RECT 11.205 161.115 12.415 161.865 ;
        RECT 12.585 161.320 17.930 161.865 ;
        RECT 11.205 160.575 11.725 161.115 ;
        RECT 11.895 160.405 12.415 160.945 ;
        RECT 14.170 160.490 14.510 161.320 ;
        RECT 18.105 161.095 21.615 161.865 ;
        RECT 21.785 161.115 22.995 161.865 ;
        RECT 23.255 161.315 23.425 161.605 ;
        RECT 23.595 161.485 23.925 161.865 ;
        RECT 23.255 161.145 23.920 161.315 ;
        RECT 11.205 159.315 12.415 160.405 ;
        RECT 15.990 159.750 16.340 161.000 ;
        RECT 18.105 160.575 19.755 161.095 ;
        RECT 19.925 160.405 21.615 160.925 ;
        RECT 21.785 160.575 22.305 161.115 ;
        RECT 22.475 160.405 22.995 160.945 ;
        RECT 12.585 159.315 17.930 159.750 ;
        RECT 18.105 159.315 21.615 160.405 ;
        RECT 21.785 159.315 22.995 160.405 ;
        RECT 23.170 160.325 23.520 160.975 ;
        RECT 23.690 160.155 23.920 161.145 ;
        RECT 23.255 159.985 23.920 160.155 ;
        RECT 23.255 159.485 23.425 159.985 ;
        RECT 23.595 159.315 23.925 159.815 ;
        RECT 24.095 159.485 24.280 161.605 ;
        RECT 24.535 161.405 24.785 161.865 ;
        RECT 24.955 161.415 25.290 161.585 ;
        RECT 25.485 161.415 26.160 161.585 ;
        RECT 24.955 161.275 25.125 161.415 ;
        RECT 24.450 160.285 24.730 161.235 ;
        RECT 24.900 161.145 25.125 161.275 ;
        RECT 24.900 160.040 25.070 161.145 ;
        RECT 25.295 160.995 25.820 161.215 ;
        RECT 25.240 160.230 25.480 160.825 ;
        RECT 25.650 160.295 25.820 160.995 ;
        RECT 25.990 160.635 26.160 161.415 ;
        RECT 26.480 161.365 26.850 161.865 ;
        RECT 27.030 161.415 27.435 161.585 ;
        RECT 27.605 161.415 28.390 161.585 ;
        RECT 27.030 161.185 27.200 161.415 ;
        RECT 26.370 160.885 27.200 161.185 ;
        RECT 27.585 160.915 28.050 161.245 ;
        RECT 26.370 160.855 26.570 160.885 ;
        RECT 26.690 160.635 26.860 160.705 ;
        RECT 25.990 160.465 26.860 160.635 ;
        RECT 26.350 160.375 26.860 160.465 ;
        RECT 24.900 159.910 25.205 160.040 ;
        RECT 25.650 159.930 26.180 160.295 ;
        RECT 24.520 159.315 24.785 159.775 ;
        RECT 24.955 159.485 25.205 159.910 ;
        RECT 26.350 159.760 26.520 160.375 ;
        RECT 25.415 159.590 26.520 159.760 ;
        RECT 26.690 159.315 26.860 160.115 ;
        RECT 27.030 159.815 27.200 160.885 ;
        RECT 27.370 159.985 27.560 160.705 ;
        RECT 27.730 159.955 28.050 160.915 ;
        RECT 28.220 160.955 28.390 161.415 ;
        RECT 28.665 161.335 28.875 161.865 ;
        RECT 29.135 161.125 29.465 161.650 ;
        RECT 29.635 161.255 29.805 161.865 ;
        RECT 29.975 161.210 30.305 161.645 ;
        RECT 30.475 161.350 30.645 161.865 ;
        RECT 30.985 161.320 36.330 161.865 ;
        RECT 29.975 161.125 30.355 161.210 ;
        RECT 29.265 160.955 29.465 161.125 ;
        RECT 30.130 161.085 30.355 161.125 ;
        RECT 28.220 160.625 29.095 160.955 ;
        RECT 29.265 160.625 30.015 160.955 ;
        RECT 27.030 159.485 27.280 159.815 ;
        RECT 28.220 159.785 28.390 160.625 ;
        RECT 29.265 160.420 29.455 160.625 ;
        RECT 30.185 160.505 30.355 161.085 ;
        RECT 30.140 160.455 30.355 160.505 ;
        RECT 32.570 160.490 32.910 161.320 ;
        RECT 36.965 161.140 37.255 161.865 ;
        RECT 37.425 161.125 37.740 161.500 ;
        RECT 37.995 161.125 38.165 161.865 ;
        RECT 38.415 161.295 38.585 161.500 ;
        RECT 38.810 161.465 39.185 161.865 ;
        RECT 39.355 161.295 39.525 161.645 ;
        RECT 39.710 161.465 40.040 161.865 ;
        RECT 40.210 161.295 40.380 161.645 ;
        RECT 40.550 161.465 40.930 161.865 ;
        RECT 38.415 161.125 38.915 161.295 ;
        RECT 39.355 161.125 40.950 161.295 ;
        RECT 41.120 161.190 41.395 161.535 ;
        RECT 28.560 160.045 29.455 160.420 ;
        RECT 29.965 160.375 30.355 160.455 ;
        RECT 27.505 159.615 28.390 159.785 ;
        RECT 28.570 159.315 28.885 159.815 ;
        RECT 29.115 159.485 29.455 160.045 ;
        RECT 29.625 159.315 29.795 160.325 ;
        RECT 29.965 159.530 30.295 160.375 ;
        RECT 30.465 159.315 30.635 160.230 ;
        RECT 34.390 159.750 34.740 161.000 ;
        RECT 30.985 159.315 36.330 159.750 ;
        RECT 36.965 159.315 37.255 160.480 ;
        RECT 37.425 160.085 37.595 161.125 ;
        RECT 37.765 160.255 38.115 160.955 ;
        RECT 38.285 160.625 38.575 160.955 ;
        RECT 38.745 160.875 38.915 161.125 ;
        RECT 40.780 160.955 40.950 161.125 ;
        RECT 38.745 160.705 39.170 160.875 ;
        RECT 38.745 160.425 38.915 160.705 ;
        RECT 39.565 160.535 39.735 160.955 ;
        RECT 39.955 160.625 40.610 160.955 ;
        RECT 40.780 160.625 41.055 160.955 ;
        RECT 38.330 160.255 38.915 160.425 ;
        RECT 39.085 160.365 39.735 160.535 ;
        RECT 40.780 160.455 40.950 160.625 ;
        RECT 41.225 160.455 41.395 161.190 ;
        RECT 41.565 161.095 43.235 161.865 ;
        RECT 41.565 160.575 42.315 161.095 ;
        RECT 43.925 161.045 44.135 161.865 ;
        RECT 44.305 161.065 44.635 161.695 ;
        RECT 39.085 160.085 39.255 160.365 ;
        RECT 40.290 160.285 40.950 160.455 ;
        RECT 40.290 160.165 40.460 160.285 ;
        RECT 37.425 159.915 39.255 160.085 ;
        RECT 39.425 159.995 40.460 160.165 ;
        RECT 37.425 159.495 37.685 159.915 ;
        RECT 39.425 159.745 39.595 159.995 ;
        RECT 37.855 159.315 38.185 159.745 ;
        RECT 38.850 159.575 39.595 159.745 ;
        RECT 39.785 159.655 40.460 159.825 ;
        RECT 39.820 159.495 40.460 159.655 ;
        RECT 40.630 159.315 40.910 160.115 ;
        RECT 41.120 159.485 41.395 160.455 ;
        RECT 42.485 160.405 43.235 160.925 ;
        RECT 44.305 160.465 44.555 161.065 ;
        RECT 44.805 161.045 45.035 161.865 ;
        RECT 45.245 161.095 48.755 161.865 ;
        RECT 49.845 161.365 50.185 161.865 ;
        RECT 44.725 160.625 45.055 160.875 ;
        RECT 45.245 160.575 46.895 161.095 ;
        RECT 41.565 159.315 43.235 160.405 ;
        RECT 43.925 159.315 44.135 160.455 ;
        RECT 44.305 159.485 44.635 160.465 ;
        RECT 44.805 159.315 45.035 160.455 ;
        RECT 47.065 160.405 48.755 160.925 ;
        RECT 49.845 160.625 50.185 161.195 ;
        RECT 50.355 160.955 50.600 161.645 ;
        RECT 50.795 161.365 51.125 161.865 ;
        RECT 51.325 161.295 51.495 161.645 ;
        RECT 51.670 161.465 52.000 161.865 ;
        RECT 52.170 161.295 52.340 161.645 ;
        RECT 52.510 161.465 52.890 161.865 ;
        RECT 51.325 161.125 52.910 161.295 ;
        RECT 53.080 161.190 53.355 161.535 ;
        RECT 52.740 160.955 52.910 161.125 ;
        RECT 50.355 160.625 51.010 160.955 ;
        RECT 45.245 159.315 48.755 160.405 ;
        RECT 49.845 159.315 50.185 160.390 ;
        RECT 50.355 160.030 50.595 160.625 ;
        RECT 50.790 160.165 51.110 160.455 ;
        RECT 51.280 160.335 52.020 160.955 ;
        RECT 52.190 160.625 52.570 160.955 ;
        RECT 52.740 160.625 53.015 160.955 ;
        RECT 52.740 160.455 52.910 160.625 ;
        RECT 53.185 160.455 53.355 161.190 ;
        RECT 53.525 161.095 55.195 161.865 ;
        RECT 55.415 161.210 55.745 161.645 ;
        RECT 55.915 161.255 56.085 161.865 ;
        RECT 55.365 161.125 55.745 161.210 ;
        RECT 56.255 161.125 56.585 161.650 ;
        RECT 56.845 161.335 57.055 161.865 ;
        RECT 57.330 161.415 58.115 161.585 ;
        RECT 58.285 161.415 58.690 161.585 ;
        RECT 53.525 160.575 54.275 161.095 ;
        RECT 55.365 161.085 55.590 161.125 ;
        RECT 52.250 160.285 52.910 160.455 ;
        RECT 52.250 160.165 52.420 160.285 ;
        RECT 50.790 159.995 52.420 160.165 ;
        RECT 50.370 159.535 52.420 159.825 ;
        RECT 52.590 159.315 52.870 160.115 ;
        RECT 53.080 159.485 53.355 160.455 ;
        RECT 54.445 160.405 55.195 160.925 ;
        RECT 53.525 159.315 55.195 160.405 ;
        RECT 55.365 160.505 55.535 161.085 ;
        RECT 56.255 160.955 56.455 161.125 ;
        RECT 57.330 160.955 57.500 161.415 ;
        RECT 55.705 160.625 56.455 160.955 ;
        RECT 56.625 160.625 57.500 160.955 ;
        RECT 55.365 160.455 55.580 160.505 ;
        RECT 55.365 160.375 55.755 160.455 ;
        RECT 55.425 159.530 55.755 160.375 ;
        RECT 56.265 160.420 56.455 160.625 ;
        RECT 55.925 159.315 56.095 160.325 ;
        RECT 56.265 160.045 57.160 160.420 ;
        RECT 56.265 159.485 56.605 160.045 ;
        RECT 56.835 159.315 57.150 159.815 ;
        RECT 57.330 159.785 57.500 160.625 ;
        RECT 57.670 160.915 58.135 161.245 ;
        RECT 58.520 161.185 58.690 161.415 ;
        RECT 58.870 161.365 59.240 161.865 ;
        RECT 59.560 161.415 60.235 161.585 ;
        RECT 60.430 161.415 60.765 161.585 ;
        RECT 57.670 159.955 57.990 160.915 ;
        RECT 58.520 160.885 59.350 161.185 ;
        RECT 58.160 159.985 58.350 160.705 ;
        RECT 58.520 159.815 58.690 160.885 ;
        RECT 59.150 160.855 59.350 160.885 ;
        RECT 58.860 160.635 59.030 160.705 ;
        RECT 59.560 160.635 59.730 161.415 ;
        RECT 60.595 161.275 60.765 161.415 ;
        RECT 60.935 161.405 61.185 161.865 ;
        RECT 58.860 160.465 59.730 160.635 ;
        RECT 59.900 160.995 60.425 161.215 ;
        RECT 60.595 161.145 60.820 161.275 ;
        RECT 58.860 160.375 59.370 160.465 ;
        RECT 57.330 159.615 58.215 159.785 ;
        RECT 58.440 159.485 58.690 159.815 ;
        RECT 58.860 159.315 59.030 160.115 ;
        RECT 59.200 159.760 59.370 160.375 ;
        RECT 59.900 160.295 60.070 160.995 ;
        RECT 59.540 159.930 60.070 160.295 ;
        RECT 60.240 160.230 60.480 160.825 ;
        RECT 60.650 160.040 60.820 161.145 ;
        RECT 60.990 160.285 61.270 161.235 ;
        RECT 60.515 159.910 60.820 160.040 ;
        RECT 59.200 159.590 60.305 159.760 ;
        RECT 60.515 159.485 60.765 159.910 ;
        RECT 60.935 159.315 61.200 159.775 ;
        RECT 61.440 159.485 61.625 161.605 ;
        RECT 61.795 161.485 62.125 161.865 ;
        RECT 62.295 161.315 62.465 161.605 ;
        RECT 61.800 161.145 62.465 161.315 ;
        RECT 61.800 160.155 62.030 161.145 ;
        RECT 62.725 161.140 63.015 161.865 ;
        RECT 63.185 161.190 63.445 161.695 ;
        RECT 63.625 161.485 63.955 161.865 ;
        RECT 64.135 161.315 64.305 161.695 ;
        RECT 62.200 160.325 62.550 160.975 ;
        RECT 61.800 159.985 62.465 160.155 ;
        RECT 61.795 159.315 62.125 159.815 ;
        RECT 62.295 159.485 62.465 159.985 ;
        RECT 62.725 159.315 63.015 160.480 ;
        RECT 63.185 160.390 63.355 161.190 ;
        RECT 63.640 161.145 64.305 161.315 ;
        RECT 63.640 160.890 63.810 161.145 ;
        RECT 64.565 161.115 65.775 161.865 ;
        RECT 65.945 161.125 66.305 161.500 ;
        RECT 66.570 161.125 66.740 161.865 ;
        RECT 67.020 161.295 67.190 161.500 ;
        RECT 67.020 161.125 67.560 161.295 ;
        RECT 63.525 160.560 63.810 160.890 ;
        RECT 64.045 160.595 64.375 160.965 ;
        RECT 64.565 160.575 65.085 161.115 ;
        RECT 63.640 160.415 63.810 160.560 ;
        RECT 63.185 159.485 63.455 160.390 ;
        RECT 63.640 160.245 64.305 160.415 ;
        RECT 65.255 160.405 65.775 160.945 ;
        RECT 63.625 159.315 63.955 160.075 ;
        RECT 64.135 159.485 64.305 160.245 ;
        RECT 64.565 159.315 65.775 160.405 ;
        RECT 65.945 160.470 66.200 161.125 ;
        RECT 66.370 160.625 66.720 160.955 ;
        RECT 66.890 160.625 67.220 160.955 ;
        RECT 65.945 159.485 66.285 160.470 ;
        RECT 66.455 160.085 66.720 160.625 ;
        RECT 67.390 160.425 67.560 161.125 ;
        RECT 66.935 160.255 67.560 160.425 ;
        RECT 67.730 160.495 67.900 161.695 ;
        RECT 68.130 161.215 68.460 161.695 ;
        RECT 68.630 161.395 68.800 161.865 ;
        RECT 68.970 161.215 69.300 161.680 ;
        RECT 68.130 161.045 69.300 161.215 ;
        RECT 70.085 161.125 70.470 161.695 ;
        RECT 70.640 161.405 70.965 161.865 ;
        RECT 71.485 161.235 71.765 161.695 ;
        RECT 68.070 160.665 68.640 160.875 ;
        RECT 68.810 160.665 69.455 160.875 ;
        RECT 67.730 160.085 68.435 160.495 ;
        RECT 70.085 160.455 70.365 161.125 ;
        RECT 70.640 161.065 71.765 161.235 ;
        RECT 70.640 160.955 71.090 161.065 ;
        RECT 70.535 160.625 71.090 160.955 ;
        RECT 71.955 160.895 72.355 161.695 ;
        RECT 72.755 161.405 73.025 161.865 ;
        RECT 73.195 161.235 73.480 161.695 ;
        RECT 66.455 159.915 68.435 160.085 ;
        RECT 66.455 159.315 66.865 159.745 ;
        RECT 67.610 159.315 67.940 159.735 ;
        RECT 68.110 159.485 68.435 159.915 ;
        RECT 68.910 159.315 69.240 160.415 ;
        RECT 70.085 159.485 70.470 160.455 ;
        RECT 70.640 160.165 71.090 160.625 ;
        RECT 71.260 160.335 72.355 160.895 ;
        RECT 70.640 159.945 71.765 160.165 ;
        RECT 70.640 159.315 70.965 159.775 ;
        RECT 71.485 159.485 71.765 159.945 ;
        RECT 71.955 159.485 72.355 160.335 ;
        RECT 72.525 161.065 73.480 161.235 ;
        RECT 73.775 161.140 74.105 161.650 ;
        RECT 74.275 161.465 74.605 161.865 ;
        RECT 75.655 161.295 75.985 161.635 ;
        RECT 76.155 161.465 76.485 161.865 ;
        RECT 72.525 160.165 72.735 161.065 ;
        RECT 72.905 160.335 73.595 160.895 ;
        RECT 73.775 160.375 73.965 161.140 ;
        RECT 74.275 161.125 76.640 161.295 ;
        RECT 74.275 160.955 74.445 161.125 ;
        RECT 74.135 160.625 74.445 160.955 ;
        RECT 74.615 160.625 74.920 160.955 ;
        RECT 72.525 159.945 73.480 160.165 ;
        RECT 72.755 159.315 73.025 159.775 ;
        RECT 73.195 159.485 73.480 159.945 ;
        RECT 73.775 159.525 74.105 160.375 ;
        RECT 74.275 159.315 74.525 160.455 ;
        RECT 74.705 160.295 74.920 160.625 ;
        RECT 75.095 160.295 75.380 160.955 ;
        RECT 75.575 160.295 75.840 160.955 ;
        RECT 76.055 160.295 76.300 160.955 ;
        RECT 76.470 160.125 76.640 161.125 ;
        RECT 76.985 161.045 77.245 161.865 ;
        RECT 77.415 161.045 77.745 161.465 ;
        RECT 77.925 161.380 78.715 161.645 ;
        RECT 77.495 160.955 77.745 161.045 ;
        RECT 74.715 159.955 76.005 160.125 ;
        RECT 74.715 159.535 74.965 159.955 ;
        RECT 75.195 159.315 75.525 159.785 ;
        RECT 75.755 159.535 76.005 159.955 ;
        RECT 76.185 159.955 76.640 160.125 ;
        RECT 76.985 159.995 77.325 160.875 ;
        RECT 77.495 160.705 78.290 160.955 ;
        RECT 76.185 159.525 76.515 159.955 ;
        RECT 76.985 159.315 77.245 159.825 ;
        RECT 77.495 159.485 77.665 160.705 ;
        RECT 78.460 160.525 78.715 161.380 ;
        RECT 78.885 161.225 79.085 161.645 ;
        RECT 79.275 161.405 79.605 161.865 ;
        RECT 78.885 160.705 79.295 161.225 ;
        RECT 79.775 161.215 80.035 161.695 ;
        RECT 79.465 160.525 79.695 160.955 ;
        RECT 77.905 160.355 79.695 160.525 ;
        RECT 77.905 159.990 78.155 160.355 ;
        RECT 78.325 159.995 78.655 160.185 ;
        RECT 78.875 160.060 79.590 160.355 ;
        RECT 79.865 160.185 80.035 161.215 ;
        RECT 78.325 159.820 78.520 159.995 ;
        RECT 77.905 159.315 78.520 159.820 ;
        RECT 78.690 159.485 79.165 159.825 ;
        RECT 79.335 159.315 79.550 159.860 ;
        RECT 79.760 159.485 80.035 160.185 ;
        RECT 80.215 161.140 80.545 161.650 ;
        RECT 80.715 161.465 81.045 161.865 ;
        RECT 82.095 161.295 82.425 161.635 ;
        RECT 82.595 161.465 82.925 161.865 ;
        RECT 83.515 161.315 83.685 161.695 ;
        RECT 83.865 161.485 84.195 161.865 ;
        RECT 80.215 160.375 80.405 161.140 ;
        RECT 80.715 161.125 83.080 161.295 ;
        RECT 83.515 161.145 84.180 161.315 ;
        RECT 84.375 161.190 84.635 161.695 ;
        RECT 80.715 160.955 80.885 161.125 ;
        RECT 80.575 160.625 80.885 160.955 ;
        RECT 81.055 160.625 81.360 160.955 ;
        RECT 80.215 159.525 80.545 160.375 ;
        RECT 80.715 159.315 80.965 160.455 ;
        RECT 81.145 160.295 81.360 160.625 ;
        RECT 81.535 160.295 81.820 160.955 ;
        RECT 82.015 160.295 82.280 160.955 ;
        RECT 82.495 160.295 82.740 160.955 ;
        RECT 82.910 160.125 83.080 161.125 ;
        RECT 83.445 160.595 83.775 160.965 ;
        RECT 84.010 160.890 84.180 161.145 ;
        RECT 84.010 160.560 84.295 160.890 ;
        RECT 84.010 160.415 84.180 160.560 ;
        RECT 81.155 159.955 82.445 160.125 ;
        RECT 81.155 159.535 81.405 159.955 ;
        RECT 81.635 159.315 81.965 159.785 ;
        RECT 82.195 159.535 82.445 159.955 ;
        RECT 82.625 159.955 83.080 160.125 ;
        RECT 83.515 160.245 84.180 160.415 ;
        RECT 84.465 160.390 84.635 161.190 ;
        RECT 84.805 161.095 88.315 161.865 ;
        RECT 88.485 161.140 88.775 161.865 ;
        RECT 88.945 161.125 89.330 161.695 ;
        RECT 89.500 161.405 89.825 161.865 ;
        RECT 90.345 161.235 90.625 161.695 ;
        RECT 84.805 160.575 86.455 161.095 ;
        RECT 86.625 160.405 88.315 160.925 ;
        RECT 82.625 159.525 82.955 159.955 ;
        RECT 83.515 159.485 83.685 160.245 ;
        RECT 83.865 159.315 84.195 160.075 ;
        RECT 84.365 159.485 84.635 160.390 ;
        RECT 84.805 159.315 88.315 160.405 ;
        RECT 88.485 159.315 88.775 160.480 ;
        RECT 88.945 160.455 89.225 161.125 ;
        RECT 89.500 161.065 90.625 161.235 ;
        RECT 89.500 160.955 89.950 161.065 ;
        RECT 89.395 160.625 89.950 160.955 ;
        RECT 90.815 160.895 91.215 161.695 ;
        RECT 91.615 161.405 91.885 161.865 ;
        RECT 92.055 161.235 92.340 161.695 ;
        RECT 88.945 159.485 89.330 160.455 ;
        RECT 89.500 160.165 89.950 160.625 ;
        RECT 90.120 160.335 91.215 160.895 ;
        RECT 89.500 159.945 90.625 160.165 ;
        RECT 89.500 159.315 89.825 159.775 ;
        RECT 90.345 159.485 90.625 159.945 ;
        RECT 90.815 159.485 91.215 160.335 ;
        RECT 91.385 161.065 92.340 161.235 ;
        RECT 92.625 161.095 96.135 161.865 ;
        RECT 96.855 161.315 97.025 161.605 ;
        RECT 97.195 161.485 97.525 161.865 ;
        RECT 96.855 161.145 97.520 161.315 ;
        RECT 91.385 160.165 91.595 161.065 ;
        RECT 91.765 160.335 92.455 160.895 ;
        RECT 92.625 160.575 94.275 161.095 ;
        RECT 94.445 160.405 96.135 160.925 ;
        RECT 91.385 159.945 92.340 160.165 ;
        RECT 91.615 159.315 91.885 159.775 ;
        RECT 92.055 159.485 92.340 159.945 ;
        RECT 92.625 159.315 96.135 160.405 ;
        RECT 96.770 160.325 97.120 160.975 ;
        RECT 97.290 160.155 97.520 161.145 ;
        RECT 96.855 159.985 97.520 160.155 ;
        RECT 96.855 159.485 97.025 159.985 ;
        RECT 97.195 159.315 97.525 159.815 ;
        RECT 97.695 159.485 97.880 161.605 ;
        RECT 98.135 161.405 98.385 161.865 ;
        RECT 98.555 161.415 98.890 161.585 ;
        RECT 99.085 161.415 99.760 161.585 ;
        RECT 98.555 161.275 98.725 161.415 ;
        RECT 98.050 160.285 98.330 161.235 ;
        RECT 98.500 161.145 98.725 161.275 ;
        RECT 98.500 160.040 98.670 161.145 ;
        RECT 98.895 160.995 99.420 161.215 ;
        RECT 98.840 160.230 99.080 160.825 ;
        RECT 99.250 160.295 99.420 160.995 ;
        RECT 99.590 160.635 99.760 161.415 ;
        RECT 100.080 161.365 100.450 161.865 ;
        RECT 100.630 161.415 101.035 161.585 ;
        RECT 101.205 161.415 101.990 161.585 ;
        RECT 100.630 161.185 100.800 161.415 ;
        RECT 99.970 160.885 100.800 161.185 ;
        RECT 101.185 160.915 101.650 161.245 ;
        RECT 99.970 160.855 100.170 160.885 ;
        RECT 100.290 160.635 100.460 160.705 ;
        RECT 99.590 160.465 100.460 160.635 ;
        RECT 99.950 160.375 100.460 160.465 ;
        RECT 98.500 159.910 98.805 160.040 ;
        RECT 99.250 159.930 99.780 160.295 ;
        RECT 98.120 159.315 98.385 159.775 ;
        RECT 98.555 159.485 98.805 159.910 ;
        RECT 99.950 159.760 100.120 160.375 ;
        RECT 99.015 159.590 100.120 159.760 ;
        RECT 100.290 159.315 100.460 160.115 ;
        RECT 100.630 159.815 100.800 160.885 ;
        RECT 100.970 159.985 101.160 160.705 ;
        RECT 101.330 159.955 101.650 160.915 ;
        RECT 101.820 160.955 101.990 161.415 ;
        RECT 102.265 161.335 102.475 161.865 ;
        RECT 102.735 161.125 103.065 161.650 ;
        RECT 103.235 161.255 103.405 161.865 ;
        RECT 103.575 161.210 103.905 161.645 ;
        RECT 103.575 161.125 103.955 161.210 ;
        RECT 102.865 160.955 103.065 161.125 ;
        RECT 103.730 161.085 103.955 161.125 ;
        RECT 101.820 160.625 102.695 160.955 ;
        RECT 102.865 160.625 103.615 160.955 ;
        RECT 100.630 159.485 100.880 159.815 ;
        RECT 101.820 159.785 101.990 160.625 ;
        RECT 102.865 160.420 103.055 160.625 ;
        RECT 103.785 160.505 103.955 161.085 ;
        RECT 104.125 161.095 105.795 161.865 ;
        RECT 106.515 161.315 106.685 161.605 ;
        RECT 106.855 161.485 107.185 161.865 ;
        RECT 106.515 161.145 107.180 161.315 ;
        RECT 104.125 160.575 104.875 161.095 ;
        RECT 103.740 160.455 103.955 160.505 ;
        RECT 102.160 160.045 103.055 160.420 ;
        RECT 103.565 160.375 103.955 160.455 ;
        RECT 105.045 160.405 105.795 160.925 ;
        RECT 101.105 159.615 101.990 159.785 ;
        RECT 102.170 159.315 102.485 159.815 ;
        RECT 102.715 159.485 103.055 160.045 ;
        RECT 103.225 159.315 103.395 160.325 ;
        RECT 103.565 159.530 103.895 160.375 ;
        RECT 104.125 159.315 105.795 160.405 ;
        RECT 106.430 160.325 106.780 160.975 ;
        RECT 106.950 160.155 107.180 161.145 ;
        RECT 106.515 159.985 107.180 160.155 ;
        RECT 106.515 159.485 106.685 159.985 ;
        RECT 106.855 159.315 107.185 159.815 ;
        RECT 107.355 159.485 107.540 161.605 ;
        RECT 107.795 161.405 108.045 161.865 ;
        RECT 108.215 161.415 108.550 161.585 ;
        RECT 108.745 161.415 109.420 161.585 ;
        RECT 108.215 161.275 108.385 161.415 ;
        RECT 107.710 160.285 107.990 161.235 ;
        RECT 108.160 161.145 108.385 161.275 ;
        RECT 108.160 160.040 108.330 161.145 ;
        RECT 108.555 160.995 109.080 161.215 ;
        RECT 108.500 160.230 108.740 160.825 ;
        RECT 108.910 160.295 109.080 160.995 ;
        RECT 109.250 160.635 109.420 161.415 ;
        RECT 109.740 161.365 110.110 161.865 ;
        RECT 110.290 161.415 110.695 161.585 ;
        RECT 110.865 161.415 111.650 161.585 ;
        RECT 110.290 161.185 110.460 161.415 ;
        RECT 109.630 160.885 110.460 161.185 ;
        RECT 110.845 160.915 111.310 161.245 ;
        RECT 109.630 160.855 109.830 160.885 ;
        RECT 109.950 160.635 110.120 160.705 ;
        RECT 109.250 160.465 110.120 160.635 ;
        RECT 109.610 160.375 110.120 160.465 ;
        RECT 108.160 159.910 108.465 160.040 ;
        RECT 108.910 159.930 109.440 160.295 ;
        RECT 107.780 159.315 108.045 159.775 ;
        RECT 108.215 159.485 108.465 159.910 ;
        RECT 109.610 159.760 109.780 160.375 ;
        RECT 108.675 159.590 109.780 159.760 ;
        RECT 109.950 159.315 110.120 160.115 ;
        RECT 110.290 159.815 110.460 160.885 ;
        RECT 110.630 159.985 110.820 160.705 ;
        RECT 110.990 159.955 111.310 160.915 ;
        RECT 111.480 160.955 111.650 161.415 ;
        RECT 111.925 161.335 112.135 161.865 ;
        RECT 112.395 161.125 112.725 161.650 ;
        RECT 112.895 161.255 113.065 161.865 ;
        RECT 113.235 161.210 113.565 161.645 ;
        RECT 113.735 161.350 113.905 161.865 ;
        RECT 113.235 161.125 113.615 161.210 ;
        RECT 114.245 161.140 114.535 161.865 ;
        RECT 114.705 161.320 120.050 161.865 ;
        RECT 120.225 161.320 125.570 161.865 ;
        RECT 125.745 161.320 131.090 161.865 ;
        RECT 131.265 161.320 136.610 161.865 ;
        RECT 112.525 160.955 112.725 161.125 ;
        RECT 113.390 161.085 113.615 161.125 ;
        RECT 111.480 160.625 112.355 160.955 ;
        RECT 112.525 160.625 113.275 160.955 ;
        RECT 110.290 159.485 110.540 159.815 ;
        RECT 111.480 159.785 111.650 160.625 ;
        RECT 112.525 160.420 112.715 160.625 ;
        RECT 113.445 160.505 113.615 161.085 ;
        RECT 113.400 160.455 113.615 160.505 ;
        RECT 116.290 160.490 116.630 161.320 ;
        RECT 111.820 160.045 112.715 160.420 ;
        RECT 113.225 160.375 113.615 160.455 ;
        RECT 110.765 159.615 111.650 159.785 ;
        RECT 111.830 159.315 112.145 159.815 ;
        RECT 112.375 159.485 112.715 160.045 ;
        RECT 112.885 159.315 113.055 160.325 ;
        RECT 113.225 159.530 113.555 160.375 ;
        RECT 113.725 159.315 113.895 160.230 ;
        RECT 114.245 159.315 114.535 160.480 ;
        RECT 118.110 159.750 118.460 161.000 ;
        RECT 121.810 160.490 122.150 161.320 ;
        RECT 123.630 159.750 123.980 161.000 ;
        RECT 127.330 160.490 127.670 161.320 ;
        RECT 129.150 159.750 129.500 161.000 ;
        RECT 132.850 160.490 133.190 161.320 ;
        RECT 136.785 161.095 139.375 161.865 ;
        RECT 140.005 161.140 140.295 161.865 ;
        RECT 140.465 161.320 145.810 161.865 ;
        RECT 134.670 159.750 135.020 161.000 ;
        RECT 136.785 160.575 137.995 161.095 ;
        RECT 138.165 160.405 139.375 160.925 ;
        RECT 142.050 160.490 142.390 161.320 ;
        RECT 145.985 161.095 148.575 161.865 ;
        RECT 149.205 161.115 150.415 161.865 ;
        RECT 114.705 159.315 120.050 159.750 ;
        RECT 120.225 159.315 125.570 159.750 ;
        RECT 125.745 159.315 131.090 159.750 ;
        RECT 131.265 159.315 136.610 159.750 ;
        RECT 136.785 159.315 139.375 160.405 ;
        RECT 140.005 159.315 140.295 160.480 ;
        RECT 143.870 159.750 144.220 161.000 ;
        RECT 145.985 160.575 147.195 161.095 ;
        RECT 147.365 160.405 148.575 160.925 ;
        RECT 140.465 159.315 145.810 159.750 ;
        RECT 145.985 159.315 148.575 160.405 ;
        RECT 149.205 160.405 149.725 160.945 ;
        RECT 149.895 160.575 150.415 161.115 ;
        RECT 149.205 159.315 150.415 160.405 ;
        RECT 11.120 159.145 150.500 159.315 ;
        RECT 11.205 158.055 12.415 159.145 ;
        RECT 12.585 158.710 17.930 159.145 ;
        RECT 18.105 158.710 23.450 159.145 ;
        RECT 11.205 157.345 11.725 157.885 ;
        RECT 11.895 157.515 12.415 158.055 ;
        RECT 11.205 156.595 12.415 157.345 ;
        RECT 14.170 157.140 14.510 157.970 ;
        RECT 15.990 157.460 16.340 158.710 ;
        RECT 19.690 157.140 20.030 157.970 ;
        RECT 21.510 157.460 21.860 158.710 ;
        RECT 24.085 157.980 24.375 159.145 ;
        RECT 24.745 158.475 25.025 159.145 ;
        RECT 25.195 158.255 25.495 158.805 ;
        RECT 25.695 158.425 26.025 159.145 ;
        RECT 26.215 158.425 26.675 158.975 ;
        RECT 24.560 157.835 24.825 158.195 ;
        RECT 25.195 158.085 26.135 158.255 ;
        RECT 25.965 157.835 26.135 158.085 ;
        RECT 24.560 157.585 25.235 157.835 ;
        RECT 25.455 157.585 25.795 157.835 ;
        RECT 25.965 157.505 26.255 157.835 ;
        RECT 25.965 157.415 26.135 157.505 ;
        RECT 12.585 156.595 17.930 157.140 ;
        RECT 18.105 156.595 23.450 157.140 ;
        RECT 24.085 156.595 24.375 157.320 ;
        RECT 24.745 157.225 26.135 157.415 ;
        RECT 24.745 156.865 25.075 157.225 ;
        RECT 26.425 157.055 26.675 158.425 ;
        RECT 25.695 156.595 25.945 157.055 ;
        RECT 26.115 156.765 26.675 157.055 ;
        RECT 26.845 158.070 27.115 158.975 ;
        RECT 27.285 158.385 27.615 159.145 ;
        RECT 27.795 158.215 27.965 158.975 ;
        RECT 28.225 158.710 33.570 159.145 ;
        RECT 33.745 158.710 39.090 159.145 ;
        RECT 39.265 158.710 44.610 159.145 ;
        RECT 26.845 157.270 27.015 158.070 ;
        RECT 27.300 158.045 27.965 158.215 ;
        RECT 27.300 157.900 27.470 158.045 ;
        RECT 27.185 157.570 27.470 157.900 ;
        RECT 27.300 157.315 27.470 157.570 ;
        RECT 27.705 157.495 28.035 157.865 ;
        RECT 26.845 156.765 27.105 157.270 ;
        RECT 27.300 157.145 27.965 157.315 ;
        RECT 27.285 156.595 27.615 156.975 ;
        RECT 27.795 156.765 27.965 157.145 ;
        RECT 29.810 157.140 30.150 157.970 ;
        RECT 31.630 157.460 31.980 158.710 ;
        RECT 35.330 157.140 35.670 157.970 ;
        RECT 37.150 157.460 37.500 158.710 ;
        RECT 40.850 157.140 41.190 157.970 ;
        RECT 42.670 157.460 43.020 158.710 ;
        RECT 44.785 158.055 48.295 159.145 ;
        RECT 48.465 158.055 49.675 159.145 ;
        RECT 44.785 157.365 46.435 157.885 ;
        RECT 46.605 157.535 48.295 158.055 ;
        RECT 28.225 156.595 33.570 157.140 ;
        RECT 33.745 156.595 39.090 157.140 ;
        RECT 39.265 156.595 44.610 157.140 ;
        RECT 44.785 156.595 48.295 157.365 ;
        RECT 48.465 157.345 48.985 157.885 ;
        RECT 49.155 157.515 49.675 158.055 ;
        RECT 49.845 157.980 50.135 159.145 ;
        RECT 50.310 158.765 50.645 159.145 ;
        RECT 48.465 156.595 49.675 157.345 ;
        RECT 49.845 156.595 50.135 157.320 ;
        RECT 50.305 157.275 50.545 158.585 ;
        RECT 50.815 158.175 51.065 158.975 ;
        RECT 51.285 158.425 51.615 159.145 ;
        RECT 51.800 158.175 52.050 158.975 ;
        RECT 52.515 158.345 52.845 159.145 ;
        RECT 53.015 158.715 53.355 158.975 ;
        RECT 50.715 158.005 52.905 158.175 ;
        RECT 50.715 157.095 50.885 158.005 ;
        RECT 52.590 157.835 52.905 158.005 ;
        RECT 50.390 156.765 50.885 157.095 ;
        RECT 51.105 156.870 51.455 157.835 ;
        RECT 51.635 156.865 51.935 157.835 ;
        RECT 52.115 156.865 52.395 157.835 ;
        RECT 52.590 157.585 52.920 157.835 ;
        RECT 52.575 156.595 52.845 157.395 ;
        RECT 53.095 157.315 53.355 158.715 ;
        RECT 53.525 158.055 56.115 159.145 ;
        RECT 56.745 158.590 57.350 159.145 ;
        RECT 57.525 158.635 58.005 158.975 ;
        RECT 58.175 158.600 58.430 159.145 ;
        RECT 56.745 158.490 57.360 158.590 ;
        RECT 57.175 158.465 57.360 158.490 ;
        RECT 53.015 156.805 53.355 157.315 ;
        RECT 53.525 157.365 54.735 157.885 ;
        RECT 54.905 157.535 56.115 158.055 ;
        RECT 56.745 157.870 57.005 158.320 ;
        RECT 57.175 158.220 57.505 158.465 ;
        RECT 57.675 158.145 58.430 158.395 ;
        RECT 58.600 158.275 58.875 158.975 ;
        RECT 59.045 158.710 64.390 159.145 ;
        RECT 64.565 158.710 69.910 159.145 ;
        RECT 57.660 158.110 58.430 158.145 ;
        RECT 57.645 158.100 58.430 158.110 ;
        RECT 57.640 158.085 58.535 158.100 ;
        RECT 57.620 158.070 58.535 158.085 ;
        RECT 57.600 158.060 58.535 158.070 ;
        RECT 57.575 158.050 58.535 158.060 ;
        RECT 57.505 158.020 58.535 158.050 ;
        RECT 57.485 157.990 58.535 158.020 ;
        RECT 57.465 157.960 58.535 157.990 ;
        RECT 57.435 157.935 58.535 157.960 ;
        RECT 57.400 157.900 58.535 157.935 ;
        RECT 57.370 157.895 58.535 157.900 ;
        RECT 57.370 157.890 57.760 157.895 ;
        RECT 57.370 157.880 57.735 157.890 ;
        RECT 57.370 157.875 57.720 157.880 ;
        RECT 57.370 157.870 57.705 157.875 ;
        RECT 56.745 157.865 57.705 157.870 ;
        RECT 56.745 157.855 57.695 157.865 ;
        RECT 56.745 157.850 57.685 157.855 ;
        RECT 56.745 157.840 57.675 157.850 ;
        RECT 56.745 157.830 57.670 157.840 ;
        RECT 56.745 157.825 57.665 157.830 ;
        RECT 56.745 157.810 57.655 157.825 ;
        RECT 56.745 157.795 57.650 157.810 ;
        RECT 56.745 157.770 57.640 157.795 ;
        RECT 56.745 157.700 57.635 157.770 ;
        RECT 53.525 156.595 56.115 157.365 ;
        RECT 56.745 157.145 57.295 157.530 ;
        RECT 57.465 156.975 57.635 157.700 ;
        RECT 56.745 156.805 57.635 156.975 ;
        RECT 57.805 157.300 58.135 157.725 ;
        RECT 58.305 157.500 58.535 157.895 ;
        RECT 57.805 156.815 58.025 157.300 ;
        RECT 58.705 157.245 58.875 158.275 ;
        RECT 58.195 156.595 58.445 157.135 ;
        RECT 58.615 156.765 58.875 157.245 ;
        RECT 60.630 157.140 60.970 157.970 ;
        RECT 62.450 157.460 62.800 158.710 ;
        RECT 66.150 157.140 66.490 157.970 ;
        RECT 67.970 157.460 68.320 158.710 ;
        RECT 71.005 158.425 71.465 158.975 ;
        RECT 71.655 158.425 71.985 159.145 ;
        RECT 59.045 156.595 64.390 157.140 ;
        RECT 64.565 156.595 69.910 157.140 ;
        RECT 71.005 157.055 71.255 158.425 ;
        RECT 72.185 158.255 72.485 158.805 ;
        RECT 72.655 158.475 72.935 159.145 ;
        RECT 73.305 158.590 73.910 159.145 ;
        RECT 74.085 158.635 74.565 158.975 ;
        RECT 74.735 158.600 74.990 159.145 ;
        RECT 73.305 158.490 73.920 158.590 ;
        RECT 73.735 158.465 73.920 158.490 ;
        RECT 71.545 158.085 72.485 158.255 ;
        RECT 71.545 157.835 71.715 158.085 ;
        RECT 72.855 157.835 73.120 158.195 ;
        RECT 71.425 157.505 71.715 157.835 ;
        RECT 71.885 157.585 72.225 157.835 ;
        RECT 72.445 157.585 73.120 157.835 ;
        RECT 73.305 157.870 73.565 158.320 ;
        RECT 73.735 158.220 74.065 158.465 ;
        RECT 74.235 158.145 74.990 158.395 ;
        RECT 75.160 158.275 75.435 158.975 ;
        RECT 74.220 158.110 74.990 158.145 ;
        RECT 74.205 158.100 74.990 158.110 ;
        RECT 74.200 158.085 75.095 158.100 ;
        RECT 74.180 158.070 75.095 158.085 ;
        RECT 74.160 158.060 75.095 158.070 ;
        RECT 74.135 158.050 75.095 158.060 ;
        RECT 74.065 158.020 75.095 158.050 ;
        RECT 74.045 157.990 75.095 158.020 ;
        RECT 74.025 157.960 75.095 157.990 ;
        RECT 73.995 157.935 75.095 157.960 ;
        RECT 73.960 157.900 75.095 157.935 ;
        RECT 73.930 157.895 75.095 157.900 ;
        RECT 73.930 157.890 74.320 157.895 ;
        RECT 73.930 157.880 74.295 157.890 ;
        RECT 73.930 157.875 74.280 157.880 ;
        RECT 73.930 157.870 74.265 157.875 ;
        RECT 73.305 157.865 74.265 157.870 ;
        RECT 73.305 157.855 74.255 157.865 ;
        RECT 73.305 157.850 74.245 157.855 ;
        RECT 73.305 157.840 74.235 157.850 ;
        RECT 73.305 157.830 74.230 157.840 ;
        RECT 73.305 157.825 74.225 157.830 ;
        RECT 73.305 157.810 74.215 157.825 ;
        RECT 73.305 157.795 74.210 157.810 ;
        RECT 73.305 157.770 74.200 157.795 ;
        RECT 73.305 157.700 74.195 157.770 ;
        RECT 71.545 157.415 71.715 157.505 ;
        RECT 71.545 157.225 72.935 157.415 ;
        RECT 71.005 156.765 71.565 157.055 ;
        RECT 71.735 156.595 71.985 157.055 ;
        RECT 72.605 156.865 72.935 157.225 ;
        RECT 73.305 157.145 73.855 157.530 ;
        RECT 74.025 156.975 74.195 157.700 ;
        RECT 73.305 156.805 74.195 156.975 ;
        RECT 74.365 157.300 74.695 157.725 ;
        RECT 74.865 157.500 75.095 157.895 ;
        RECT 74.365 156.815 74.585 157.300 ;
        RECT 75.265 157.245 75.435 158.275 ;
        RECT 75.605 157.980 75.895 159.145 ;
        RECT 76.065 158.055 77.275 159.145 ;
        RECT 76.065 157.345 76.585 157.885 ;
        RECT 76.755 157.515 77.275 158.055 ;
        RECT 77.445 158.295 77.825 158.975 ;
        RECT 78.415 158.295 78.585 159.145 ;
        RECT 78.755 158.465 79.085 158.975 ;
        RECT 79.255 158.635 79.425 159.145 ;
        RECT 79.595 158.465 79.995 158.975 ;
        RECT 78.755 158.295 79.995 158.465 ;
        RECT 74.755 156.595 75.005 157.135 ;
        RECT 75.175 156.765 75.435 157.245 ;
        RECT 75.605 156.595 75.895 157.320 ;
        RECT 76.065 156.595 77.275 157.345 ;
        RECT 77.445 157.335 77.615 158.295 ;
        RECT 77.785 157.955 79.090 158.125 ;
        RECT 80.175 158.045 80.495 158.975 ;
        RECT 80.665 158.055 84.175 159.145 ;
        RECT 77.785 157.505 78.030 157.955 ;
        RECT 78.200 157.585 78.750 157.785 ;
        RECT 78.920 157.755 79.090 157.955 ;
        RECT 79.865 157.875 80.495 158.045 ;
        RECT 78.920 157.585 79.295 157.755 ;
        RECT 79.465 157.335 79.695 157.835 ;
        RECT 77.445 157.165 79.695 157.335 ;
        RECT 77.495 156.595 77.825 156.985 ;
        RECT 77.995 156.845 78.165 157.165 ;
        RECT 79.865 156.995 80.035 157.875 ;
        RECT 78.335 156.595 78.665 156.985 ;
        RECT 79.080 156.825 80.035 156.995 ;
        RECT 80.205 156.595 80.495 157.430 ;
        RECT 80.665 157.365 82.315 157.885 ;
        RECT 82.485 157.535 84.175 158.055 ;
        RECT 84.345 158.005 84.625 159.145 ;
        RECT 84.795 157.995 85.125 158.975 ;
        RECT 85.295 158.005 85.555 159.145 ;
        RECT 85.815 158.135 85.985 158.975 ;
        RECT 86.155 158.805 87.325 158.975 ;
        RECT 86.155 158.305 86.485 158.805 ;
        RECT 86.995 158.765 87.325 158.805 ;
        RECT 87.515 158.725 87.870 159.145 ;
        RECT 86.655 158.545 86.885 158.635 ;
        RECT 88.040 158.545 88.290 158.975 ;
        RECT 86.655 158.305 88.290 158.545 ;
        RECT 88.460 158.385 88.790 159.145 ;
        RECT 88.960 158.305 89.215 158.975 ;
        RECT 84.860 157.955 85.035 157.995 ;
        RECT 85.815 157.965 88.875 158.135 ;
        RECT 84.355 157.565 84.690 157.835 ;
        RECT 84.860 157.395 85.030 157.955 ;
        RECT 85.200 157.585 85.535 157.835 ;
        RECT 85.730 157.585 86.080 157.795 ;
        RECT 86.250 157.585 86.695 157.785 ;
        RECT 86.865 157.585 87.340 157.785 ;
        RECT 80.665 156.595 84.175 157.365 ;
        RECT 84.345 156.595 84.655 157.395 ;
        RECT 84.860 156.765 85.555 157.395 ;
        RECT 85.815 157.245 86.880 157.415 ;
        RECT 85.815 156.765 85.985 157.245 ;
        RECT 86.155 156.595 86.485 157.075 ;
        RECT 86.710 157.015 86.880 157.245 ;
        RECT 87.060 157.185 87.340 157.585 ;
        RECT 87.610 157.585 87.940 157.785 ;
        RECT 88.110 157.585 88.475 157.785 ;
        RECT 87.610 157.185 87.895 157.585 ;
        RECT 88.705 157.415 88.875 157.965 ;
        RECT 88.075 157.245 88.875 157.415 ;
        RECT 88.075 157.015 88.245 157.245 ;
        RECT 89.045 157.175 89.215 158.305 ;
        RECT 89.590 158.175 89.980 158.350 ;
        RECT 90.465 158.345 90.795 159.145 ;
        RECT 90.965 158.355 91.500 158.975 ;
        RECT 89.590 158.005 91.015 158.175 ;
        RECT 89.465 157.275 89.820 157.835 ;
        RECT 89.030 157.095 89.215 157.175 ;
        RECT 89.990 157.105 90.160 158.005 ;
        RECT 90.330 157.275 90.595 157.835 ;
        RECT 90.845 157.505 91.015 158.005 ;
        RECT 91.185 157.335 91.500 158.355 ;
        RECT 91.705 158.055 93.375 159.145 ;
        RECT 86.710 156.765 88.245 157.015 ;
        RECT 88.415 156.595 88.745 157.075 ;
        RECT 88.960 156.765 89.215 157.095 ;
        RECT 89.570 156.595 89.810 157.105 ;
        RECT 89.990 156.775 90.270 157.105 ;
        RECT 90.500 156.595 90.715 157.105 ;
        RECT 90.885 156.765 91.500 157.335 ;
        RECT 91.705 157.365 92.455 157.885 ;
        RECT 92.625 157.535 93.375 158.055 ;
        RECT 93.545 158.005 93.885 158.975 ;
        RECT 94.055 158.005 94.225 159.145 ;
        RECT 94.495 158.345 94.745 159.145 ;
        RECT 95.390 158.175 95.720 158.975 ;
        RECT 96.020 158.345 96.350 159.145 ;
        RECT 96.520 158.175 96.850 158.975 ;
        RECT 94.415 158.005 96.850 158.175 ;
        RECT 97.235 158.085 97.565 158.935 ;
        RECT 93.545 157.395 93.720 158.005 ;
        RECT 94.415 157.755 94.585 158.005 ;
        RECT 93.890 157.585 94.585 157.755 ;
        RECT 94.760 157.585 95.180 157.785 ;
        RECT 95.350 157.585 95.680 157.785 ;
        RECT 95.850 157.585 96.180 157.785 ;
        RECT 91.705 156.595 93.375 157.365 ;
        RECT 93.545 156.765 93.885 157.395 ;
        RECT 94.055 156.595 94.305 157.395 ;
        RECT 94.495 157.245 95.720 157.415 ;
        RECT 94.495 156.765 94.825 157.245 ;
        RECT 94.995 156.595 95.220 157.055 ;
        RECT 95.390 156.765 95.720 157.245 ;
        RECT 96.350 157.375 96.520 158.005 ;
        RECT 97.235 157.955 97.455 158.085 ;
        RECT 97.735 158.005 97.985 159.145 ;
        RECT 98.175 158.505 98.425 158.925 ;
        RECT 98.655 158.675 98.985 159.145 ;
        RECT 99.215 158.505 99.465 158.925 ;
        RECT 98.175 158.335 99.465 158.505 ;
        RECT 99.645 158.505 99.975 158.935 ;
        RECT 99.645 158.335 100.100 158.505 ;
        RECT 96.705 157.585 97.055 157.835 ;
        RECT 96.350 156.765 96.850 157.375 ;
        RECT 97.235 157.320 97.425 157.955 ;
        RECT 98.165 157.835 98.380 158.165 ;
        RECT 97.595 157.505 97.905 157.835 ;
        RECT 98.075 157.505 98.380 157.835 ;
        RECT 98.555 157.505 98.840 158.165 ;
        RECT 99.035 157.505 99.300 158.165 ;
        RECT 99.515 157.505 99.760 158.165 ;
        RECT 97.735 157.335 97.905 157.505 ;
        RECT 99.930 157.335 100.100 158.335 ;
        RECT 101.365 157.980 101.655 159.145 ;
        RECT 101.845 158.635 102.145 159.145 ;
        RECT 102.315 158.635 102.695 158.805 ;
        RECT 103.275 158.635 103.905 159.145 ;
        RECT 102.315 158.465 102.485 158.635 ;
        RECT 104.075 158.465 104.405 158.975 ;
        RECT 104.575 158.635 104.875 159.145 ;
        RECT 101.825 158.265 102.485 158.465 ;
        RECT 102.655 158.295 104.875 158.465 ;
        RECT 97.235 156.810 97.565 157.320 ;
        RECT 97.735 157.165 100.100 157.335 ;
        RECT 101.825 157.335 101.995 158.265 ;
        RECT 102.655 158.095 102.825 158.295 ;
        RECT 102.165 157.925 102.825 158.095 ;
        RECT 102.995 157.955 104.535 158.125 ;
        RECT 102.165 157.505 102.335 157.925 ;
        RECT 102.995 157.755 103.165 157.955 ;
        RECT 102.565 157.585 103.165 157.755 ;
        RECT 103.335 157.585 104.030 157.785 ;
        RECT 104.290 157.505 104.535 157.955 ;
        RECT 102.655 157.335 103.565 157.415 ;
        RECT 97.735 156.595 98.065 156.995 ;
        RECT 99.115 156.825 99.445 157.165 ;
        RECT 99.615 156.595 99.945 156.995 ;
        RECT 101.365 156.595 101.655 157.320 ;
        RECT 101.825 156.855 102.145 157.335 ;
        RECT 102.315 157.245 103.565 157.335 ;
        RECT 102.315 157.165 102.825 157.245 ;
        RECT 102.315 156.765 102.545 157.165 ;
        RECT 102.715 156.595 103.065 156.985 ;
        RECT 103.235 156.765 103.565 157.245 ;
        RECT 103.735 156.595 103.905 157.415 ;
        RECT 104.705 157.335 104.875 158.295 ;
        RECT 105.045 158.055 108.555 159.145 ;
        RECT 104.410 156.790 104.875 157.335 ;
        RECT 105.045 157.365 106.695 157.885 ;
        RECT 106.865 157.535 108.555 158.055 ;
        RECT 109.645 158.175 109.955 158.975 ;
        RECT 110.125 158.345 110.435 159.145 ;
        RECT 110.605 158.515 110.865 158.975 ;
        RECT 111.035 158.685 111.290 159.145 ;
        RECT 111.465 158.515 111.725 158.975 ;
        RECT 110.605 158.345 111.725 158.515 ;
        RECT 109.645 158.005 110.675 158.175 ;
        RECT 105.045 156.595 108.555 157.365 ;
        RECT 109.645 157.095 109.815 158.005 ;
        RECT 109.985 157.265 110.335 157.835 ;
        RECT 110.505 157.755 110.675 158.005 ;
        RECT 111.465 158.095 111.725 158.345 ;
        RECT 111.895 158.275 112.180 159.145 ;
        RECT 112.405 158.710 117.750 159.145 ;
        RECT 117.925 158.710 123.270 159.145 ;
        RECT 111.465 157.925 112.220 158.095 ;
        RECT 110.505 157.585 111.645 157.755 ;
        RECT 111.815 157.415 112.220 157.925 ;
        RECT 110.570 157.245 112.220 157.415 ;
        RECT 109.645 156.765 109.945 157.095 ;
        RECT 110.115 156.595 110.390 157.075 ;
        RECT 110.570 156.855 110.865 157.245 ;
        RECT 111.035 156.595 111.290 157.075 ;
        RECT 111.465 156.855 111.725 157.245 ;
        RECT 113.990 157.140 114.330 157.970 ;
        RECT 115.810 157.460 116.160 158.710 ;
        RECT 119.510 157.140 119.850 157.970 ;
        RECT 121.330 157.460 121.680 158.710 ;
        RECT 123.445 158.055 126.955 159.145 ;
        RECT 123.445 157.365 125.095 157.885 ;
        RECT 125.265 157.535 126.955 158.055 ;
        RECT 127.125 157.980 127.415 159.145 ;
        RECT 127.585 158.710 132.930 159.145 ;
        RECT 133.105 158.710 138.450 159.145 ;
        RECT 138.625 158.710 143.970 159.145 ;
        RECT 111.895 156.595 112.175 157.075 ;
        RECT 112.405 156.595 117.750 157.140 ;
        RECT 117.925 156.595 123.270 157.140 ;
        RECT 123.445 156.595 126.955 157.365 ;
        RECT 127.125 156.595 127.415 157.320 ;
        RECT 129.170 157.140 129.510 157.970 ;
        RECT 130.990 157.460 131.340 158.710 ;
        RECT 134.690 157.140 135.030 157.970 ;
        RECT 136.510 157.460 136.860 158.710 ;
        RECT 140.210 157.140 140.550 157.970 ;
        RECT 142.030 157.460 142.380 158.710 ;
        RECT 144.145 158.055 147.655 159.145 ;
        RECT 147.825 158.055 149.035 159.145 ;
        RECT 144.145 157.365 145.795 157.885 ;
        RECT 145.965 157.535 147.655 158.055 ;
        RECT 127.585 156.595 132.930 157.140 ;
        RECT 133.105 156.595 138.450 157.140 ;
        RECT 138.625 156.595 143.970 157.140 ;
        RECT 144.145 156.595 147.655 157.365 ;
        RECT 147.825 157.345 148.345 157.885 ;
        RECT 148.515 157.515 149.035 158.055 ;
        RECT 149.205 158.055 150.415 159.145 ;
        RECT 149.205 157.515 149.725 158.055 ;
        RECT 149.895 157.345 150.415 157.885 ;
        RECT 147.825 156.595 149.035 157.345 ;
        RECT 149.205 156.595 150.415 157.345 ;
        RECT 11.120 156.425 150.500 156.595 ;
        RECT 11.205 155.675 12.415 156.425 ;
        RECT 12.585 155.880 17.930 156.425 ;
        RECT 11.205 155.135 11.725 155.675 ;
        RECT 11.895 154.965 12.415 155.505 ;
        RECT 14.170 155.050 14.510 155.880 ;
        RECT 18.105 155.750 18.365 156.255 ;
        RECT 18.545 156.045 18.875 156.425 ;
        RECT 19.055 155.875 19.225 156.255 ;
        RECT 19.485 155.880 24.830 156.425 ;
        RECT 11.205 153.875 12.415 154.965 ;
        RECT 15.990 154.310 16.340 155.560 ;
        RECT 18.105 154.950 18.275 155.750 ;
        RECT 18.560 155.705 19.225 155.875 ;
        RECT 18.560 155.450 18.730 155.705 ;
        RECT 18.445 155.120 18.730 155.450 ;
        RECT 18.965 155.155 19.295 155.525 ;
        RECT 18.560 154.975 18.730 155.120 ;
        RECT 21.070 155.050 21.410 155.880 ;
        RECT 25.005 155.655 28.515 156.425 ;
        RECT 29.145 155.925 29.405 156.255 ;
        RECT 29.575 156.065 29.905 156.425 ;
        RECT 30.160 156.045 31.460 156.255 ;
        RECT 29.145 155.915 29.375 155.925 ;
        RECT 12.585 153.875 17.930 154.310 ;
        RECT 18.105 154.045 18.375 154.950 ;
        RECT 18.560 154.805 19.225 154.975 ;
        RECT 18.545 153.875 18.875 154.635 ;
        RECT 19.055 154.045 19.225 154.805 ;
        RECT 22.890 154.310 23.240 155.560 ;
        RECT 25.005 155.135 26.655 155.655 ;
        RECT 26.825 154.965 28.515 155.485 ;
        RECT 19.485 153.875 24.830 154.310 ;
        RECT 25.005 153.875 28.515 154.965 ;
        RECT 29.145 154.725 29.315 155.915 ;
        RECT 30.160 155.895 30.330 156.045 ;
        RECT 29.575 155.770 30.330 155.895 ;
        RECT 29.485 155.725 30.330 155.770 ;
        RECT 29.485 155.605 29.755 155.725 ;
        RECT 29.485 155.030 29.655 155.605 ;
        RECT 29.885 155.165 30.295 155.470 ;
        RECT 30.585 155.435 30.795 155.835 ;
        RECT 30.465 155.225 30.795 155.435 ;
        RECT 31.040 155.435 31.260 155.835 ;
        RECT 31.735 155.660 32.190 156.425 ;
        RECT 32.365 155.675 33.575 156.425 ;
        RECT 33.745 155.685 34.210 156.230 ;
        RECT 31.040 155.225 31.515 155.435 ;
        RECT 31.705 155.235 32.195 155.435 ;
        RECT 32.365 155.135 32.885 155.675 ;
        RECT 29.485 154.995 29.685 155.030 ;
        RECT 31.015 154.995 32.190 155.055 ;
        RECT 29.485 154.885 32.190 154.995 ;
        RECT 33.055 154.965 33.575 155.505 ;
        RECT 29.545 154.825 31.345 154.885 ;
        RECT 31.015 154.795 31.345 154.825 ;
        RECT 29.145 154.045 29.405 154.725 ;
        RECT 29.575 153.875 29.825 154.655 ;
        RECT 30.075 154.625 30.910 154.635 ;
        RECT 31.500 154.625 31.685 154.715 ;
        RECT 30.075 154.425 31.685 154.625 ;
        RECT 30.075 154.045 30.325 154.425 ;
        RECT 31.455 154.385 31.685 154.425 ;
        RECT 31.935 154.265 32.190 154.885 ;
        RECT 30.495 153.875 30.850 154.255 ;
        RECT 31.855 154.045 32.190 154.265 ;
        RECT 32.365 153.875 33.575 154.965 ;
        RECT 33.745 154.725 33.915 155.685 ;
        RECT 34.715 155.605 34.885 156.425 ;
        RECT 35.055 155.775 35.385 156.255 ;
        RECT 35.555 156.035 35.905 156.425 ;
        RECT 36.075 155.855 36.305 156.255 ;
        RECT 35.795 155.775 36.305 155.855 ;
        RECT 35.055 155.685 36.305 155.775 ;
        RECT 36.475 155.685 36.795 156.165 ;
        RECT 36.965 155.700 37.255 156.425 ;
        RECT 35.055 155.605 35.965 155.685 ;
        RECT 34.085 155.065 34.330 155.515 ;
        RECT 34.590 155.235 35.285 155.435 ;
        RECT 35.455 155.265 36.055 155.435 ;
        RECT 35.455 155.065 35.625 155.265 ;
        RECT 36.285 155.095 36.455 155.515 ;
        RECT 34.085 154.895 35.625 155.065 ;
        RECT 35.795 154.925 36.455 155.095 ;
        RECT 35.795 154.725 35.965 154.925 ;
        RECT 36.625 154.755 36.795 155.685 ;
        RECT 37.425 155.675 38.635 156.425 ;
        RECT 38.815 155.915 39.265 156.425 ;
        RECT 39.540 156.005 40.845 156.255 ;
        RECT 41.025 156.025 41.355 156.425 ;
        RECT 40.665 155.855 40.845 156.005 ;
        RECT 37.425 155.135 37.945 155.675 ;
        RECT 33.745 154.555 35.965 154.725 ;
        RECT 36.135 154.555 36.795 154.755 ;
        RECT 33.745 153.875 34.045 154.385 ;
        RECT 34.215 154.045 34.545 154.555 ;
        RECT 36.135 154.385 36.305 154.555 ;
        RECT 34.715 153.875 35.345 154.385 ;
        RECT 35.925 154.215 36.305 154.385 ;
        RECT 36.475 153.875 36.775 154.385 ;
        RECT 36.965 153.875 37.255 155.040 ;
        RECT 38.115 154.965 38.635 155.505 ;
        RECT 38.845 155.235 39.295 155.745 ;
        RECT 39.710 155.435 39.960 155.835 ;
        RECT 39.485 155.235 39.960 155.435 ;
        RECT 40.210 155.435 40.420 155.835 ;
        RECT 40.665 155.685 41.395 155.855 ;
        RECT 41.585 155.695 41.875 156.425 ;
        RECT 40.210 155.235 40.560 155.435 ;
        RECT 40.730 155.185 41.055 155.515 ;
        RECT 37.425 153.875 38.635 154.965 ;
        RECT 38.815 155.015 40.560 155.065 ;
        RECT 41.225 155.015 41.395 155.685 ;
        RECT 41.575 155.185 41.875 155.515 ;
        RECT 42.055 155.495 42.285 156.135 ;
        RECT 42.465 155.875 42.775 156.245 ;
        RECT 42.955 156.055 43.625 156.425 ;
        RECT 42.465 155.675 43.695 155.875 ;
        RECT 42.055 155.185 42.580 155.495 ;
        RECT 42.760 155.185 43.225 155.495 ;
        RECT 38.815 154.885 41.395 155.015 ;
        RECT 43.405 155.005 43.695 155.675 ;
        RECT 38.815 154.215 39.145 154.885 ;
        RECT 40.335 154.845 41.395 154.885 ;
        RECT 41.585 154.765 42.745 155.005 ;
        RECT 39.315 154.675 40.195 154.715 ;
        RECT 39.315 154.475 40.845 154.675 ;
        RECT 39.315 154.425 39.930 154.475 ;
        RECT 39.315 154.385 39.545 154.425 ;
        RECT 40.675 154.345 40.845 154.475 ;
        RECT 39.655 154.215 39.985 154.255 ;
        RECT 38.815 154.045 39.985 154.215 ;
        RECT 40.155 153.875 40.530 154.255 ;
        RECT 41.080 153.875 41.345 154.655 ;
        RECT 41.585 154.055 41.845 154.765 ;
        RECT 42.015 153.875 42.345 154.585 ;
        RECT 42.515 154.055 42.745 154.765 ;
        RECT 42.925 154.785 43.695 155.005 ;
        RECT 42.925 154.055 43.195 154.785 ;
        RECT 43.375 153.875 43.715 154.605 ;
        RECT 43.885 154.055 44.145 156.245 ;
        RECT 44.485 155.865 44.815 156.255 ;
        RECT 44.985 156.035 46.170 156.205 ;
        RECT 46.430 155.955 46.600 156.425 ;
        RECT 44.485 155.685 44.995 155.865 ;
        RECT 44.325 155.225 44.655 155.515 ;
        RECT 44.825 155.055 44.995 155.685 ;
        RECT 45.400 155.775 45.785 155.865 ;
        RECT 46.770 155.775 47.100 156.240 ;
        RECT 45.400 155.605 47.100 155.775 ;
        RECT 47.270 155.605 47.440 156.425 ;
        RECT 47.610 155.605 48.295 156.245 ;
        RECT 48.705 155.955 48.875 156.425 ;
        RECT 49.545 155.955 49.715 156.425 ;
        RECT 49.980 156.035 51.210 156.255 ;
        RECT 49.045 155.785 49.375 155.865 ;
        RECT 50.405 155.785 50.735 155.865 ;
        RECT 45.165 155.225 45.495 155.435 ;
        RECT 45.675 155.185 46.055 155.435 ;
        RECT 44.480 154.885 45.565 155.055 ;
        RECT 44.480 154.045 44.780 154.885 ;
        RECT 44.975 153.875 45.225 154.715 ;
        RECT 45.395 154.635 45.565 154.885 ;
        RECT 45.735 154.805 46.055 155.185 ;
        RECT 46.245 155.225 46.730 155.435 ;
        RECT 46.920 155.225 47.370 155.435 ;
        RECT 47.540 155.225 47.875 155.435 ;
        RECT 46.245 155.065 46.620 155.225 ;
        RECT 46.225 154.895 46.620 155.065 ;
        RECT 47.540 155.055 47.710 155.225 ;
        RECT 46.245 154.805 46.620 154.895 ;
        RECT 46.790 154.885 47.710 155.055 ;
        RECT 46.790 154.635 46.960 154.885 ;
        RECT 45.395 154.465 46.960 154.635 ;
        RECT 45.815 154.045 46.620 154.465 ;
        RECT 47.130 153.875 47.460 154.715 ;
        RECT 48.045 154.635 48.295 155.605 ;
        RECT 48.465 155.605 50.735 155.785 ;
        RECT 50.960 155.785 51.210 156.035 ;
        RECT 51.380 155.955 51.550 156.425 ;
        RECT 51.720 155.785 52.050 156.255 ;
        RECT 52.320 155.955 52.490 156.425 ;
        RECT 50.960 155.605 52.050 155.785 ;
        RECT 52.660 155.785 52.990 156.255 ;
        RECT 53.160 155.955 53.330 156.425 ;
        RECT 53.500 155.785 53.830 156.255 ;
        RECT 54.000 155.955 54.170 156.425 ;
        RECT 52.660 155.605 54.240 155.785 ;
        RECT 48.465 155.095 48.875 155.605 ;
        RECT 49.085 155.265 49.745 155.435 ;
        RECT 48.465 154.885 49.335 155.095 ;
        RECT 49.575 155.065 49.745 155.265 ;
        RECT 50.270 155.235 50.940 155.435 ;
        RECT 51.130 155.235 52.650 155.435 ;
        RECT 52.820 155.235 53.315 155.435 ;
        RECT 53.485 155.235 53.815 155.435 ;
        RECT 52.480 155.065 52.650 155.235 ;
        RECT 53.485 155.065 53.655 155.235 ;
        RECT 49.575 154.895 52.310 155.065 ;
        RECT 52.480 154.895 53.655 155.065 ;
        RECT 47.630 154.045 48.295 154.635 ;
        RECT 48.665 154.215 48.915 154.715 ;
        RECT 49.085 154.385 49.335 154.885 ;
        RECT 52.140 154.725 52.310 154.895 ;
        RECT 54.070 154.725 54.240 155.605 ;
        RECT 54.445 155.655 56.115 156.425 ;
        RECT 54.445 155.135 55.195 155.655 ;
        RECT 56.285 155.625 56.595 156.425 ;
        RECT 56.800 155.625 57.495 156.255 ;
        RECT 57.665 155.675 58.875 156.425 ;
        RECT 59.135 155.875 59.305 156.255 ;
        RECT 59.485 156.045 59.815 156.425 ;
        RECT 59.135 155.705 59.800 155.875 ;
        RECT 59.995 155.750 60.255 156.255 ;
        RECT 55.365 154.965 56.115 155.485 ;
        RECT 56.295 155.185 56.630 155.455 ;
        RECT 56.800 155.025 56.970 155.625 ;
        RECT 57.140 155.185 57.475 155.435 ;
        RECT 57.665 155.135 58.185 155.675 ;
        RECT 49.505 154.555 51.970 154.725 ;
        RECT 52.140 154.555 54.240 154.725 ;
        RECT 49.505 154.215 50.275 154.555 ;
        RECT 48.665 154.045 50.275 154.215 ;
        RECT 50.445 153.875 50.750 154.375 ;
        RECT 50.920 154.045 51.170 154.555 ;
        RECT 51.760 154.385 51.970 154.555 ;
        RECT 52.700 154.385 52.950 154.555 ;
        RECT 51.340 153.875 51.590 154.375 ;
        RECT 51.760 154.045 52.075 154.385 ;
        RECT 53.125 154.375 53.295 154.385 ;
        RECT 54.045 154.375 54.215 154.385 ;
        RECT 52.280 154.215 52.530 154.375 ;
        RECT 53.120 154.215 53.370 154.375 ;
        RECT 52.280 154.045 53.370 154.215 ;
        RECT 53.540 153.875 53.790 154.375 ;
        RECT 53.960 154.045 54.240 154.375 ;
        RECT 54.445 153.875 56.115 154.965 ;
        RECT 56.285 153.875 56.565 155.015 ;
        RECT 56.735 154.045 57.065 155.025 ;
        RECT 57.235 153.875 57.495 155.015 ;
        RECT 58.355 154.965 58.875 155.505 ;
        RECT 59.065 155.155 59.395 155.525 ;
        RECT 59.630 155.450 59.800 155.705 ;
        RECT 59.630 155.120 59.915 155.450 ;
        RECT 59.630 154.975 59.800 155.120 ;
        RECT 57.665 153.875 58.875 154.965 ;
        RECT 59.135 154.805 59.800 154.975 ;
        RECT 60.085 154.950 60.255 155.750 ;
        RECT 60.425 155.655 62.095 156.425 ;
        RECT 62.725 155.700 63.015 156.425 ;
        RECT 64.195 155.875 64.365 156.165 ;
        RECT 64.535 156.045 64.865 156.425 ;
        RECT 64.195 155.705 64.860 155.875 ;
        RECT 60.425 155.135 61.175 155.655 ;
        RECT 61.345 154.965 62.095 155.485 ;
        RECT 59.135 154.045 59.305 154.805 ;
        RECT 59.485 153.875 59.815 154.635 ;
        RECT 59.985 154.045 60.255 154.950 ;
        RECT 60.425 153.875 62.095 154.965 ;
        RECT 62.725 153.875 63.015 155.040 ;
        RECT 64.110 154.885 64.460 155.535 ;
        RECT 64.630 154.715 64.860 155.705 ;
        RECT 64.195 154.545 64.860 154.715 ;
        RECT 64.195 154.045 64.365 154.545 ;
        RECT 64.535 153.875 64.865 154.375 ;
        RECT 65.035 154.045 65.220 156.165 ;
        RECT 65.475 155.965 65.725 156.425 ;
        RECT 65.895 155.975 66.230 156.145 ;
        RECT 66.425 155.975 67.100 156.145 ;
        RECT 65.895 155.835 66.065 155.975 ;
        RECT 65.390 154.845 65.670 155.795 ;
        RECT 65.840 155.705 66.065 155.835 ;
        RECT 65.840 154.600 66.010 155.705 ;
        RECT 66.235 155.555 66.760 155.775 ;
        RECT 66.180 154.790 66.420 155.385 ;
        RECT 66.590 154.855 66.760 155.555 ;
        RECT 66.930 155.195 67.100 155.975 ;
        RECT 67.420 155.925 67.790 156.425 ;
        RECT 67.970 155.975 68.375 156.145 ;
        RECT 68.545 155.975 69.330 156.145 ;
        RECT 67.970 155.745 68.140 155.975 ;
        RECT 67.310 155.445 68.140 155.745 ;
        RECT 68.525 155.475 68.990 155.805 ;
        RECT 67.310 155.415 67.510 155.445 ;
        RECT 67.630 155.195 67.800 155.265 ;
        RECT 66.930 155.025 67.800 155.195 ;
        RECT 67.290 154.935 67.800 155.025 ;
        RECT 65.840 154.470 66.145 154.600 ;
        RECT 66.590 154.490 67.120 154.855 ;
        RECT 65.460 153.875 65.725 154.335 ;
        RECT 65.895 154.045 66.145 154.470 ;
        RECT 67.290 154.320 67.460 154.935 ;
        RECT 66.355 154.150 67.460 154.320 ;
        RECT 67.630 153.875 67.800 154.675 ;
        RECT 67.970 154.375 68.140 155.445 ;
        RECT 68.310 154.545 68.500 155.265 ;
        RECT 68.670 154.515 68.990 155.475 ;
        RECT 69.160 155.515 69.330 155.975 ;
        RECT 69.605 155.895 69.815 156.425 ;
        RECT 70.075 155.685 70.405 156.210 ;
        RECT 70.575 155.815 70.745 156.425 ;
        RECT 70.915 155.770 71.245 156.205 ;
        RECT 71.415 155.910 71.585 156.425 ;
        RECT 72.390 155.895 72.680 156.245 ;
        RECT 72.875 156.065 73.205 156.425 ;
        RECT 73.375 155.895 73.605 156.200 ;
        RECT 70.915 155.685 71.295 155.770 ;
        RECT 72.390 155.725 73.605 155.895 ;
        RECT 70.205 155.515 70.405 155.685 ;
        RECT 71.070 155.645 71.295 155.685 ;
        RECT 69.160 155.185 70.035 155.515 ;
        RECT 70.205 155.185 70.955 155.515 ;
        RECT 67.970 154.045 68.220 154.375 ;
        RECT 69.160 154.345 69.330 155.185 ;
        RECT 70.205 154.980 70.395 155.185 ;
        RECT 71.125 155.065 71.295 155.645 ;
        RECT 73.795 155.555 73.965 156.120 ;
        RECT 74.225 155.880 79.570 156.425 ;
        RECT 72.450 155.405 72.710 155.515 ;
        RECT 72.445 155.235 72.710 155.405 ;
        RECT 72.450 155.185 72.710 155.235 ;
        RECT 72.890 155.185 73.275 155.515 ;
        RECT 73.445 155.385 73.965 155.555 ;
        RECT 71.080 155.015 71.295 155.065 ;
        RECT 69.500 154.605 70.395 154.980 ;
        RECT 70.905 154.935 71.295 155.015 ;
        RECT 68.445 154.175 69.330 154.345 ;
        RECT 69.510 153.875 69.825 154.375 ;
        RECT 70.055 154.045 70.395 154.605 ;
        RECT 70.565 153.875 70.735 154.885 ;
        RECT 70.905 154.090 71.235 154.935 ;
        RECT 71.405 153.875 71.575 154.790 ;
        RECT 72.390 153.875 72.710 155.015 ;
        RECT 72.890 154.135 73.085 155.185 ;
        RECT 73.445 155.005 73.615 155.385 ;
        RECT 73.265 154.725 73.615 155.005 ;
        RECT 73.805 154.855 74.050 155.215 ;
        RECT 75.810 155.050 76.150 155.880 ;
        RECT 79.745 155.655 83.255 156.425 ;
        RECT 83.425 156.045 84.315 156.215 ;
        RECT 73.265 154.045 73.595 154.725 ;
        RECT 73.795 153.875 74.050 154.675 ;
        RECT 77.630 154.310 77.980 155.560 ;
        RECT 79.745 155.135 81.395 155.655 ;
        RECT 83.425 155.490 83.975 155.875 ;
        RECT 81.565 154.965 83.255 155.485 ;
        RECT 84.145 155.320 84.315 156.045 ;
        RECT 74.225 153.875 79.570 154.310 ;
        RECT 79.745 153.875 83.255 154.965 ;
        RECT 83.425 155.250 84.315 155.320 ;
        RECT 84.485 155.745 84.705 156.205 ;
        RECT 84.875 155.885 85.125 156.425 ;
        RECT 85.295 155.775 85.555 156.255 ;
        RECT 84.485 155.720 84.735 155.745 ;
        RECT 84.485 155.295 84.815 155.720 ;
        RECT 83.425 155.225 84.320 155.250 ;
        RECT 83.425 155.210 84.330 155.225 ;
        RECT 83.425 155.195 84.335 155.210 ;
        RECT 83.425 155.190 84.345 155.195 ;
        RECT 83.425 155.180 84.350 155.190 ;
        RECT 83.425 155.170 84.355 155.180 ;
        RECT 83.425 155.165 84.365 155.170 ;
        RECT 83.425 155.155 84.375 155.165 ;
        RECT 83.425 155.150 84.385 155.155 ;
        RECT 83.425 154.700 83.685 155.150 ;
        RECT 84.050 155.145 84.385 155.150 ;
        RECT 84.050 155.140 84.400 155.145 ;
        RECT 84.050 155.130 84.415 155.140 ;
        RECT 84.050 155.125 84.440 155.130 ;
        RECT 84.985 155.125 85.215 155.520 ;
        RECT 84.050 155.120 85.215 155.125 ;
        RECT 84.080 155.085 85.215 155.120 ;
        RECT 84.115 155.060 85.215 155.085 ;
        RECT 84.145 155.030 85.215 155.060 ;
        RECT 84.165 155.000 85.215 155.030 ;
        RECT 84.185 154.970 85.215 155.000 ;
        RECT 84.255 154.960 85.215 154.970 ;
        RECT 84.280 154.950 85.215 154.960 ;
        RECT 84.300 154.935 85.215 154.950 ;
        RECT 84.320 154.920 85.215 154.935 ;
        RECT 84.325 154.910 85.110 154.920 ;
        RECT 84.340 154.875 85.110 154.910 ;
        RECT 83.855 154.555 84.185 154.800 ;
        RECT 84.355 154.625 85.110 154.875 ;
        RECT 85.385 154.745 85.555 155.775 ;
        RECT 85.725 155.675 86.935 156.425 ;
        RECT 85.725 155.135 86.245 155.675 ;
        RECT 87.115 155.615 87.385 156.425 ;
        RECT 87.555 155.615 87.885 156.255 ;
        RECT 88.055 155.615 88.295 156.425 ;
        RECT 88.485 155.700 88.775 156.425 ;
        RECT 88.945 155.655 92.455 156.425 ;
        RECT 92.710 155.855 92.885 156.255 ;
        RECT 93.055 156.045 93.385 156.425 ;
        RECT 93.630 155.925 93.860 156.255 ;
        RECT 92.710 155.685 93.340 155.855 ;
        RECT 86.415 154.965 86.935 155.505 ;
        RECT 87.105 155.185 87.455 155.435 ;
        RECT 87.625 155.015 87.795 155.615 ;
        RECT 87.965 155.185 88.315 155.435 ;
        RECT 88.945 155.135 90.595 155.655 ;
        RECT 93.170 155.515 93.340 155.685 ;
        RECT 83.855 154.530 84.040 154.555 ;
        RECT 83.425 154.430 84.040 154.530 ;
        RECT 83.425 153.875 84.030 154.430 ;
        RECT 84.205 154.045 84.685 154.385 ;
        RECT 84.855 153.875 85.110 154.420 ;
        RECT 85.280 154.045 85.555 154.745 ;
        RECT 85.725 153.875 86.935 154.965 ;
        RECT 87.115 153.875 87.445 155.015 ;
        RECT 87.625 154.845 88.305 155.015 ;
        RECT 87.975 154.060 88.305 154.845 ;
        RECT 88.485 153.875 88.775 155.040 ;
        RECT 90.765 154.965 92.455 155.485 ;
        RECT 88.945 153.875 92.455 154.965 ;
        RECT 92.625 154.835 92.990 155.515 ;
        RECT 93.170 155.185 93.520 155.515 ;
        RECT 93.170 154.665 93.340 155.185 ;
        RECT 92.710 154.495 93.340 154.665 ;
        RECT 93.690 154.635 93.860 155.925 ;
        RECT 94.060 154.815 94.340 156.090 ;
        RECT 94.565 155.065 94.835 156.090 ;
        RECT 95.295 156.045 95.625 156.425 ;
        RECT 95.795 156.170 96.130 156.215 ;
        RECT 94.525 154.895 94.835 155.065 ;
        RECT 94.565 154.815 94.835 154.895 ;
        RECT 95.025 154.815 95.365 155.845 ;
        RECT 95.795 155.705 96.135 156.170 ;
        RECT 95.535 155.185 95.795 155.515 ;
        RECT 95.535 154.635 95.705 155.185 ;
        RECT 95.965 155.015 96.135 155.705 ;
        RECT 92.710 154.045 92.885 154.495 ;
        RECT 93.690 154.465 95.705 154.635 ;
        RECT 93.055 153.875 93.385 154.315 ;
        RECT 93.690 154.045 93.860 154.465 ;
        RECT 94.095 153.875 94.765 154.285 ;
        RECT 94.980 154.045 95.150 154.465 ;
        RECT 95.350 153.875 95.680 154.285 ;
        RECT 95.875 154.045 96.135 155.015 ;
        RECT 96.305 155.775 96.565 156.255 ;
        RECT 96.735 155.965 97.065 156.425 ;
        RECT 97.255 155.785 97.455 156.205 ;
        RECT 96.305 154.745 96.475 155.775 ;
        RECT 96.645 155.085 96.875 155.515 ;
        RECT 97.045 155.265 97.455 155.785 ;
        RECT 97.625 155.940 98.415 156.205 ;
        RECT 97.625 155.085 97.880 155.940 ;
        RECT 98.595 155.605 98.925 156.025 ;
        RECT 99.095 155.605 99.355 156.425 ;
        RECT 100.445 155.775 100.705 156.255 ;
        RECT 100.875 155.885 101.125 156.425 ;
        RECT 98.595 155.515 98.845 155.605 ;
        RECT 98.050 155.265 98.845 155.515 ;
        RECT 96.645 154.915 98.435 155.085 ;
        RECT 96.305 154.045 96.580 154.745 ;
        RECT 96.750 154.620 97.465 154.915 ;
        RECT 97.685 154.555 98.015 154.745 ;
        RECT 96.790 153.875 97.005 154.420 ;
        RECT 97.175 154.045 97.650 154.385 ;
        RECT 97.820 154.380 98.015 154.555 ;
        RECT 98.185 154.550 98.435 154.915 ;
        RECT 97.820 153.875 98.435 154.380 ;
        RECT 98.675 154.045 98.845 155.265 ;
        RECT 99.015 154.555 99.355 155.435 ;
        RECT 100.445 154.745 100.615 155.775 ;
        RECT 101.295 155.720 101.515 156.205 ;
        RECT 100.785 155.125 101.015 155.520 ;
        RECT 101.185 155.295 101.515 155.720 ;
        RECT 101.685 156.045 102.575 156.215 ;
        RECT 101.685 155.320 101.855 156.045 ;
        RECT 102.745 155.880 108.090 156.425 ;
        RECT 102.025 155.490 102.575 155.875 ;
        RECT 101.685 155.250 102.575 155.320 ;
        RECT 101.680 155.225 102.575 155.250 ;
        RECT 101.670 155.210 102.575 155.225 ;
        RECT 101.665 155.195 102.575 155.210 ;
        RECT 101.655 155.190 102.575 155.195 ;
        RECT 101.650 155.180 102.575 155.190 ;
        RECT 101.645 155.170 102.575 155.180 ;
        RECT 101.635 155.165 102.575 155.170 ;
        RECT 101.625 155.155 102.575 155.165 ;
        RECT 101.615 155.150 102.575 155.155 ;
        RECT 101.615 155.145 101.950 155.150 ;
        RECT 101.600 155.140 101.950 155.145 ;
        RECT 101.585 155.130 101.950 155.140 ;
        RECT 101.560 155.125 101.950 155.130 ;
        RECT 100.785 155.120 101.950 155.125 ;
        RECT 100.785 155.085 101.920 155.120 ;
        RECT 100.785 155.060 101.885 155.085 ;
        RECT 100.785 155.030 101.855 155.060 ;
        RECT 100.785 155.000 101.835 155.030 ;
        RECT 100.785 154.970 101.815 155.000 ;
        RECT 100.785 154.960 101.745 154.970 ;
        RECT 100.785 154.950 101.720 154.960 ;
        RECT 100.785 154.935 101.700 154.950 ;
        RECT 100.785 154.920 101.680 154.935 ;
        RECT 100.890 154.910 101.675 154.920 ;
        RECT 100.890 154.875 101.660 154.910 ;
        RECT 99.095 153.875 99.355 154.385 ;
        RECT 100.445 154.045 100.720 154.745 ;
        RECT 100.890 154.625 101.645 154.875 ;
        RECT 101.815 154.555 102.145 154.800 ;
        RECT 102.315 154.700 102.575 155.150 ;
        RECT 104.330 155.050 104.670 155.880 ;
        RECT 108.265 155.625 108.960 156.255 ;
        RECT 109.165 155.625 109.475 156.425 ;
        RECT 109.645 155.655 113.155 156.425 ;
        RECT 114.245 155.700 114.535 156.425 ;
        RECT 114.705 155.880 120.050 156.425 ;
        RECT 120.225 155.880 125.570 156.425 ;
        RECT 125.745 155.880 131.090 156.425 ;
        RECT 131.265 155.880 136.610 156.425 ;
        RECT 101.960 154.530 102.145 154.555 ;
        RECT 101.960 154.430 102.575 154.530 ;
        RECT 100.890 153.875 101.145 154.420 ;
        RECT 101.315 154.045 101.795 154.385 ;
        RECT 101.970 153.875 102.575 154.430 ;
        RECT 106.150 154.310 106.500 155.560 ;
        RECT 108.285 155.185 108.620 155.435 ;
        RECT 108.790 155.025 108.960 155.625 ;
        RECT 109.130 155.185 109.465 155.455 ;
        RECT 109.645 155.135 111.295 155.655 ;
        RECT 102.745 153.875 108.090 154.310 ;
        RECT 108.265 153.875 108.525 155.015 ;
        RECT 108.695 154.045 109.025 155.025 ;
        RECT 109.195 153.875 109.475 155.015 ;
        RECT 111.465 154.965 113.155 155.485 ;
        RECT 116.290 155.050 116.630 155.880 ;
        RECT 109.645 153.875 113.155 154.965 ;
        RECT 114.245 153.875 114.535 155.040 ;
        RECT 118.110 154.310 118.460 155.560 ;
        RECT 121.810 155.050 122.150 155.880 ;
        RECT 123.630 154.310 123.980 155.560 ;
        RECT 127.330 155.050 127.670 155.880 ;
        RECT 129.150 154.310 129.500 155.560 ;
        RECT 132.850 155.050 133.190 155.880 ;
        RECT 136.785 155.655 139.375 156.425 ;
        RECT 140.005 155.700 140.295 156.425 ;
        RECT 140.465 155.880 145.810 156.425 ;
        RECT 134.670 154.310 135.020 155.560 ;
        RECT 136.785 155.135 137.995 155.655 ;
        RECT 138.165 154.965 139.375 155.485 ;
        RECT 142.050 155.050 142.390 155.880 ;
        RECT 145.985 155.655 148.575 156.425 ;
        RECT 149.205 155.675 150.415 156.425 ;
        RECT 114.705 153.875 120.050 154.310 ;
        RECT 120.225 153.875 125.570 154.310 ;
        RECT 125.745 153.875 131.090 154.310 ;
        RECT 131.265 153.875 136.610 154.310 ;
        RECT 136.785 153.875 139.375 154.965 ;
        RECT 140.005 153.875 140.295 155.040 ;
        RECT 143.870 154.310 144.220 155.560 ;
        RECT 145.985 155.135 147.195 155.655 ;
        RECT 147.365 154.965 148.575 155.485 ;
        RECT 140.465 153.875 145.810 154.310 ;
        RECT 145.985 153.875 148.575 154.965 ;
        RECT 149.205 154.965 149.725 155.505 ;
        RECT 149.895 155.135 150.415 155.675 ;
        RECT 149.205 153.875 150.415 154.965 ;
        RECT 11.120 153.705 150.500 153.875 ;
        RECT 11.205 152.615 12.415 153.705 ;
        RECT 12.585 152.615 15.175 153.705 ;
        RECT 15.895 153.035 16.065 153.535 ;
        RECT 16.235 153.205 16.565 153.705 ;
        RECT 15.895 152.865 16.560 153.035 ;
        RECT 11.205 151.905 11.725 152.445 ;
        RECT 11.895 152.075 12.415 152.615 ;
        RECT 12.585 151.925 13.795 152.445 ;
        RECT 13.965 152.095 15.175 152.615 ;
        RECT 15.810 152.045 16.160 152.695 ;
        RECT 11.205 151.155 12.415 151.905 ;
        RECT 12.585 151.155 15.175 151.925 ;
        RECT 16.330 151.875 16.560 152.865 ;
        RECT 15.895 151.705 16.560 151.875 ;
        RECT 15.895 151.415 16.065 151.705 ;
        RECT 16.235 151.155 16.565 151.535 ;
        RECT 16.735 151.415 16.920 153.535 ;
        RECT 17.160 153.245 17.425 153.705 ;
        RECT 17.595 153.110 17.845 153.535 ;
        RECT 18.055 153.260 19.160 153.430 ;
        RECT 17.540 152.980 17.845 153.110 ;
        RECT 17.090 151.785 17.370 152.735 ;
        RECT 17.540 151.875 17.710 152.980 ;
        RECT 17.880 152.195 18.120 152.790 ;
        RECT 18.290 152.725 18.820 153.090 ;
        RECT 18.290 152.025 18.460 152.725 ;
        RECT 18.990 152.645 19.160 153.260 ;
        RECT 19.330 152.905 19.500 153.705 ;
        RECT 19.670 153.205 19.920 153.535 ;
        RECT 20.145 153.235 21.030 153.405 ;
        RECT 18.990 152.555 19.500 152.645 ;
        RECT 17.540 151.745 17.765 151.875 ;
        RECT 17.935 151.805 18.460 152.025 ;
        RECT 18.630 152.385 19.500 152.555 ;
        RECT 17.175 151.155 17.425 151.615 ;
        RECT 17.595 151.605 17.765 151.745 ;
        RECT 18.630 151.605 18.800 152.385 ;
        RECT 19.330 152.315 19.500 152.385 ;
        RECT 19.010 152.135 19.210 152.165 ;
        RECT 19.670 152.135 19.840 153.205 ;
        RECT 20.010 152.315 20.200 153.035 ;
        RECT 19.010 151.835 19.840 152.135 ;
        RECT 20.370 152.105 20.690 153.065 ;
        RECT 17.595 151.435 17.930 151.605 ;
        RECT 18.125 151.435 18.800 151.605 ;
        RECT 19.120 151.155 19.490 151.655 ;
        RECT 19.670 151.605 19.840 151.835 ;
        RECT 20.225 151.775 20.690 152.105 ;
        RECT 20.860 152.395 21.030 153.235 ;
        RECT 21.210 153.205 21.525 153.705 ;
        RECT 21.755 152.975 22.095 153.535 ;
        RECT 21.200 152.600 22.095 152.975 ;
        RECT 22.265 152.695 22.435 153.705 ;
        RECT 21.905 152.395 22.095 152.600 ;
        RECT 22.605 152.645 22.935 153.490 ;
        RECT 22.605 152.565 22.995 152.645 ;
        RECT 22.780 152.515 22.995 152.565 ;
        RECT 24.085 152.540 24.375 153.705 ;
        RECT 24.545 153.195 24.845 153.705 ;
        RECT 25.015 153.025 25.345 153.535 ;
        RECT 25.515 153.195 26.145 153.705 ;
        RECT 26.725 153.195 27.105 153.365 ;
        RECT 27.275 153.195 27.575 153.705 ;
        RECT 26.935 153.025 27.105 153.195 ;
        RECT 24.545 152.855 26.765 153.025 ;
        RECT 20.860 152.065 21.735 152.395 ;
        RECT 21.905 152.065 22.655 152.395 ;
        RECT 20.860 151.605 21.030 152.065 ;
        RECT 21.905 151.895 22.105 152.065 ;
        RECT 22.825 151.935 22.995 152.515 ;
        RECT 22.770 151.895 22.995 151.935 ;
        RECT 19.670 151.435 20.075 151.605 ;
        RECT 20.245 151.435 21.030 151.605 ;
        RECT 21.305 151.155 21.515 151.685 ;
        RECT 21.775 151.370 22.105 151.895 ;
        RECT 22.615 151.810 22.995 151.895 ;
        RECT 24.545 151.895 24.715 152.855 ;
        RECT 24.885 152.515 26.425 152.685 ;
        RECT 24.885 152.065 25.130 152.515 ;
        RECT 25.390 152.145 26.085 152.345 ;
        RECT 26.255 152.315 26.425 152.515 ;
        RECT 26.595 152.655 26.765 152.855 ;
        RECT 26.935 152.825 27.595 153.025 ;
        RECT 26.595 152.485 27.255 152.655 ;
        RECT 26.255 152.145 26.855 152.315 ;
        RECT 27.085 152.065 27.255 152.485 ;
        RECT 22.275 151.155 22.445 151.765 ;
        RECT 22.615 151.375 22.945 151.810 ;
        RECT 24.085 151.155 24.375 151.880 ;
        RECT 24.545 151.350 25.010 151.895 ;
        RECT 25.515 151.155 25.685 151.975 ;
        RECT 25.855 151.895 26.765 151.975 ;
        RECT 27.425 151.895 27.595 152.825 ;
        RECT 27.765 152.615 29.435 153.705 ;
        RECT 25.855 151.805 27.105 151.895 ;
        RECT 25.855 151.325 26.185 151.805 ;
        RECT 26.595 151.725 27.105 151.805 ;
        RECT 26.355 151.155 26.705 151.545 ;
        RECT 26.875 151.325 27.105 151.725 ;
        RECT 27.275 151.415 27.595 151.895 ;
        RECT 27.765 151.925 28.515 152.445 ;
        RECT 28.685 152.095 29.435 152.615 ;
        RECT 29.605 152.855 29.865 153.535 ;
        RECT 30.035 152.925 30.285 153.705 ;
        RECT 30.535 153.155 30.785 153.535 ;
        RECT 30.955 153.325 31.310 153.705 ;
        RECT 32.315 153.315 32.650 153.535 ;
        RECT 31.915 153.155 32.145 153.195 ;
        RECT 30.535 152.955 32.145 153.155 ;
        RECT 30.535 152.945 31.370 152.955 ;
        RECT 31.960 152.865 32.145 152.955 ;
        RECT 27.765 151.155 29.435 151.925 ;
        RECT 29.605 151.665 29.775 152.855 ;
        RECT 31.475 152.755 31.805 152.785 ;
        RECT 30.005 152.695 31.805 152.755 ;
        RECT 32.395 152.695 32.650 153.315 ;
        RECT 32.825 153.270 38.170 153.705 ;
        RECT 29.945 152.585 32.650 152.695 ;
        RECT 29.945 152.550 30.145 152.585 ;
        RECT 29.945 151.975 30.115 152.550 ;
        RECT 31.475 152.525 32.650 152.585 ;
        RECT 30.345 152.110 30.755 152.415 ;
        RECT 30.925 152.145 31.255 152.355 ;
        RECT 29.945 151.855 30.215 151.975 ;
        RECT 29.945 151.810 30.790 151.855 ;
        RECT 30.035 151.685 30.790 151.810 ;
        RECT 31.045 151.745 31.255 152.145 ;
        RECT 31.500 152.145 31.975 152.355 ;
        RECT 32.165 152.145 32.655 152.345 ;
        RECT 31.500 151.745 31.720 152.145 ;
        RECT 29.605 151.655 29.835 151.665 ;
        RECT 29.605 151.325 29.865 151.655 ;
        RECT 30.620 151.535 30.790 151.685 ;
        RECT 30.035 151.155 30.365 151.515 ;
        RECT 30.620 151.325 31.920 151.535 ;
        RECT 32.195 151.155 32.650 151.920 ;
        RECT 34.410 151.700 34.750 152.530 ;
        RECT 36.230 152.020 36.580 153.270 ;
        RECT 38.345 152.615 40.935 153.705 ;
        RECT 38.345 151.925 39.555 152.445 ;
        RECT 39.725 152.095 40.935 152.615 ;
        RECT 41.575 152.735 41.905 153.535 ;
        RECT 42.075 152.905 42.305 153.705 ;
        RECT 42.475 152.735 42.805 153.535 ;
        RECT 41.575 152.565 42.805 152.735 ;
        RECT 42.975 152.565 43.230 153.705 ;
        RECT 44.325 152.565 44.605 153.705 ;
        RECT 41.565 152.065 41.875 152.395 ;
        RECT 32.825 151.155 38.170 151.700 ;
        RECT 38.345 151.155 40.935 151.925 ;
        RECT 41.575 151.665 41.905 151.895 ;
        RECT 42.080 151.835 42.455 152.395 ;
        RECT 42.625 151.665 42.805 152.565 ;
        RECT 44.775 152.555 45.105 153.535 ;
        RECT 45.275 152.565 45.535 153.705 ;
        RECT 45.705 152.615 49.215 153.705 ;
        RECT 42.990 151.815 43.210 152.395 ;
        RECT 44.335 152.125 44.670 152.395 ;
        RECT 44.840 151.955 45.010 152.555 ;
        RECT 45.180 152.145 45.515 152.395 ;
        RECT 41.575 151.325 42.805 151.665 ;
        RECT 42.975 151.155 43.230 151.645 ;
        RECT 44.325 151.155 44.635 151.955 ;
        RECT 44.840 151.325 45.535 151.955 ;
        RECT 45.705 151.925 47.355 152.445 ;
        RECT 47.525 152.095 49.215 152.615 ;
        RECT 49.845 152.540 50.135 153.705 ;
        RECT 50.305 152.615 51.975 153.705 ;
        RECT 50.305 151.925 51.055 152.445 ;
        RECT 51.225 152.095 51.975 152.615 ;
        RECT 52.645 152.755 52.935 153.525 ;
        RECT 53.505 153.165 53.765 153.525 ;
        RECT 53.935 153.335 54.265 153.705 ;
        RECT 54.435 153.165 54.695 153.525 ;
        RECT 53.505 152.935 54.695 153.165 ;
        RECT 54.885 152.985 55.215 153.705 ;
        RECT 55.385 152.755 55.650 153.525 ;
        RECT 52.645 152.575 55.140 152.755 ;
        RECT 52.615 152.065 52.885 152.395 ;
        RECT 53.065 152.065 53.500 152.395 ;
        RECT 53.680 152.065 54.255 152.395 ;
        RECT 54.435 152.065 54.715 152.395 ;
        RECT 45.705 151.155 49.215 151.925 ;
        RECT 49.845 151.155 50.135 151.880 ;
        RECT 50.305 151.155 51.975 151.925 ;
        RECT 54.915 151.885 55.140 152.575 ;
        RECT 52.655 151.695 55.140 151.885 ;
        RECT 52.655 151.335 52.880 151.695 ;
        RECT 53.060 151.155 53.390 151.525 ;
        RECT 53.570 151.335 53.825 151.695 ;
        RECT 54.390 151.155 55.135 151.525 ;
        RECT 55.315 151.335 55.650 152.755 ;
        RECT 55.825 152.615 57.035 153.705 ;
        RECT 57.385 152.790 57.555 153.705 ;
        RECT 57.725 152.645 58.055 153.490 ;
        RECT 58.225 152.695 58.395 153.705 ;
        RECT 58.565 152.975 58.905 153.535 ;
        RECT 59.135 153.205 59.450 153.705 ;
        RECT 59.630 153.235 60.515 153.405 ;
        RECT 55.825 151.905 56.345 152.445 ;
        RECT 56.515 152.075 57.035 152.615 ;
        RECT 57.665 152.565 58.055 152.645 ;
        RECT 58.565 152.600 59.460 152.975 ;
        RECT 57.665 152.515 57.880 152.565 ;
        RECT 57.665 151.935 57.835 152.515 ;
        RECT 58.565 152.395 58.755 152.600 ;
        RECT 59.630 152.395 59.800 153.235 ;
        RECT 60.740 153.205 60.990 153.535 ;
        RECT 58.005 152.065 58.755 152.395 ;
        RECT 58.925 152.065 59.800 152.395 ;
        RECT 55.825 151.155 57.035 151.905 ;
        RECT 57.665 151.895 57.890 151.935 ;
        RECT 58.555 151.895 58.755 152.065 ;
        RECT 57.665 151.810 58.045 151.895 ;
        RECT 57.375 151.155 57.545 151.670 ;
        RECT 57.715 151.375 58.045 151.810 ;
        RECT 58.215 151.155 58.385 151.765 ;
        RECT 58.555 151.370 58.885 151.895 ;
        RECT 59.145 151.155 59.355 151.685 ;
        RECT 59.630 151.605 59.800 152.065 ;
        RECT 59.970 152.105 60.290 153.065 ;
        RECT 60.460 152.315 60.650 153.035 ;
        RECT 60.820 152.135 60.990 153.205 ;
        RECT 61.160 152.905 61.330 153.705 ;
        RECT 61.500 153.260 62.605 153.430 ;
        RECT 61.500 152.645 61.670 153.260 ;
        RECT 62.815 153.110 63.065 153.535 ;
        RECT 63.235 153.245 63.500 153.705 ;
        RECT 61.840 152.725 62.370 153.090 ;
        RECT 62.815 152.980 63.120 153.110 ;
        RECT 61.160 152.555 61.670 152.645 ;
        RECT 61.160 152.385 62.030 152.555 ;
        RECT 61.160 152.315 61.330 152.385 ;
        RECT 61.450 152.135 61.650 152.165 ;
        RECT 59.970 151.775 60.435 152.105 ;
        RECT 60.820 151.835 61.650 152.135 ;
        RECT 60.820 151.605 60.990 151.835 ;
        RECT 59.630 151.435 60.415 151.605 ;
        RECT 60.585 151.435 60.990 151.605 ;
        RECT 61.170 151.155 61.540 151.655 ;
        RECT 61.860 151.605 62.030 152.385 ;
        RECT 62.200 152.025 62.370 152.725 ;
        RECT 62.540 152.195 62.780 152.790 ;
        RECT 62.200 151.805 62.725 152.025 ;
        RECT 62.950 151.875 63.120 152.980 ;
        RECT 62.895 151.745 63.120 151.875 ;
        RECT 63.290 151.785 63.570 152.735 ;
        RECT 62.895 151.605 63.065 151.745 ;
        RECT 61.860 151.435 62.535 151.605 ;
        RECT 62.730 151.435 63.065 151.605 ;
        RECT 63.235 151.155 63.485 151.615 ;
        RECT 63.740 151.415 63.925 153.535 ;
        RECT 64.095 153.205 64.425 153.705 ;
        RECT 64.595 153.035 64.765 153.535 ;
        RECT 64.100 152.865 64.765 153.035 ;
        RECT 64.100 151.875 64.330 152.865 ;
        RECT 64.500 152.045 64.850 152.695 ;
        RECT 65.025 152.565 65.315 153.705 ;
        RECT 65.485 152.985 65.935 153.535 ;
        RECT 66.125 152.985 66.455 153.705 ;
        RECT 64.100 151.705 64.765 151.875 ;
        RECT 64.095 151.155 64.425 151.535 ;
        RECT 64.595 151.415 64.765 151.705 ;
        RECT 65.025 151.155 65.315 151.955 ;
        RECT 65.485 151.615 65.735 152.985 ;
        RECT 66.665 152.815 66.965 153.365 ;
        RECT 67.135 153.035 67.415 153.705 ;
        RECT 66.025 152.645 66.965 152.815 ;
        RECT 66.025 152.395 66.195 152.645 ;
        RECT 67.300 152.395 67.615 152.835 ;
        RECT 67.785 152.615 71.295 153.705 ;
        RECT 65.905 152.065 66.195 152.395 ;
        RECT 66.365 152.145 66.695 152.395 ;
        RECT 66.925 152.145 67.615 152.395 ;
        RECT 66.025 151.975 66.195 152.065 ;
        RECT 66.025 151.785 67.415 151.975 ;
        RECT 65.485 151.325 66.035 151.615 ;
        RECT 66.205 151.155 66.455 151.615 ;
        RECT 67.085 151.425 67.415 151.785 ;
        RECT 67.785 151.925 69.435 152.445 ;
        RECT 69.605 152.095 71.295 152.615 ;
        RECT 67.785 151.155 71.295 151.925 ;
        RECT 71.935 151.335 72.195 153.525 ;
        RECT 72.365 152.975 72.705 153.705 ;
        RECT 72.885 152.795 73.155 153.525 ;
        RECT 72.385 152.575 73.155 152.795 ;
        RECT 73.335 152.815 73.565 153.525 ;
        RECT 73.735 152.995 74.065 153.705 ;
        RECT 74.235 152.815 74.495 153.525 ;
        RECT 73.335 152.575 74.495 152.815 ;
        RECT 72.385 151.905 72.675 152.575 ;
        RECT 75.605 152.540 75.895 153.705 ;
        RECT 76.125 152.565 76.335 153.705 ;
        RECT 76.505 152.555 76.835 153.535 ;
        RECT 77.005 152.565 77.235 153.705 ;
        RECT 77.445 153.195 77.745 153.705 ;
        RECT 77.915 153.025 78.245 153.535 ;
        RECT 78.415 153.195 79.045 153.705 ;
        RECT 79.625 153.195 80.005 153.365 ;
        RECT 80.175 153.195 80.475 153.705 ;
        RECT 79.835 153.025 80.005 153.195 ;
        RECT 77.445 152.855 79.665 153.025 ;
        RECT 72.855 152.085 73.320 152.395 ;
        RECT 73.500 152.085 74.025 152.395 ;
        RECT 72.385 151.705 73.615 151.905 ;
        RECT 72.455 151.155 73.125 151.525 ;
        RECT 73.305 151.335 73.615 151.705 ;
        RECT 73.795 151.445 74.025 152.085 ;
        RECT 74.205 152.065 74.505 152.395 ;
        RECT 74.205 151.155 74.495 151.885 ;
        RECT 75.605 151.155 75.895 151.880 ;
        RECT 76.125 151.155 76.335 151.975 ;
        RECT 76.505 151.955 76.755 152.555 ;
        RECT 76.925 152.145 77.255 152.395 ;
        RECT 76.505 151.325 76.835 151.955 ;
        RECT 77.005 151.155 77.235 151.975 ;
        RECT 77.445 151.895 77.615 152.855 ;
        RECT 77.785 152.515 79.325 152.685 ;
        RECT 77.785 152.065 78.030 152.515 ;
        RECT 78.290 152.145 78.985 152.345 ;
        RECT 79.155 152.315 79.325 152.515 ;
        RECT 79.495 152.655 79.665 152.855 ;
        RECT 79.835 152.825 80.495 153.025 ;
        RECT 79.495 152.485 80.155 152.655 ;
        RECT 79.155 152.145 79.755 152.315 ;
        RECT 79.985 152.065 80.155 152.485 ;
        RECT 77.445 151.350 77.910 151.895 ;
        RECT 78.415 151.155 78.585 151.975 ;
        RECT 78.755 151.895 79.665 151.975 ;
        RECT 80.325 151.895 80.495 152.825 ;
        RECT 80.665 152.615 83.255 153.705 ;
        RECT 78.755 151.805 80.005 151.895 ;
        RECT 78.755 151.325 79.085 151.805 ;
        RECT 79.495 151.725 80.005 151.805 ;
        RECT 79.255 151.155 79.605 151.545 ;
        RECT 79.775 151.325 80.005 151.725 ;
        RECT 80.175 151.415 80.495 151.895 ;
        RECT 80.665 151.925 81.875 152.445 ;
        RECT 82.045 152.095 83.255 152.615 ;
        RECT 83.895 152.735 84.225 153.535 ;
        RECT 84.395 152.905 84.625 153.705 ;
        RECT 84.795 152.735 85.125 153.535 ;
        RECT 83.895 152.565 85.125 152.735 ;
        RECT 85.295 152.565 85.550 153.705 ;
        RECT 85.735 153.095 86.065 153.525 ;
        RECT 86.245 153.265 86.440 153.705 ;
        RECT 86.610 153.095 86.940 153.525 ;
        RECT 85.735 152.925 86.940 153.095 ;
        RECT 85.735 152.595 86.630 152.925 ;
        RECT 87.110 152.755 87.385 153.525 ;
        RECT 86.800 152.565 87.385 152.755 ;
        RECT 87.565 152.615 91.075 153.705 ;
        RECT 83.885 152.065 84.195 152.395 ;
        RECT 80.665 151.155 83.255 151.925 ;
        RECT 83.895 151.665 84.225 151.895 ;
        RECT 84.400 151.835 84.775 152.395 ;
        RECT 84.945 151.665 85.125 152.565 ;
        RECT 85.310 151.815 85.530 152.395 ;
        RECT 85.740 152.065 86.035 152.395 ;
        RECT 86.215 152.065 86.630 152.395 ;
        RECT 83.895 151.325 85.125 151.665 ;
        RECT 85.295 151.155 85.550 151.645 ;
        RECT 85.735 151.155 86.035 151.885 ;
        RECT 86.215 151.445 86.445 152.065 ;
        RECT 86.800 151.895 86.975 152.565 ;
        RECT 86.645 151.715 86.975 151.895 ;
        RECT 87.145 151.745 87.385 152.395 ;
        RECT 87.565 151.925 89.215 152.445 ;
        RECT 89.385 152.095 91.075 152.615 ;
        RECT 92.165 152.565 92.505 153.535 ;
        RECT 92.675 152.565 92.845 153.705 ;
        RECT 93.115 152.905 93.365 153.705 ;
        RECT 94.010 152.735 94.340 153.535 ;
        RECT 94.640 152.905 94.970 153.705 ;
        RECT 95.140 152.735 95.470 153.535 ;
        RECT 93.035 152.565 95.470 152.735 ;
        RECT 95.845 152.565 96.120 153.535 ;
        RECT 96.330 152.905 96.610 153.705 ;
        RECT 96.780 153.195 98.830 153.485 ;
        RECT 96.780 152.855 98.410 153.025 ;
        RECT 96.780 152.735 96.950 152.855 ;
        RECT 96.290 152.565 96.950 152.735 ;
        RECT 92.165 151.955 92.340 152.565 ;
        RECT 93.035 152.315 93.205 152.565 ;
        RECT 92.510 152.145 93.205 152.315 ;
        RECT 93.380 152.145 93.800 152.345 ;
        RECT 93.970 152.145 94.300 152.345 ;
        RECT 94.470 152.145 94.800 152.345 ;
        RECT 86.645 151.335 86.870 151.715 ;
        RECT 87.040 151.155 87.370 151.545 ;
        RECT 87.565 151.155 91.075 151.925 ;
        RECT 92.165 151.325 92.505 151.955 ;
        RECT 92.675 151.155 92.925 151.955 ;
        RECT 93.115 151.805 94.340 151.975 ;
        RECT 93.115 151.325 93.445 151.805 ;
        RECT 93.615 151.155 93.840 151.615 ;
        RECT 94.010 151.325 94.340 151.805 ;
        RECT 94.970 151.935 95.140 152.565 ;
        RECT 95.325 152.145 95.675 152.395 ;
        RECT 94.970 151.325 95.470 151.935 ;
        RECT 95.845 151.830 96.015 152.565 ;
        RECT 96.290 152.395 96.460 152.565 ;
        RECT 96.185 152.065 96.460 152.395 ;
        RECT 96.630 152.065 97.010 152.395 ;
        RECT 97.180 152.065 97.920 152.685 ;
        RECT 98.090 152.565 98.410 152.855 ;
        RECT 98.605 152.395 98.845 152.990 ;
        RECT 99.015 152.630 99.355 153.705 ;
        RECT 99.525 152.615 101.195 153.705 ;
        RECT 98.190 152.065 98.845 152.395 ;
        RECT 96.290 151.895 96.460 152.065 ;
        RECT 95.845 151.485 96.120 151.830 ;
        RECT 96.290 151.725 97.875 151.895 ;
        RECT 96.310 151.155 96.690 151.555 ;
        RECT 96.860 151.375 97.030 151.725 ;
        RECT 97.200 151.155 97.530 151.555 ;
        RECT 97.705 151.375 97.875 151.725 ;
        RECT 98.075 151.155 98.405 151.655 ;
        RECT 98.600 151.375 98.845 152.065 ;
        RECT 99.015 151.825 99.355 152.395 ;
        RECT 99.525 151.925 100.275 152.445 ;
        RECT 100.445 152.095 101.195 152.615 ;
        RECT 101.365 152.540 101.655 153.705 ;
        RECT 101.835 152.895 102.130 153.705 ;
        RECT 102.310 152.395 102.555 153.535 ;
        RECT 102.730 152.895 102.990 153.705 ;
        RECT 103.590 153.700 109.865 153.705 ;
        RECT 103.170 152.395 103.420 153.530 ;
        RECT 103.590 152.905 103.850 153.700 ;
        RECT 104.020 152.805 104.280 153.530 ;
        RECT 104.450 152.975 104.710 153.700 ;
        RECT 104.880 152.805 105.140 153.530 ;
        RECT 105.310 152.975 105.570 153.700 ;
        RECT 105.740 152.805 106.000 153.530 ;
        RECT 106.170 152.975 106.430 153.700 ;
        RECT 106.600 152.805 106.860 153.530 ;
        RECT 107.030 152.975 107.275 153.700 ;
        RECT 107.445 152.805 107.705 153.530 ;
        RECT 107.890 152.975 108.135 153.700 ;
        RECT 108.305 152.805 108.565 153.530 ;
        RECT 108.750 152.975 108.995 153.700 ;
        RECT 109.165 152.805 109.425 153.530 ;
        RECT 109.610 152.975 109.865 153.700 ;
        RECT 104.020 152.790 109.425 152.805 ;
        RECT 110.035 152.790 110.325 153.530 ;
        RECT 110.495 152.960 110.765 153.705 ;
        RECT 104.020 152.565 110.765 152.790 ;
        RECT 111.085 152.645 111.415 153.490 ;
        RECT 111.585 152.695 111.755 153.705 ;
        RECT 111.925 152.975 112.265 153.535 ;
        RECT 112.495 153.205 112.810 153.705 ;
        RECT 112.990 153.235 113.875 153.405 ;
        RECT 99.015 151.155 99.355 151.655 ;
        RECT 99.525 151.155 101.195 151.925 ;
        RECT 101.365 151.155 101.655 151.880 ;
        RECT 101.825 151.835 102.140 152.395 ;
        RECT 102.310 152.145 109.430 152.395 ;
        RECT 101.825 151.155 102.130 151.665 ;
        RECT 102.310 151.335 102.560 152.145 ;
        RECT 102.730 151.155 102.990 151.680 ;
        RECT 103.170 151.335 103.420 152.145 ;
        RECT 109.600 151.975 110.765 152.565 ;
        RECT 104.020 151.805 110.765 151.975 ;
        RECT 111.025 152.565 111.415 152.645 ;
        RECT 111.925 152.600 112.820 152.975 ;
        RECT 111.025 152.515 111.240 152.565 ;
        RECT 111.025 151.935 111.195 152.515 ;
        RECT 111.925 152.395 112.115 152.600 ;
        RECT 112.990 152.395 113.160 153.235 ;
        RECT 114.100 153.205 114.350 153.535 ;
        RECT 111.365 152.065 112.115 152.395 ;
        RECT 112.285 152.065 113.160 152.395 ;
        RECT 111.025 151.895 111.250 151.935 ;
        RECT 111.915 151.895 112.115 152.065 ;
        RECT 111.025 151.810 111.405 151.895 ;
        RECT 103.590 151.155 103.850 151.715 ;
        RECT 104.020 151.350 104.280 151.805 ;
        RECT 104.450 151.155 104.710 151.635 ;
        RECT 104.880 151.350 105.140 151.805 ;
        RECT 105.310 151.155 105.570 151.635 ;
        RECT 105.740 151.350 106.000 151.805 ;
        RECT 106.170 151.155 106.415 151.635 ;
        RECT 106.585 151.350 106.860 151.805 ;
        RECT 107.030 151.155 107.275 151.635 ;
        RECT 107.445 151.350 107.705 151.805 ;
        RECT 107.885 151.155 108.135 151.635 ;
        RECT 108.305 151.350 108.565 151.805 ;
        RECT 108.745 151.155 108.995 151.635 ;
        RECT 109.165 151.350 109.425 151.805 ;
        RECT 109.605 151.155 109.865 151.635 ;
        RECT 110.035 151.350 110.295 151.805 ;
        RECT 110.465 151.155 110.765 151.635 ;
        RECT 111.075 151.375 111.405 151.810 ;
        RECT 111.575 151.155 111.745 151.765 ;
        RECT 111.915 151.370 112.245 151.895 ;
        RECT 112.505 151.155 112.715 151.685 ;
        RECT 112.990 151.605 113.160 152.065 ;
        RECT 113.330 152.105 113.650 153.065 ;
        RECT 113.820 152.315 114.010 153.035 ;
        RECT 114.180 152.135 114.350 153.205 ;
        RECT 114.520 152.905 114.690 153.705 ;
        RECT 114.860 153.260 115.965 153.430 ;
        RECT 114.860 152.645 115.030 153.260 ;
        RECT 116.175 153.110 116.425 153.535 ;
        RECT 116.595 153.245 116.860 153.705 ;
        RECT 115.200 152.725 115.730 153.090 ;
        RECT 116.175 152.980 116.480 153.110 ;
        RECT 114.520 152.555 115.030 152.645 ;
        RECT 114.520 152.385 115.390 152.555 ;
        RECT 114.520 152.315 114.690 152.385 ;
        RECT 114.810 152.135 115.010 152.165 ;
        RECT 113.330 151.775 113.795 152.105 ;
        RECT 114.180 151.835 115.010 152.135 ;
        RECT 114.180 151.605 114.350 151.835 ;
        RECT 112.990 151.435 113.775 151.605 ;
        RECT 113.945 151.435 114.350 151.605 ;
        RECT 114.530 151.155 114.900 151.655 ;
        RECT 115.220 151.605 115.390 152.385 ;
        RECT 115.560 152.025 115.730 152.725 ;
        RECT 115.900 152.195 116.140 152.790 ;
        RECT 115.560 151.805 116.085 152.025 ;
        RECT 116.310 151.875 116.480 152.980 ;
        RECT 116.255 151.745 116.480 151.875 ;
        RECT 116.650 151.785 116.930 152.735 ;
        RECT 116.255 151.605 116.425 151.745 ;
        RECT 115.220 151.435 115.895 151.605 ;
        RECT 116.090 151.435 116.425 151.605 ;
        RECT 116.595 151.155 116.845 151.615 ;
        RECT 117.100 151.415 117.285 153.535 ;
        RECT 117.455 153.205 117.785 153.705 ;
        RECT 117.955 153.035 118.125 153.535 ;
        RECT 118.385 153.270 123.730 153.705 ;
        RECT 117.460 152.865 118.125 153.035 ;
        RECT 117.460 151.875 117.690 152.865 ;
        RECT 117.860 152.045 118.210 152.695 ;
        RECT 117.460 151.705 118.125 151.875 ;
        RECT 117.455 151.155 117.785 151.535 ;
        RECT 117.955 151.415 118.125 151.705 ;
        RECT 119.970 151.700 120.310 152.530 ;
        RECT 121.790 152.020 122.140 153.270 ;
        RECT 123.905 152.615 126.495 153.705 ;
        RECT 123.905 151.925 125.115 152.445 ;
        RECT 125.285 152.095 126.495 152.615 ;
        RECT 127.125 152.540 127.415 153.705 ;
        RECT 127.585 153.270 132.930 153.705 ;
        RECT 133.105 153.270 138.450 153.705 ;
        RECT 138.625 153.270 143.970 153.705 ;
        RECT 118.385 151.155 123.730 151.700 ;
        RECT 123.905 151.155 126.495 151.925 ;
        RECT 127.125 151.155 127.415 151.880 ;
        RECT 129.170 151.700 129.510 152.530 ;
        RECT 130.990 152.020 131.340 153.270 ;
        RECT 134.690 151.700 135.030 152.530 ;
        RECT 136.510 152.020 136.860 153.270 ;
        RECT 140.210 151.700 140.550 152.530 ;
        RECT 142.030 152.020 142.380 153.270 ;
        RECT 144.145 152.615 147.655 153.705 ;
        RECT 147.825 152.615 149.035 153.705 ;
        RECT 144.145 151.925 145.795 152.445 ;
        RECT 145.965 152.095 147.655 152.615 ;
        RECT 127.585 151.155 132.930 151.700 ;
        RECT 133.105 151.155 138.450 151.700 ;
        RECT 138.625 151.155 143.970 151.700 ;
        RECT 144.145 151.155 147.655 151.925 ;
        RECT 147.825 151.905 148.345 152.445 ;
        RECT 148.515 152.075 149.035 152.615 ;
        RECT 149.205 152.615 150.415 153.705 ;
        RECT 149.205 152.075 149.725 152.615 ;
        RECT 149.895 151.905 150.415 152.445 ;
        RECT 147.825 151.155 149.035 151.905 ;
        RECT 149.205 151.155 150.415 151.905 ;
        RECT 11.120 150.985 150.500 151.155 ;
        RECT 11.205 150.235 12.415 150.985 ;
        RECT 12.585 150.440 17.930 150.985 ;
        RECT 19.025 150.525 19.585 150.815 ;
        RECT 19.755 150.525 20.005 150.985 ;
        RECT 11.205 149.695 11.725 150.235 ;
        RECT 11.895 149.525 12.415 150.065 ;
        RECT 14.170 149.610 14.510 150.440 ;
        RECT 11.205 148.435 12.415 149.525 ;
        RECT 15.990 148.870 16.340 150.120 ;
        RECT 19.025 149.155 19.275 150.525 ;
        RECT 20.625 150.355 20.955 150.715 ;
        RECT 21.325 150.440 26.670 150.985 ;
        RECT 19.565 150.165 20.955 150.355 ;
        RECT 19.565 150.075 19.735 150.165 ;
        RECT 19.445 149.745 19.735 150.075 ;
        RECT 19.905 149.745 20.245 149.995 ;
        RECT 20.465 149.745 21.140 149.995 ;
        RECT 19.565 149.495 19.735 149.745 ;
        RECT 19.565 149.325 20.505 149.495 ;
        RECT 20.875 149.385 21.140 149.745 ;
        RECT 22.910 149.610 23.250 150.440 ;
        RECT 26.845 150.215 30.355 150.985 ;
        RECT 30.525 150.235 31.735 150.985 ;
        RECT 31.905 150.245 32.225 150.725 ;
        RECT 32.395 150.415 32.625 150.815 ;
        RECT 32.795 150.595 33.145 150.985 ;
        RECT 32.395 150.335 32.905 150.415 ;
        RECT 33.315 150.335 33.645 150.815 ;
        RECT 32.395 150.245 33.645 150.335 ;
        RECT 12.585 148.435 17.930 148.870 ;
        RECT 19.025 148.605 19.485 149.155 ;
        RECT 19.675 148.435 20.005 149.155 ;
        RECT 20.205 148.775 20.505 149.325 ;
        RECT 20.675 148.435 20.955 149.105 ;
        RECT 24.730 148.870 25.080 150.120 ;
        RECT 26.845 149.695 28.495 150.215 ;
        RECT 28.665 149.525 30.355 150.045 ;
        RECT 30.525 149.695 31.045 150.235 ;
        RECT 31.215 149.525 31.735 150.065 ;
        RECT 21.325 148.435 26.670 148.870 ;
        RECT 26.845 148.435 30.355 149.525 ;
        RECT 30.525 148.435 31.735 149.525 ;
        RECT 31.905 149.315 32.075 150.245 ;
        RECT 32.735 150.165 33.645 150.245 ;
        RECT 33.815 150.165 33.985 150.985 ;
        RECT 34.490 150.245 34.955 150.790 ;
        RECT 32.245 149.655 32.415 150.075 ;
        RECT 32.645 149.825 33.245 149.995 ;
        RECT 32.245 149.485 32.905 149.655 ;
        RECT 31.905 149.115 32.565 149.315 ;
        RECT 32.735 149.285 32.905 149.485 ;
        RECT 33.075 149.625 33.245 149.825 ;
        RECT 33.415 149.795 34.110 149.995 ;
        RECT 34.370 149.625 34.615 150.075 ;
        RECT 33.075 149.455 34.615 149.625 ;
        RECT 34.785 149.285 34.955 150.245 ;
        RECT 35.125 150.215 36.795 150.985 ;
        RECT 36.965 150.260 37.255 150.985 ;
        RECT 37.425 150.235 38.635 150.985 ;
        RECT 35.125 149.695 35.875 150.215 ;
        RECT 36.045 149.525 36.795 150.045 ;
        RECT 37.425 149.695 37.945 150.235 ;
        RECT 38.805 150.185 39.115 150.985 ;
        RECT 39.320 150.185 40.015 150.815 ;
        RECT 41.105 150.185 41.415 150.985 ;
        RECT 41.620 150.185 42.315 150.815 ;
        RECT 42.485 150.440 47.830 150.985 ;
        RECT 39.320 150.135 39.495 150.185 ;
        RECT 32.735 149.115 34.955 149.285 ;
        RECT 32.395 148.945 32.565 149.115 ;
        RECT 31.925 148.435 32.225 148.945 ;
        RECT 32.395 148.775 32.775 148.945 ;
        RECT 33.355 148.435 33.985 148.945 ;
        RECT 34.155 148.605 34.485 149.115 ;
        RECT 34.655 148.435 34.955 148.945 ;
        RECT 35.125 148.435 36.795 149.525 ;
        RECT 36.965 148.435 37.255 149.600 ;
        RECT 38.115 149.525 38.635 150.065 ;
        RECT 38.815 149.745 39.150 150.015 ;
        RECT 39.320 149.585 39.490 150.135 ;
        RECT 39.660 149.745 39.995 149.995 ;
        RECT 41.115 149.745 41.450 150.015 ;
        RECT 41.620 149.585 41.790 150.185 ;
        RECT 41.960 149.745 42.295 149.995 ;
        RECT 44.070 149.610 44.410 150.440 ;
        RECT 48.005 150.215 50.595 150.985 ;
        RECT 37.425 148.435 38.635 149.525 ;
        RECT 38.805 148.435 39.085 149.575 ;
        RECT 39.255 148.605 39.585 149.585 ;
        RECT 39.755 148.435 40.015 149.575 ;
        RECT 41.105 148.435 41.385 149.575 ;
        RECT 41.555 148.605 41.885 149.585 ;
        RECT 42.055 148.435 42.315 149.575 ;
        RECT 45.890 148.870 46.240 150.120 ;
        RECT 48.005 149.695 49.215 150.215 ;
        RECT 49.385 149.525 50.595 150.045 ;
        RECT 42.485 148.435 47.830 148.870 ;
        RECT 48.005 148.435 50.595 149.525 ;
        RECT 51.245 149.405 51.475 150.745 ;
        RECT 51.655 149.905 51.885 150.805 ;
        RECT 52.085 150.205 52.330 150.985 ;
        RECT 52.500 150.445 52.930 150.805 ;
        RECT 53.510 150.615 54.240 150.985 ;
        RECT 52.500 150.255 54.240 150.445 ;
        RECT 52.500 150.025 52.720 150.255 ;
        RECT 51.655 149.225 51.995 149.905 ;
        RECT 51.245 149.025 51.995 149.225 ;
        RECT 52.175 149.725 52.720 150.025 ;
        RECT 51.245 148.635 51.485 149.025 ;
        RECT 51.655 148.435 52.005 148.845 ;
        RECT 52.175 148.615 52.505 149.725 ;
        RECT 52.890 149.455 53.315 150.075 ;
        RECT 53.510 149.455 53.770 150.075 ;
        RECT 53.980 149.745 54.240 150.255 ;
        RECT 52.675 149.085 53.700 149.285 ;
        RECT 52.675 148.615 52.855 149.085 ;
        RECT 53.025 148.435 53.355 148.915 ;
        RECT 53.530 148.615 53.700 149.085 ;
        RECT 53.965 148.435 54.250 149.575 ;
        RECT 54.440 148.615 54.720 150.805 ;
        RECT 54.905 150.440 60.250 150.985 ;
        RECT 56.490 149.610 56.830 150.440 ;
        RECT 60.425 150.215 62.095 150.985 ;
        RECT 62.725 150.260 63.015 150.985 ;
        RECT 63.185 150.440 68.530 150.985 ;
        RECT 68.705 150.440 74.050 150.985 ;
        RECT 74.775 150.645 74.945 150.680 ;
        RECT 74.745 150.475 74.945 150.645 ;
        RECT 58.310 148.870 58.660 150.120 ;
        RECT 60.425 149.695 61.175 150.215 ;
        RECT 61.345 149.525 62.095 150.045 ;
        RECT 64.770 149.610 65.110 150.440 ;
        RECT 54.905 148.435 60.250 148.870 ;
        RECT 60.425 148.435 62.095 149.525 ;
        RECT 62.725 148.435 63.015 149.600 ;
        RECT 66.590 148.870 66.940 150.120 ;
        RECT 70.290 149.610 70.630 150.440 ;
        RECT 72.110 148.870 72.460 150.120 ;
        RECT 74.775 150.115 74.945 150.475 ;
        RECT 75.135 150.455 75.365 150.760 ;
        RECT 75.535 150.625 75.865 150.985 ;
        RECT 76.060 150.455 76.350 150.805 ;
        RECT 75.135 150.285 76.350 150.455 ;
        RECT 76.525 150.440 81.870 150.985 ;
        RECT 82.045 150.440 87.390 150.985 ;
        RECT 74.775 149.945 75.295 150.115 ;
        RECT 74.690 149.415 74.935 149.775 ;
        RECT 75.125 149.565 75.295 149.945 ;
        RECT 75.465 149.745 75.850 150.075 ;
        RECT 76.030 149.965 76.290 150.075 ;
        RECT 76.030 149.795 76.295 149.965 ;
        RECT 76.030 149.745 76.290 149.795 ;
        RECT 75.125 149.285 75.475 149.565 ;
        RECT 63.185 148.435 68.530 148.870 ;
        RECT 68.705 148.435 74.050 148.870 ;
        RECT 74.690 148.435 74.945 149.235 ;
        RECT 75.145 148.605 75.475 149.285 ;
        RECT 75.655 148.695 75.850 149.745 ;
        RECT 78.110 149.610 78.450 150.440 ;
        RECT 76.030 148.435 76.350 149.575 ;
        RECT 79.930 148.870 80.280 150.120 ;
        RECT 83.630 149.610 83.970 150.440 ;
        RECT 88.485 150.260 88.775 150.985 ;
        RECT 88.945 150.215 92.455 150.985 ;
        RECT 93.175 150.335 93.345 150.815 ;
        RECT 93.515 150.505 93.845 150.985 ;
        RECT 94.070 150.565 95.605 150.815 ;
        RECT 94.070 150.335 94.240 150.565 ;
        RECT 85.450 148.870 85.800 150.120 ;
        RECT 88.945 149.695 90.595 150.215 ;
        RECT 93.175 150.165 94.240 150.335 ;
        RECT 76.525 148.435 81.870 148.870 ;
        RECT 82.045 148.435 87.390 148.870 ;
        RECT 88.485 148.435 88.775 149.600 ;
        RECT 90.765 149.525 92.455 150.045 ;
        RECT 94.420 149.995 94.700 150.395 ;
        RECT 93.090 149.785 93.440 149.995 ;
        RECT 93.610 149.795 94.055 149.995 ;
        RECT 94.225 149.795 94.700 149.995 ;
        RECT 94.970 149.995 95.255 150.395 ;
        RECT 95.435 150.335 95.605 150.565 ;
        RECT 95.775 150.505 96.105 150.985 ;
        RECT 96.320 150.485 96.575 150.815 ;
        RECT 96.365 150.475 96.575 150.485 ;
        RECT 96.390 150.405 96.575 150.475 ;
        RECT 95.435 150.165 96.235 150.335 ;
        RECT 94.970 149.795 95.300 149.995 ;
        RECT 95.470 149.795 95.835 149.995 ;
        RECT 96.065 149.615 96.235 150.165 ;
        RECT 88.945 148.435 92.455 149.525 ;
        RECT 93.175 149.445 96.235 149.615 ;
        RECT 93.175 148.605 93.345 149.445 ;
        RECT 96.405 149.275 96.575 150.405 ;
        RECT 96.855 150.115 97.025 150.680 ;
        RECT 97.215 150.455 97.445 150.760 ;
        RECT 97.615 150.625 97.945 150.985 ;
        RECT 98.140 150.455 98.430 150.805 ;
        RECT 97.215 150.285 98.430 150.455 ;
        RECT 98.605 150.215 101.195 150.985 ;
        RECT 96.855 149.945 97.375 150.115 ;
        RECT 96.770 149.415 97.015 149.775 ;
        RECT 97.205 149.565 97.375 149.945 ;
        RECT 97.545 149.745 97.930 150.075 ;
        RECT 98.110 149.965 98.370 150.075 ;
        RECT 98.110 149.795 98.375 149.965 ;
        RECT 98.110 149.745 98.370 149.795 ;
        RECT 97.205 149.285 97.555 149.565 ;
        RECT 93.515 148.775 93.845 149.275 ;
        RECT 94.015 149.035 95.650 149.275 ;
        RECT 94.015 148.945 94.245 149.035 ;
        RECT 94.355 148.775 94.685 148.815 ;
        RECT 93.515 148.605 94.685 148.775 ;
        RECT 94.875 148.435 95.230 148.855 ;
        RECT 95.400 148.605 95.650 149.035 ;
        RECT 95.820 148.435 96.150 149.195 ;
        RECT 96.320 148.605 96.575 149.275 ;
        RECT 96.770 148.435 97.025 149.235 ;
        RECT 97.225 148.605 97.555 149.285 ;
        RECT 97.735 148.695 97.930 149.745 ;
        RECT 98.605 149.695 99.815 150.215 ;
        RECT 101.825 150.150 102.115 150.985 ;
        RECT 102.285 150.585 103.240 150.755 ;
        RECT 103.655 150.595 103.985 150.985 ;
        RECT 98.110 148.435 98.430 149.575 ;
        RECT 99.985 149.525 101.195 150.045 ;
        RECT 102.285 149.705 102.455 150.585 ;
        RECT 104.155 150.415 104.325 150.735 ;
        RECT 104.495 150.595 104.825 150.985 ;
        RECT 102.625 150.245 104.875 150.415 ;
        RECT 102.625 149.745 102.855 150.245 ;
        RECT 103.025 149.825 103.400 149.995 ;
        RECT 98.605 148.435 101.195 149.525 ;
        RECT 101.825 149.535 102.455 149.705 ;
        RECT 103.230 149.625 103.400 149.825 ;
        RECT 103.570 149.795 104.120 149.995 ;
        RECT 104.290 149.625 104.535 150.075 ;
        RECT 101.825 148.605 102.145 149.535 ;
        RECT 103.230 149.455 104.535 149.625 ;
        RECT 104.705 149.285 104.875 150.245 ;
        RECT 106.170 150.205 106.670 150.815 ;
        RECT 105.965 149.745 106.315 149.995 ;
        RECT 106.500 149.575 106.670 150.205 ;
        RECT 107.300 150.335 107.630 150.815 ;
        RECT 107.800 150.525 108.025 150.985 ;
        RECT 108.195 150.335 108.525 150.815 ;
        RECT 107.300 150.165 108.525 150.335 ;
        RECT 108.715 150.185 108.965 150.985 ;
        RECT 109.135 150.185 109.475 150.815 ;
        RECT 109.655 150.645 110.845 150.815 ;
        RECT 109.655 150.475 109.965 150.645 ;
        RECT 106.840 149.795 107.170 149.995 ;
        RECT 107.340 149.795 107.670 149.995 ;
        RECT 107.840 149.795 108.260 149.995 ;
        RECT 108.435 149.825 109.130 149.995 ;
        RECT 108.435 149.575 108.605 149.825 ;
        RECT 109.300 149.575 109.475 150.185 ;
        RECT 109.650 149.670 109.965 150.305 ;
        RECT 102.325 149.115 103.565 149.285 ;
        RECT 102.325 148.605 102.725 149.115 ;
        RECT 102.895 148.435 103.065 148.945 ;
        RECT 103.235 148.605 103.565 149.115 ;
        RECT 103.735 148.435 103.905 149.285 ;
        RECT 104.495 148.605 104.875 149.285 ;
        RECT 106.170 149.405 108.605 149.575 ;
        RECT 106.170 148.605 106.500 149.405 ;
        RECT 106.670 148.435 107.000 149.235 ;
        RECT 107.300 148.605 107.630 149.405 ;
        RECT 108.275 148.435 108.525 149.235 ;
        RECT 108.795 148.435 108.965 149.575 ;
        RECT 109.135 148.605 109.475 149.575 ;
        RECT 109.655 148.435 109.965 149.500 ;
        RECT 110.135 149.285 110.345 150.475 ;
        RECT 110.515 150.355 110.845 150.645 ;
        RECT 111.085 150.525 111.255 150.985 ;
        RECT 111.485 150.355 111.815 150.815 ;
        RECT 111.995 150.525 112.165 150.985 ;
        RECT 112.345 150.355 112.675 150.815 ;
        RECT 110.515 150.185 112.675 150.355 ;
        RECT 112.905 150.165 113.135 150.985 ;
        RECT 113.305 150.185 113.635 150.815 ;
        RECT 110.685 149.625 111.180 149.995 ;
        RECT 111.360 149.795 112.160 149.995 ;
        RECT 112.330 149.625 112.660 150.015 ;
        RECT 112.885 149.745 113.215 149.995 ;
        RECT 110.625 149.455 112.660 149.625 ;
        RECT 113.385 149.585 113.635 150.185 ;
        RECT 113.805 150.165 114.015 150.985 ;
        RECT 114.245 150.260 114.535 150.985 ;
        RECT 114.795 150.435 114.965 150.815 ;
        RECT 115.145 150.605 115.475 150.985 ;
        RECT 114.795 150.265 115.460 150.435 ;
        RECT 115.655 150.310 115.915 150.815 ;
        RECT 116.255 150.470 116.425 150.985 ;
        RECT 116.595 150.330 116.925 150.765 ;
        RECT 117.095 150.375 117.265 150.985 ;
        RECT 114.725 149.715 115.055 150.085 ;
        RECT 115.290 150.010 115.460 150.265 ;
        RECT 115.290 149.680 115.575 150.010 ;
        RECT 110.135 149.105 111.785 149.285 ;
        RECT 110.135 148.605 110.370 149.105 ;
        RECT 111.485 148.945 111.785 149.105 ;
        RECT 110.540 148.435 110.870 148.895 ;
        RECT 111.065 148.775 111.255 148.935 ;
        RECT 111.955 148.775 112.175 149.285 ;
        RECT 111.065 148.605 112.175 148.775 ;
        RECT 112.345 148.435 112.675 149.285 ;
        RECT 112.905 148.435 113.135 149.575 ;
        RECT 113.305 148.605 113.635 149.585 ;
        RECT 113.805 148.435 114.015 149.575 ;
        RECT 114.245 148.435 114.535 149.600 ;
        RECT 115.290 149.535 115.460 149.680 ;
        RECT 114.795 149.365 115.460 149.535 ;
        RECT 115.745 149.510 115.915 150.310 ;
        RECT 114.795 148.605 114.965 149.365 ;
        RECT 115.145 148.435 115.475 149.195 ;
        RECT 115.645 148.605 115.915 149.510 ;
        RECT 116.545 150.245 116.925 150.330 ;
        RECT 117.435 150.245 117.765 150.770 ;
        RECT 118.025 150.455 118.235 150.985 ;
        RECT 118.510 150.535 119.295 150.705 ;
        RECT 119.465 150.535 119.870 150.705 ;
        RECT 116.545 150.205 116.770 150.245 ;
        RECT 116.545 149.625 116.715 150.205 ;
        RECT 117.435 150.075 117.635 150.245 ;
        RECT 118.510 150.075 118.680 150.535 ;
        RECT 116.885 149.745 117.635 150.075 ;
        RECT 117.805 149.745 118.680 150.075 ;
        RECT 116.545 149.575 116.760 149.625 ;
        RECT 116.545 149.495 116.935 149.575 ;
        RECT 116.265 148.435 116.435 149.350 ;
        RECT 116.605 148.650 116.935 149.495 ;
        RECT 117.445 149.540 117.635 149.745 ;
        RECT 117.105 148.435 117.275 149.445 ;
        RECT 117.445 149.165 118.340 149.540 ;
        RECT 117.445 148.605 117.785 149.165 ;
        RECT 118.015 148.435 118.330 148.935 ;
        RECT 118.510 148.905 118.680 149.745 ;
        RECT 118.850 150.035 119.315 150.365 ;
        RECT 119.700 150.305 119.870 150.535 ;
        RECT 120.050 150.485 120.420 150.985 ;
        RECT 120.740 150.535 121.415 150.705 ;
        RECT 121.610 150.535 121.945 150.705 ;
        RECT 118.850 149.075 119.170 150.035 ;
        RECT 119.700 150.005 120.530 150.305 ;
        RECT 119.340 149.105 119.530 149.825 ;
        RECT 119.700 148.935 119.870 150.005 ;
        RECT 120.330 149.975 120.530 150.005 ;
        RECT 120.040 149.755 120.210 149.825 ;
        RECT 120.740 149.755 120.910 150.535 ;
        RECT 121.775 150.395 121.945 150.535 ;
        RECT 122.115 150.525 122.365 150.985 ;
        RECT 120.040 149.585 120.910 149.755 ;
        RECT 121.080 150.115 121.605 150.335 ;
        RECT 121.775 150.265 122.000 150.395 ;
        RECT 120.040 149.495 120.550 149.585 ;
        RECT 118.510 148.735 119.395 148.905 ;
        RECT 119.620 148.605 119.870 148.935 ;
        RECT 120.040 148.435 120.210 149.235 ;
        RECT 120.380 148.880 120.550 149.495 ;
        RECT 121.080 149.415 121.250 150.115 ;
        RECT 120.720 149.050 121.250 149.415 ;
        RECT 121.420 149.350 121.660 149.945 ;
        RECT 121.830 149.160 122.000 150.265 ;
        RECT 122.170 149.405 122.450 150.355 ;
        RECT 121.695 149.030 122.000 149.160 ;
        RECT 120.380 148.710 121.485 148.880 ;
        RECT 121.695 148.605 121.945 149.030 ;
        RECT 122.115 148.435 122.380 148.895 ;
        RECT 122.620 148.605 122.805 150.725 ;
        RECT 122.975 150.605 123.305 150.985 ;
        RECT 123.475 150.435 123.645 150.725 ;
        RECT 123.905 150.440 129.250 150.985 ;
        RECT 129.425 150.440 134.770 150.985 ;
        RECT 122.980 150.265 123.645 150.435 ;
        RECT 122.980 149.275 123.210 150.265 ;
        RECT 123.380 149.445 123.730 150.095 ;
        RECT 125.490 149.610 125.830 150.440 ;
        RECT 122.980 149.105 123.645 149.275 ;
        RECT 122.975 148.435 123.305 148.935 ;
        RECT 123.475 148.605 123.645 149.105 ;
        RECT 127.310 148.870 127.660 150.120 ;
        RECT 131.010 149.610 131.350 150.440 ;
        RECT 134.945 150.215 138.455 150.985 ;
        RECT 138.625 150.235 139.835 150.985 ;
        RECT 140.005 150.260 140.295 150.985 ;
        RECT 140.465 150.440 145.810 150.985 ;
        RECT 132.830 148.870 133.180 150.120 ;
        RECT 134.945 149.695 136.595 150.215 ;
        RECT 136.765 149.525 138.455 150.045 ;
        RECT 138.625 149.695 139.145 150.235 ;
        RECT 139.315 149.525 139.835 150.065 ;
        RECT 142.050 149.610 142.390 150.440 ;
        RECT 145.985 150.215 148.575 150.985 ;
        RECT 149.205 150.235 150.415 150.985 ;
        RECT 123.905 148.435 129.250 148.870 ;
        RECT 129.425 148.435 134.770 148.870 ;
        RECT 134.945 148.435 138.455 149.525 ;
        RECT 138.625 148.435 139.835 149.525 ;
        RECT 140.005 148.435 140.295 149.600 ;
        RECT 143.870 148.870 144.220 150.120 ;
        RECT 145.985 149.695 147.195 150.215 ;
        RECT 147.365 149.525 148.575 150.045 ;
        RECT 140.465 148.435 145.810 148.870 ;
        RECT 145.985 148.435 148.575 149.525 ;
        RECT 149.205 149.525 149.725 150.065 ;
        RECT 149.895 149.695 150.415 150.235 ;
        RECT 149.205 148.435 150.415 149.525 ;
        RECT 11.120 148.265 150.500 148.435 ;
        RECT 11.205 147.175 12.415 148.265 ;
        RECT 12.585 147.830 17.930 148.265 ;
        RECT 11.205 146.465 11.725 147.005 ;
        RECT 11.895 146.635 12.415 147.175 ;
        RECT 11.205 145.715 12.415 146.465 ;
        RECT 14.170 146.260 14.510 147.090 ;
        RECT 15.990 146.580 16.340 147.830 ;
        RECT 18.655 147.645 18.825 148.075 ;
        RECT 18.995 147.815 19.325 148.265 ;
        RECT 18.655 147.415 19.330 147.645 ;
        RECT 18.625 146.395 18.925 147.245 ;
        RECT 19.095 146.765 19.330 147.415 ;
        RECT 19.500 147.105 19.785 148.050 ;
        RECT 19.965 147.795 20.650 148.265 ;
        RECT 19.960 147.275 20.655 147.585 ;
        RECT 20.830 147.210 21.135 147.995 ;
        RECT 21.415 147.645 21.585 148.075 ;
        RECT 21.755 147.815 22.085 148.265 ;
        RECT 21.415 147.415 22.090 147.645 ;
        RECT 19.500 146.955 20.360 147.105 ;
        RECT 20.925 147.075 21.135 147.210 ;
        RECT 19.500 146.935 20.785 146.955 ;
        RECT 19.095 146.435 19.630 146.765 ;
        RECT 19.800 146.575 20.785 146.935 ;
        RECT 19.095 146.285 19.315 146.435 ;
        RECT 12.585 145.715 17.930 146.260 ;
        RECT 18.570 145.715 18.905 146.220 ;
        RECT 19.075 145.910 19.315 146.285 ;
        RECT 19.800 146.240 19.970 146.575 ;
        RECT 20.960 146.405 21.135 147.075 ;
        RECT 19.595 146.045 19.970 146.240 ;
        RECT 19.595 145.900 19.765 146.045 ;
        RECT 20.330 145.715 20.725 146.210 ;
        RECT 20.895 145.885 21.135 146.405 ;
        RECT 21.385 146.395 21.685 147.245 ;
        RECT 21.855 146.765 22.090 147.415 ;
        RECT 22.260 147.105 22.545 148.050 ;
        RECT 22.725 147.795 23.410 148.265 ;
        RECT 22.720 147.275 23.415 147.585 ;
        RECT 23.590 147.210 23.895 147.995 ;
        RECT 22.260 146.955 23.120 147.105 ;
        RECT 22.260 146.935 23.545 146.955 ;
        RECT 21.855 146.435 22.390 146.765 ;
        RECT 22.560 146.575 23.545 146.935 ;
        RECT 21.855 146.285 22.075 146.435 ;
        RECT 21.330 145.715 21.665 146.220 ;
        RECT 21.835 145.910 22.075 146.285 ;
        RECT 22.560 146.240 22.730 146.575 ;
        RECT 23.720 146.405 23.895 147.210 ;
        RECT 24.085 147.100 24.375 148.265 ;
        RECT 24.555 147.125 24.885 148.265 ;
        RECT 25.415 147.295 25.745 148.080 ;
        RECT 26.225 147.625 26.555 148.055 ;
        RECT 25.065 147.125 25.745 147.295 ;
        RECT 26.100 147.455 26.555 147.625 ;
        RECT 26.735 147.625 26.985 148.045 ;
        RECT 27.215 147.795 27.545 148.265 ;
        RECT 27.775 147.625 28.025 148.045 ;
        RECT 26.735 147.455 28.025 147.625 ;
        RECT 24.545 146.705 24.895 146.955 ;
        RECT 25.065 146.525 25.235 147.125 ;
        RECT 25.405 146.705 25.755 146.955 ;
        RECT 22.355 146.045 22.730 146.240 ;
        RECT 22.355 145.900 22.525 146.045 ;
        RECT 23.090 145.715 23.485 146.210 ;
        RECT 23.655 145.885 23.895 146.405 ;
        RECT 24.085 145.715 24.375 146.440 ;
        RECT 24.555 145.715 24.825 146.525 ;
        RECT 24.995 145.885 25.325 146.525 ;
        RECT 25.495 145.715 25.735 146.525 ;
        RECT 26.100 146.455 26.270 147.455 ;
        RECT 26.440 146.625 26.685 147.285 ;
        RECT 26.900 146.625 27.165 147.285 ;
        RECT 27.360 146.625 27.645 147.285 ;
        RECT 27.820 146.955 28.035 147.285 ;
        RECT 28.215 147.125 28.465 148.265 ;
        RECT 28.635 147.205 28.965 148.055 ;
        RECT 27.820 146.625 28.125 146.955 ;
        RECT 28.295 146.625 28.605 146.955 ;
        RECT 28.295 146.455 28.465 146.625 ;
        RECT 26.100 146.285 28.465 146.455 ;
        RECT 28.775 146.440 28.965 147.205 ;
        RECT 26.255 145.715 26.585 146.115 ;
        RECT 26.755 145.945 27.085 146.285 ;
        RECT 28.135 145.715 28.465 146.115 ;
        RECT 28.635 145.930 28.965 146.440 ;
        RECT 29.145 147.110 29.485 148.095 ;
        RECT 29.655 147.835 30.065 148.265 ;
        RECT 30.810 147.845 31.140 148.265 ;
        RECT 31.310 147.665 31.635 148.095 ;
        RECT 29.655 147.495 31.635 147.665 ;
        RECT 29.145 146.455 29.400 147.110 ;
        RECT 29.655 146.955 29.920 147.495 ;
        RECT 30.135 147.155 30.760 147.325 ;
        RECT 29.570 146.625 29.920 146.955 ;
        RECT 30.090 146.625 30.420 146.955 ;
        RECT 30.590 146.455 30.760 147.155 ;
        RECT 29.145 146.080 29.505 146.455 ;
        RECT 29.770 145.715 29.940 146.455 ;
        RECT 30.220 146.285 30.760 146.455 ;
        RECT 30.930 147.085 31.635 147.495 ;
        RECT 32.110 147.165 32.440 148.265 ;
        RECT 32.825 147.175 36.335 148.265 ;
        RECT 36.505 147.175 37.715 148.265 ;
        RECT 37.975 147.595 38.145 148.095 ;
        RECT 38.315 147.765 38.645 148.265 ;
        RECT 37.975 147.425 38.640 147.595 ;
        RECT 30.220 146.080 30.390 146.285 ;
        RECT 30.930 145.885 31.100 147.085 ;
        RECT 31.270 146.705 31.840 146.915 ;
        RECT 32.010 146.705 32.655 146.915 ;
        RECT 31.330 146.365 32.500 146.535 ;
        RECT 31.330 145.885 31.660 146.365 ;
        RECT 31.830 145.715 32.000 146.185 ;
        RECT 32.170 145.900 32.500 146.365 ;
        RECT 32.825 146.485 34.475 147.005 ;
        RECT 34.645 146.655 36.335 147.175 ;
        RECT 32.825 145.715 36.335 146.485 ;
        RECT 36.505 146.465 37.025 147.005 ;
        RECT 37.195 146.635 37.715 147.175 ;
        RECT 37.890 146.605 38.240 147.255 ;
        RECT 36.505 145.715 37.715 146.465 ;
        RECT 38.410 146.435 38.640 147.425 ;
        RECT 37.975 146.265 38.640 146.435 ;
        RECT 37.975 145.975 38.145 146.265 ;
        RECT 38.315 145.715 38.645 146.095 ;
        RECT 38.815 145.975 39.000 148.095 ;
        RECT 39.240 147.805 39.505 148.265 ;
        RECT 39.675 147.670 39.925 148.095 ;
        RECT 40.135 147.820 41.240 147.990 ;
        RECT 39.620 147.540 39.925 147.670 ;
        RECT 39.170 146.345 39.450 147.295 ;
        RECT 39.620 146.435 39.790 147.540 ;
        RECT 39.960 146.755 40.200 147.350 ;
        RECT 40.370 147.285 40.900 147.650 ;
        RECT 40.370 146.585 40.540 147.285 ;
        RECT 41.070 147.205 41.240 147.820 ;
        RECT 41.410 147.465 41.580 148.265 ;
        RECT 41.750 147.765 42.000 148.095 ;
        RECT 42.225 147.795 43.110 147.965 ;
        RECT 41.070 147.115 41.580 147.205 ;
        RECT 39.620 146.305 39.845 146.435 ;
        RECT 40.015 146.365 40.540 146.585 ;
        RECT 40.710 146.945 41.580 147.115 ;
        RECT 39.255 145.715 39.505 146.175 ;
        RECT 39.675 146.165 39.845 146.305 ;
        RECT 40.710 146.165 40.880 146.945 ;
        RECT 41.410 146.875 41.580 146.945 ;
        RECT 41.090 146.695 41.290 146.725 ;
        RECT 41.750 146.695 41.920 147.765 ;
        RECT 42.090 146.875 42.280 147.595 ;
        RECT 41.090 146.395 41.920 146.695 ;
        RECT 42.450 146.665 42.770 147.625 ;
        RECT 39.675 145.995 40.010 146.165 ;
        RECT 40.205 145.995 40.880 146.165 ;
        RECT 41.200 145.715 41.570 146.215 ;
        RECT 41.750 146.165 41.920 146.395 ;
        RECT 42.305 146.335 42.770 146.665 ;
        RECT 42.940 146.955 43.110 147.795 ;
        RECT 43.290 147.765 43.605 148.265 ;
        RECT 43.835 147.535 44.175 148.095 ;
        RECT 43.280 147.160 44.175 147.535 ;
        RECT 44.345 147.255 44.515 148.265 ;
        RECT 43.985 146.955 44.175 147.160 ;
        RECT 44.685 147.205 45.015 148.050 ;
        RECT 45.740 147.475 46.275 148.095 ;
        RECT 44.685 147.125 45.075 147.205 ;
        RECT 44.860 147.075 45.075 147.125 ;
        RECT 42.940 146.625 43.815 146.955 ;
        RECT 43.985 146.625 44.735 146.955 ;
        RECT 42.940 146.165 43.110 146.625 ;
        RECT 43.985 146.455 44.185 146.625 ;
        RECT 44.905 146.495 45.075 147.075 ;
        RECT 44.850 146.455 45.075 146.495 ;
        RECT 41.750 145.995 42.155 146.165 ;
        RECT 42.325 145.995 43.110 146.165 ;
        RECT 43.385 145.715 43.595 146.245 ;
        RECT 43.855 145.930 44.185 146.455 ;
        RECT 44.695 146.370 45.075 146.455 ;
        RECT 45.740 146.455 46.055 147.475 ;
        RECT 46.445 147.465 46.775 148.265 ;
        RECT 47.260 147.295 47.650 147.470 ;
        RECT 46.225 147.125 47.650 147.295 ;
        RECT 48.095 147.335 48.265 148.095 ;
        RECT 48.480 147.505 48.810 148.265 ;
        RECT 48.095 147.165 48.810 147.335 ;
        RECT 48.980 147.190 49.235 148.095 ;
        RECT 46.225 146.625 46.395 147.125 ;
        RECT 44.355 145.715 44.525 146.325 ;
        RECT 44.695 145.935 45.025 146.370 ;
        RECT 45.740 145.885 46.355 146.455 ;
        RECT 46.645 146.395 46.910 146.955 ;
        RECT 47.080 146.225 47.250 147.125 ;
        RECT 47.420 146.395 47.775 146.955 ;
        RECT 48.005 146.615 48.360 146.985 ;
        RECT 48.640 146.955 48.810 147.165 ;
        RECT 48.640 146.625 48.895 146.955 ;
        RECT 48.640 146.435 48.810 146.625 ;
        RECT 49.065 146.460 49.235 147.190 ;
        RECT 49.410 147.115 49.670 148.265 ;
        RECT 49.845 147.100 50.135 148.265 ;
        RECT 50.775 147.125 51.105 148.265 ;
        RECT 51.635 147.295 51.965 148.080 ;
        RECT 52.155 147.545 52.485 148.265 ;
        RECT 51.285 147.125 51.965 147.295 ;
        RECT 50.765 146.705 51.115 146.955 ;
        RECT 48.095 146.265 48.810 146.435 ;
        RECT 46.525 145.715 46.740 146.225 ;
        RECT 46.970 145.895 47.250 146.225 ;
        RECT 47.430 145.715 47.670 146.225 ;
        RECT 48.095 145.885 48.265 146.265 ;
        RECT 48.480 145.715 48.810 146.095 ;
        RECT 48.980 145.885 49.235 146.460 ;
        RECT 49.410 145.715 49.670 146.555 ;
        RECT 51.285 146.525 51.455 147.125 ;
        RECT 51.625 146.705 51.975 146.955 ;
        RECT 52.145 146.905 52.375 147.245 ;
        RECT 52.665 146.905 52.880 148.020 ;
        RECT 53.075 147.320 53.405 148.095 ;
        RECT 53.575 147.490 54.285 148.265 ;
        RECT 53.075 147.105 54.225 147.320 ;
        RECT 52.145 146.705 52.475 146.905 ;
        RECT 52.665 146.725 53.115 146.905 ;
        RECT 52.785 146.705 53.115 146.725 ;
        RECT 53.285 146.705 53.755 146.935 ;
        RECT 53.940 146.535 54.225 147.105 ;
        RECT 54.455 146.660 54.735 148.095 ;
        RECT 49.845 145.715 50.135 146.440 ;
        RECT 50.775 145.715 51.045 146.525 ;
        RECT 51.215 145.885 51.545 146.525 ;
        RECT 51.715 145.715 51.955 146.525 ;
        RECT 52.145 146.345 53.325 146.535 ;
        RECT 52.145 145.885 52.485 146.345 ;
        RECT 52.995 146.265 53.325 146.345 ;
        RECT 53.515 146.345 54.225 146.535 ;
        RECT 53.515 146.205 53.815 146.345 ;
        RECT 53.500 146.195 53.815 146.205 ;
        RECT 53.490 146.185 53.815 146.195 ;
        RECT 53.480 146.180 53.815 146.185 ;
        RECT 52.655 145.715 52.825 146.175 ;
        RECT 53.475 146.170 53.815 146.180 ;
        RECT 53.470 146.165 53.815 146.170 ;
        RECT 53.465 146.155 53.815 146.165 ;
        RECT 53.460 146.150 53.815 146.155 ;
        RECT 53.455 145.885 53.815 146.150 ;
        RECT 54.055 145.715 54.225 146.175 ;
        RECT 54.395 145.885 54.735 146.660 ;
        RECT 55.825 147.415 56.205 148.095 ;
        RECT 56.795 147.415 56.965 148.265 ;
        RECT 57.135 147.585 57.465 148.095 ;
        RECT 57.635 147.755 57.805 148.265 ;
        RECT 57.975 147.585 58.375 148.095 ;
        RECT 57.135 147.415 58.375 147.585 ;
        RECT 55.825 146.455 55.995 147.415 ;
        RECT 56.165 147.075 57.470 147.245 ;
        RECT 58.555 147.165 58.875 148.095 ;
        RECT 56.165 146.625 56.410 147.075 ;
        RECT 56.580 146.705 57.130 146.905 ;
        RECT 57.300 146.875 57.470 147.075 ;
        RECT 58.245 146.995 58.875 147.165 ;
        RECT 59.515 147.655 59.845 148.085 ;
        RECT 60.025 147.825 60.220 148.265 ;
        RECT 60.390 147.655 60.720 148.085 ;
        RECT 59.515 147.485 60.720 147.655 ;
        RECT 59.515 147.155 60.410 147.485 ;
        RECT 60.890 147.315 61.165 148.085 ;
        RECT 60.580 147.125 61.165 147.315 ;
        RECT 61.345 147.155 61.605 148.095 ;
        RECT 61.775 147.865 62.105 148.265 ;
        RECT 63.250 148.000 63.505 148.095 ;
        RECT 62.365 147.830 63.505 148.000 ;
        RECT 63.675 147.885 64.005 148.055 ;
        RECT 62.365 147.605 62.535 147.830 ;
        RECT 61.775 147.435 62.535 147.605 ;
        RECT 63.250 147.695 63.505 147.830 ;
        RECT 57.300 146.705 57.675 146.875 ;
        RECT 57.845 146.455 58.075 146.955 ;
        RECT 55.825 146.285 58.075 146.455 ;
        RECT 55.875 145.715 56.205 146.105 ;
        RECT 56.375 145.965 56.545 146.285 ;
        RECT 58.245 146.115 58.415 146.995 ;
        RECT 59.520 146.625 59.815 146.955 ;
        RECT 59.995 146.625 60.410 146.955 ;
        RECT 56.715 145.715 57.045 146.105 ;
        RECT 57.460 145.945 58.415 146.115 ;
        RECT 58.585 145.715 58.875 146.550 ;
        RECT 59.515 145.715 59.815 146.445 ;
        RECT 59.995 146.005 60.225 146.625 ;
        RECT 60.580 146.455 60.755 147.125 ;
        RECT 60.425 146.275 60.755 146.455 ;
        RECT 60.925 146.305 61.165 146.955 ;
        RECT 61.345 146.440 61.520 147.155 ;
        RECT 61.775 146.955 61.945 147.435 ;
        RECT 62.800 147.345 62.970 147.535 ;
        RECT 63.250 147.525 63.660 147.695 ;
        RECT 61.690 146.625 61.945 146.955 ;
        RECT 62.170 146.625 62.500 147.245 ;
        RECT 62.800 147.175 63.320 147.345 ;
        RECT 62.670 146.625 62.960 147.005 ;
        RECT 63.150 146.455 63.320 147.175 ;
        RECT 60.425 145.895 60.650 146.275 ;
        RECT 60.820 145.715 61.150 146.105 ;
        RECT 61.345 145.885 61.605 146.440 ;
        RECT 62.440 146.285 63.320 146.455 ;
        RECT 63.490 146.500 63.660 147.525 ;
        RECT 63.835 147.635 64.005 147.885 ;
        RECT 64.175 147.805 64.425 148.265 ;
        RECT 64.595 147.635 64.775 148.095 ;
        RECT 63.835 147.465 64.775 147.635 ;
        RECT 63.860 146.985 64.340 147.285 ;
        RECT 63.490 146.330 63.840 146.500 ;
        RECT 64.080 146.395 64.340 146.985 ;
        RECT 64.540 146.395 64.800 147.285 ;
        RECT 65.035 147.205 65.365 148.055 ;
        RECT 65.035 146.440 65.225 147.205 ;
        RECT 65.535 147.125 65.785 148.265 ;
        RECT 65.975 147.625 66.225 148.045 ;
        RECT 66.455 147.795 66.785 148.265 ;
        RECT 67.015 147.625 67.265 148.045 ;
        RECT 65.975 147.455 67.265 147.625 ;
        RECT 67.445 147.625 67.775 148.055 ;
        RECT 67.445 147.455 67.900 147.625 ;
        RECT 65.965 146.955 66.180 147.285 ;
        RECT 65.395 146.625 65.705 146.955 ;
        RECT 65.875 146.625 66.180 146.955 ;
        RECT 66.355 146.625 66.640 147.285 ;
        RECT 66.835 146.625 67.100 147.285 ;
        RECT 67.315 146.625 67.560 147.285 ;
        RECT 65.535 146.455 65.705 146.625 ;
        RECT 67.730 146.455 67.900 147.455 ;
        RECT 61.775 145.715 62.205 146.160 ;
        RECT 62.440 145.885 62.610 146.285 ;
        RECT 62.780 145.715 63.500 146.115 ;
        RECT 63.670 145.885 63.840 146.330 ;
        RECT 64.415 145.715 64.815 146.225 ;
        RECT 65.035 145.930 65.365 146.440 ;
        RECT 65.535 146.285 67.900 146.455 ;
        RECT 68.710 147.315 68.975 148.085 ;
        RECT 69.145 147.545 69.475 148.265 ;
        RECT 69.665 147.725 69.925 148.085 ;
        RECT 70.095 147.895 70.425 148.265 ;
        RECT 70.595 147.725 70.855 148.085 ;
        RECT 69.665 147.495 70.855 147.725 ;
        RECT 71.425 147.315 71.715 148.085 ;
        RECT 65.535 145.715 65.865 146.115 ;
        RECT 66.915 145.945 67.245 146.285 ;
        RECT 67.415 145.715 67.745 146.115 ;
        RECT 68.710 145.895 69.045 147.315 ;
        RECT 69.220 147.135 71.715 147.315 ;
        RECT 71.925 147.175 75.435 148.265 ;
        RECT 69.220 146.445 69.445 147.135 ;
        RECT 69.645 146.625 69.925 146.955 ;
        RECT 70.105 146.625 70.680 146.955 ;
        RECT 70.860 146.625 71.295 146.955 ;
        RECT 71.475 146.625 71.745 146.955 ;
        RECT 71.925 146.485 73.575 147.005 ;
        RECT 73.745 146.655 75.435 147.175 ;
        RECT 75.605 147.100 75.895 148.265 ;
        RECT 76.985 147.295 77.295 148.095 ;
        RECT 77.465 147.465 77.775 148.265 ;
        RECT 77.945 147.635 78.205 148.095 ;
        RECT 78.375 147.805 78.630 148.265 ;
        RECT 78.805 147.635 79.065 148.095 ;
        RECT 77.945 147.465 79.065 147.635 ;
        RECT 76.985 147.125 78.015 147.295 ;
        RECT 69.220 146.255 71.705 146.445 ;
        RECT 69.225 145.715 69.970 146.085 ;
        RECT 70.535 145.895 70.790 146.255 ;
        RECT 70.970 145.715 71.300 146.085 ;
        RECT 71.480 145.895 71.705 146.255 ;
        RECT 71.925 145.715 75.435 146.485 ;
        RECT 75.605 145.715 75.895 146.440 ;
        RECT 76.985 146.215 77.155 147.125 ;
        RECT 77.325 146.385 77.675 146.955 ;
        RECT 77.845 146.875 78.015 147.125 ;
        RECT 78.805 147.215 79.065 147.465 ;
        RECT 79.235 147.395 79.520 148.265 ;
        RECT 78.805 147.045 79.560 147.215 ;
        RECT 77.845 146.705 78.985 146.875 ;
        RECT 79.155 146.535 79.560 147.045 ;
        RECT 77.910 146.365 79.560 146.535 ;
        RECT 79.745 147.125 80.085 148.095 ;
        RECT 80.255 147.125 80.425 148.265 ;
        RECT 80.695 147.465 80.945 148.265 ;
        RECT 81.590 147.295 81.920 148.095 ;
        RECT 82.220 147.465 82.550 148.265 ;
        RECT 82.720 147.295 83.050 148.095 ;
        RECT 80.615 147.125 83.050 147.295 ;
        RECT 83.425 147.175 85.095 148.265 ;
        RECT 85.725 147.755 86.025 148.265 ;
        RECT 86.195 147.585 86.525 148.095 ;
        RECT 86.695 147.755 87.325 148.265 ;
        RECT 87.905 147.755 88.285 147.925 ;
        RECT 88.455 147.755 88.755 148.265 ;
        RECT 88.945 147.830 94.290 148.265 ;
        RECT 88.115 147.585 88.285 147.755 ;
        RECT 79.745 147.075 79.975 147.125 ;
        RECT 79.745 146.515 79.920 147.075 ;
        RECT 80.615 146.875 80.785 147.125 ;
        RECT 80.090 146.705 80.785 146.875 ;
        RECT 80.960 146.705 81.380 146.905 ;
        RECT 81.550 146.705 81.880 146.905 ;
        RECT 82.050 146.705 82.380 146.905 ;
        RECT 76.985 145.885 77.285 146.215 ;
        RECT 77.455 145.715 77.730 146.195 ;
        RECT 77.910 145.975 78.205 146.365 ;
        RECT 78.375 145.715 78.630 146.195 ;
        RECT 78.805 145.975 79.065 146.365 ;
        RECT 79.235 145.715 79.515 146.195 ;
        RECT 79.745 145.885 80.085 146.515 ;
        RECT 80.255 145.715 80.505 146.515 ;
        RECT 80.695 146.365 81.920 146.535 ;
        RECT 80.695 145.885 81.025 146.365 ;
        RECT 81.195 145.715 81.420 146.175 ;
        RECT 81.590 145.885 81.920 146.365 ;
        RECT 82.550 146.495 82.720 147.125 ;
        RECT 82.905 146.705 83.255 146.955 ;
        RECT 82.550 145.885 83.050 146.495 ;
        RECT 83.425 146.485 84.175 147.005 ;
        RECT 84.345 146.655 85.095 147.175 ;
        RECT 85.725 147.415 87.945 147.585 ;
        RECT 83.425 145.715 85.095 146.485 ;
        RECT 85.725 146.455 85.895 147.415 ;
        RECT 86.065 147.075 87.605 147.245 ;
        RECT 86.065 146.625 86.310 147.075 ;
        RECT 86.570 146.705 87.265 146.905 ;
        RECT 87.435 146.875 87.605 147.075 ;
        RECT 87.775 147.215 87.945 147.415 ;
        RECT 88.115 147.385 88.775 147.585 ;
        RECT 87.775 147.045 88.435 147.215 ;
        RECT 87.435 146.705 88.035 146.875 ;
        RECT 88.265 146.625 88.435 147.045 ;
        RECT 85.725 145.910 86.190 146.455 ;
        RECT 86.695 145.715 86.865 146.535 ;
        RECT 87.035 146.455 87.945 146.535 ;
        RECT 88.605 146.455 88.775 147.385 ;
        RECT 87.035 146.365 88.285 146.455 ;
        RECT 87.035 145.885 87.365 146.365 ;
        RECT 87.775 146.285 88.285 146.365 ;
        RECT 87.535 145.715 87.885 146.105 ;
        RECT 88.055 145.885 88.285 146.285 ;
        RECT 88.455 145.975 88.775 146.455 ;
        RECT 90.530 146.260 90.870 147.090 ;
        RECT 92.350 146.580 92.700 147.830 ;
        RECT 94.465 147.175 97.975 148.265 ;
        RECT 98.145 147.175 99.355 148.265 ;
        RECT 94.465 146.485 96.115 147.005 ;
        RECT 96.285 146.655 97.975 147.175 ;
        RECT 88.945 145.715 94.290 146.260 ;
        RECT 94.465 145.715 97.975 146.485 ;
        RECT 98.145 146.465 98.665 147.005 ;
        RECT 98.835 146.635 99.355 147.175 ;
        RECT 99.565 147.125 99.795 148.265 ;
        RECT 99.965 147.115 100.295 148.095 ;
        RECT 100.465 147.125 100.675 148.265 ;
        RECT 99.545 146.705 99.875 146.955 ;
        RECT 98.145 145.715 99.355 146.465 ;
        RECT 99.565 145.715 99.795 146.535 ;
        RECT 100.045 146.515 100.295 147.115 ;
        RECT 101.365 147.100 101.655 148.265 ;
        RECT 101.825 147.595 102.140 148.095 ;
        RECT 102.310 147.765 102.560 148.265 ;
        RECT 102.730 147.595 102.980 148.095 ;
        RECT 103.150 147.765 103.400 148.265 ;
        RECT 103.570 147.595 103.820 148.095 ;
        RECT 104.130 147.755 104.380 148.095 ;
        RECT 104.550 147.765 104.800 148.265 ;
        RECT 104.970 147.925 106.095 148.095 ;
        RECT 104.970 147.755 105.295 147.925 ;
        RECT 105.845 147.765 106.095 147.925 ;
        RECT 106.365 147.765 106.615 148.265 ;
        RECT 101.825 147.585 103.820 147.595 ;
        RECT 105.465 147.595 105.675 147.755 ;
        RECT 106.785 147.595 107.035 147.755 ;
        RECT 101.825 147.415 105.220 147.585 ;
        RECT 105.465 147.425 107.035 147.595 ;
        RECT 107.205 147.425 107.635 148.265 ;
        RECT 99.965 145.885 100.295 146.515 ;
        RECT 100.465 145.715 100.675 146.535 ;
        RECT 101.825 146.525 102.055 147.415 ;
        RECT 105.050 147.255 105.220 147.415 ;
        RECT 106.785 147.255 107.035 147.425 ;
        RECT 102.530 147.075 104.840 147.245 ;
        RECT 105.050 147.085 106.545 147.255 ;
        RECT 102.530 146.915 102.700 147.075 ;
        RECT 102.225 146.705 102.700 146.915 ;
        RECT 104.670 146.915 104.840 147.075 ;
        RECT 102.995 146.705 104.445 146.905 ;
        RECT 104.670 146.705 105.695 146.915 ;
        RECT 106.375 146.875 106.545 147.085 ;
        RECT 106.785 147.045 107.635 147.255 ;
        RECT 107.805 147.125 108.065 148.265 ;
        RECT 108.235 147.115 108.565 148.095 ;
        RECT 108.735 147.125 109.015 148.265 ;
        RECT 109.645 147.755 109.945 148.265 ;
        RECT 110.115 147.585 110.445 148.095 ;
        RECT 110.615 147.755 111.245 148.265 ;
        RECT 111.825 147.755 112.205 147.925 ;
        RECT 112.375 147.755 112.675 148.265 ;
        RECT 113.330 147.875 113.665 148.095 ;
        RECT 114.670 147.885 115.025 148.265 ;
        RECT 112.035 147.585 112.205 147.755 ;
        RECT 109.645 147.415 111.865 147.585 ;
        RECT 106.375 146.705 107.035 146.875 ;
        RECT 101.365 145.715 101.655 146.440 ;
        RECT 101.825 146.275 102.600 146.525 ;
        RECT 102.770 146.355 103.860 146.535 ;
        RECT 102.770 146.105 103.020 146.355 ;
        RECT 101.845 145.885 103.020 146.105 ;
        RECT 103.190 145.715 103.360 146.185 ;
        RECT 103.530 145.885 103.860 146.355 ;
        RECT 104.170 145.715 104.340 146.535 ;
        RECT 104.510 146.355 107.075 146.535 ;
        RECT 104.510 145.885 104.840 146.355 ;
        RECT 105.010 145.715 105.180 146.185 ;
        RECT 105.350 145.885 105.715 146.355 ;
        RECT 106.745 146.275 107.075 146.355 ;
        RECT 105.885 145.715 106.055 146.185 ;
        RECT 107.245 146.105 107.635 147.045 ;
        RECT 107.825 146.705 108.160 146.955 ;
        RECT 108.330 146.515 108.500 147.115 ;
        RECT 108.670 146.685 109.005 146.955 ;
        RECT 106.325 145.935 107.635 146.105 ;
        RECT 107.805 145.885 108.500 146.515 ;
        RECT 108.705 145.715 109.015 146.515 ;
        RECT 109.645 146.455 109.815 147.415 ;
        RECT 109.985 147.075 111.525 147.245 ;
        RECT 109.985 146.625 110.230 147.075 ;
        RECT 110.490 146.705 111.185 146.905 ;
        RECT 111.355 146.875 111.525 147.075 ;
        RECT 111.695 147.215 111.865 147.415 ;
        RECT 112.035 147.385 112.695 147.585 ;
        RECT 111.695 147.045 112.355 147.215 ;
        RECT 111.355 146.705 111.955 146.875 ;
        RECT 112.185 146.625 112.355 147.045 ;
        RECT 109.645 145.910 110.110 146.455 ;
        RECT 110.615 145.715 110.785 146.535 ;
        RECT 110.955 146.455 111.865 146.535 ;
        RECT 112.525 146.455 112.695 147.385 ;
        RECT 113.330 147.255 113.585 147.875 ;
        RECT 113.835 147.715 114.065 147.755 ;
        RECT 115.195 147.715 115.445 148.095 ;
        RECT 113.835 147.515 115.445 147.715 ;
        RECT 113.835 147.425 114.020 147.515 ;
        RECT 114.610 147.505 115.445 147.515 ;
        RECT 115.695 147.485 115.945 148.265 ;
        RECT 116.115 147.415 116.375 148.095 ;
        RECT 114.175 147.315 114.505 147.345 ;
        RECT 114.175 147.255 115.975 147.315 ;
        RECT 113.330 147.145 116.035 147.255 ;
        RECT 113.330 147.085 114.505 147.145 ;
        RECT 115.835 147.110 116.035 147.145 ;
        RECT 113.325 146.705 113.815 146.905 ;
        RECT 114.005 146.705 114.480 146.915 ;
        RECT 110.955 146.365 112.205 146.455 ;
        RECT 110.955 145.885 111.285 146.365 ;
        RECT 111.695 146.285 112.205 146.365 ;
        RECT 111.455 145.715 111.805 146.105 ;
        RECT 111.975 145.885 112.205 146.285 ;
        RECT 112.375 145.975 112.695 146.455 ;
        RECT 113.330 145.715 113.785 146.480 ;
        RECT 114.260 146.305 114.480 146.705 ;
        RECT 114.725 146.705 115.055 146.915 ;
        RECT 114.725 146.305 114.935 146.705 ;
        RECT 115.225 146.670 115.635 146.975 ;
        RECT 115.865 146.535 116.035 147.110 ;
        RECT 115.765 146.415 116.035 146.535 ;
        RECT 115.190 146.370 116.035 146.415 ;
        RECT 115.190 146.245 115.945 146.370 ;
        RECT 115.190 146.095 115.360 146.245 ;
        RECT 116.205 146.215 116.375 147.415 ;
        RECT 114.060 145.885 115.360 146.095 ;
        RECT 115.615 145.715 115.945 146.075 ;
        RECT 116.115 145.885 116.375 146.215 ;
        RECT 116.545 147.545 117.005 148.095 ;
        RECT 117.195 147.545 117.525 148.265 ;
        RECT 116.545 146.175 116.795 147.545 ;
        RECT 117.725 147.375 118.025 147.925 ;
        RECT 118.195 147.595 118.475 148.265 ;
        RECT 118.845 147.830 124.190 148.265 ;
        RECT 117.085 147.205 118.025 147.375 ;
        RECT 117.085 146.955 117.255 147.205 ;
        RECT 118.395 146.955 118.660 147.315 ;
        RECT 116.965 146.625 117.255 146.955 ;
        RECT 117.425 146.705 117.765 146.955 ;
        RECT 117.985 146.705 118.660 146.955 ;
        RECT 117.085 146.535 117.255 146.625 ;
        RECT 117.085 146.345 118.475 146.535 ;
        RECT 116.545 145.885 117.105 146.175 ;
        RECT 117.275 145.715 117.525 146.175 ;
        RECT 118.145 145.985 118.475 146.345 ;
        RECT 120.430 146.260 120.770 147.090 ;
        RECT 122.250 146.580 122.600 147.830 ;
        RECT 124.365 147.175 126.955 148.265 ;
        RECT 124.365 146.485 125.575 147.005 ;
        RECT 125.745 146.655 126.955 147.175 ;
        RECT 127.125 147.100 127.415 148.265 ;
        RECT 127.585 147.830 132.930 148.265 ;
        RECT 133.105 147.830 138.450 148.265 ;
        RECT 138.625 147.830 143.970 148.265 ;
        RECT 118.845 145.715 124.190 146.260 ;
        RECT 124.365 145.715 126.955 146.485 ;
        RECT 127.125 145.715 127.415 146.440 ;
        RECT 129.170 146.260 129.510 147.090 ;
        RECT 130.990 146.580 131.340 147.830 ;
        RECT 134.690 146.260 135.030 147.090 ;
        RECT 136.510 146.580 136.860 147.830 ;
        RECT 140.210 146.260 140.550 147.090 ;
        RECT 142.030 146.580 142.380 147.830 ;
        RECT 144.145 147.175 147.655 148.265 ;
        RECT 147.825 147.175 149.035 148.265 ;
        RECT 144.145 146.485 145.795 147.005 ;
        RECT 145.965 146.655 147.655 147.175 ;
        RECT 127.585 145.715 132.930 146.260 ;
        RECT 133.105 145.715 138.450 146.260 ;
        RECT 138.625 145.715 143.970 146.260 ;
        RECT 144.145 145.715 147.655 146.485 ;
        RECT 147.825 146.465 148.345 147.005 ;
        RECT 148.515 146.635 149.035 147.175 ;
        RECT 149.205 147.175 150.415 148.265 ;
        RECT 149.205 146.635 149.725 147.175 ;
        RECT 149.895 146.465 150.415 147.005 ;
        RECT 147.825 145.715 149.035 146.465 ;
        RECT 149.205 145.715 150.415 146.465 ;
        RECT 11.120 145.545 150.500 145.715 ;
        RECT 11.205 144.795 12.415 145.545 ;
        RECT 12.585 145.000 17.930 145.545 ;
        RECT 18.105 145.000 23.450 145.545 ;
        RECT 24.110 145.155 24.440 145.545 ;
        RECT 11.205 144.255 11.725 144.795 ;
        RECT 11.895 144.085 12.415 144.625 ;
        RECT 14.170 144.170 14.510 145.000 ;
        RECT 11.205 142.995 12.415 144.085 ;
        RECT 15.990 143.430 16.340 144.680 ;
        RECT 19.690 144.170 20.030 145.000 ;
        RECT 24.610 144.985 24.835 145.365 ;
        RECT 21.510 143.430 21.860 144.680 ;
        RECT 24.095 144.305 24.335 144.955 ;
        RECT 24.505 144.805 24.835 144.985 ;
        RECT 24.505 144.135 24.680 144.805 ;
        RECT 25.035 144.635 25.265 145.255 ;
        RECT 25.445 144.815 25.745 145.545 ;
        RECT 26.435 145.155 26.765 145.545 ;
        RECT 26.935 144.975 27.105 145.295 ;
        RECT 27.275 145.155 27.605 145.545 ;
        RECT 28.020 145.145 28.975 145.315 ;
        RECT 26.385 144.805 28.635 144.975 ;
        RECT 24.850 144.305 25.265 144.635 ;
        RECT 25.445 144.305 25.740 144.635 ;
        RECT 24.095 143.945 24.680 144.135 ;
        RECT 12.585 142.995 17.930 143.430 ;
        RECT 18.105 142.995 23.450 143.430 ;
        RECT 24.095 143.175 24.370 143.945 ;
        RECT 24.850 143.775 25.745 144.105 ;
        RECT 24.540 143.605 25.745 143.775 ;
        RECT 24.540 143.175 24.870 143.605 ;
        RECT 25.040 142.995 25.235 143.435 ;
        RECT 25.415 143.175 25.745 143.605 ;
        RECT 26.385 143.845 26.555 144.805 ;
        RECT 26.725 144.185 26.970 144.635 ;
        RECT 27.140 144.355 27.690 144.555 ;
        RECT 27.860 144.385 28.235 144.555 ;
        RECT 27.860 144.185 28.030 144.385 ;
        RECT 28.405 144.305 28.635 144.805 ;
        RECT 26.725 144.015 28.030 144.185 ;
        RECT 28.805 144.265 28.975 145.145 ;
        RECT 29.145 144.710 29.435 145.545 ;
        RECT 29.605 145.000 34.950 145.545 ;
        RECT 28.805 144.095 29.435 144.265 ;
        RECT 31.190 144.170 31.530 145.000 ;
        RECT 35.125 144.775 36.795 145.545 ;
        RECT 36.965 144.820 37.255 145.545 ;
        RECT 37.625 144.915 37.955 145.275 ;
        RECT 38.575 145.085 38.825 145.545 ;
        RECT 38.995 145.085 39.555 145.375 ;
        RECT 26.385 143.165 26.765 143.845 ;
        RECT 27.355 142.995 27.525 143.845 ;
        RECT 27.695 143.675 28.935 143.845 ;
        RECT 27.695 143.165 28.025 143.675 ;
        RECT 28.195 142.995 28.365 143.505 ;
        RECT 28.535 143.165 28.935 143.675 ;
        RECT 29.115 143.165 29.435 144.095 ;
        RECT 33.010 143.430 33.360 144.680 ;
        RECT 35.125 144.255 35.875 144.775 ;
        RECT 37.625 144.725 39.015 144.915 ;
        RECT 38.845 144.635 39.015 144.725 ;
        RECT 36.045 144.085 36.795 144.605 ;
        RECT 37.440 144.305 38.115 144.555 ;
        RECT 38.335 144.305 38.675 144.555 ;
        RECT 38.845 144.305 39.135 144.635 ;
        RECT 29.605 142.995 34.950 143.430 ;
        RECT 35.125 142.995 36.795 144.085 ;
        RECT 36.965 142.995 37.255 144.160 ;
        RECT 37.440 143.945 37.705 144.305 ;
        RECT 38.845 144.055 39.015 144.305 ;
        RECT 38.075 143.885 39.015 144.055 ;
        RECT 37.625 142.995 37.905 143.665 ;
        RECT 38.075 143.335 38.375 143.885 ;
        RECT 39.305 143.715 39.555 145.085 ;
        RECT 38.575 142.995 38.905 143.715 ;
        RECT 39.095 143.165 39.555 143.715 ;
        RECT 39.725 144.870 39.985 145.375 ;
        RECT 40.165 145.165 40.495 145.545 ;
        RECT 40.675 144.995 40.845 145.375 ;
        RECT 41.105 145.000 46.450 145.545 ;
        RECT 39.725 144.070 39.895 144.870 ;
        RECT 40.180 144.825 40.845 144.995 ;
        RECT 40.180 144.570 40.350 144.825 ;
        RECT 40.065 144.240 40.350 144.570 ;
        RECT 40.585 144.275 40.915 144.645 ;
        RECT 40.180 144.095 40.350 144.240 ;
        RECT 42.690 144.170 43.030 145.000 ;
        RECT 46.625 144.775 50.135 145.545 ;
        RECT 50.775 144.895 51.105 145.360 ;
        RECT 51.275 145.075 51.445 145.545 ;
        RECT 51.620 145.145 51.950 145.375 ;
        RECT 51.700 144.895 51.870 145.145 ;
        RECT 52.155 144.985 52.325 145.375 ;
        RECT 39.725 143.165 39.995 144.070 ;
        RECT 40.180 143.925 40.845 144.095 ;
        RECT 40.165 142.995 40.495 143.755 ;
        RECT 40.675 143.165 40.845 143.925 ;
        RECT 44.510 143.430 44.860 144.680 ;
        RECT 46.625 144.255 48.275 144.775 ;
        RECT 50.775 144.725 51.870 144.895 ;
        RECT 52.085 144.805 52.325 144.985 ;
        RECT 52.670 144.975 52.860 145.135 ;
        RECT 52.550 144.805 52.860 144.975 ;
        RECT 53.080 144.805 53.355 145.545 ;
        RECT 53.525 145.000 58.870 145.545 ;
        RECT 48.445 144.085 50.135 144.605 ;
        RECT 50.765 144.345 51.245 144.555 ;
        RECT 51.415 144.345 51.915 144.555 ;
        RECT 52.085 144.175 52.255 144.805 ;
        RECT 52.550 144.635 52.720 144.805 ;
        RECT 41.105 142.995 46.450 143.430 ;
        RECT 46.625 142.995 50.135 144.085 ;
        RECT 50.795 142.995 51.170 144.095 ;
        RECT 51.645 144.005 52.255 144.175 ;
        RECT 52.425 144.095 52.720 144.635 ;
        RECT 52.905 144.285 53.355 144.635 ;
        RECT 51.645 143.165 51.970 144.005 ;
        RECT 52.425 143.925 52.915 144.095 ;
        RECT 52.140 142.995 52.470 143.755 ;
        RECT 52.640 143.420 52.915 143.925 ;
        RECT 53.085 143.185 53.355 144.285 ;
        RECT 55.110 144.170 55.450 145.000 ;
        RECT 59.045 144.795 60.255 145.545 ;
        RECT 60.625 144.915 60.955 145.275 ;
        RECT 61.575 145.085 61.825 145.545 ;
        RECT 61.995 145.085 62.555 145.375 ;
        RECT 56.930 143.430 57.280 144.680 ;
        RECT 59.045 144.255 59.565 144.795 ;
        RECT 60.625 144.725 62.015 144.915 ;
        RECT 61.845 144.635 62.015 144.725 ;
        RECT 59.735 144.085 60.255 144.625 ;
        RECT 53.525 142.995 58.870 143.430 ;
        RECT 59.045 142.995 60.255 144.085 ;
        RECT 60.440 144.305 61.115 144.555 ;
        RECT 61.335 144.305 61.675 144.555 ;
        RECT 61.845 144.305 62.135 144.635 ;
        RECT 60.440 143.945 60.705 144.305 ;
        RECT 61.845 144.055 62.015 144.305 ;
        RECT 61.075 143.885 62.015 144.055 ;
        RECT 60.625 142.995 60.905 143.665 ;
        RECT 61.075 143.335 61.375 143.885 ;
        RECT 62.305 143.715 62.555 145.085 ;
        RECT 62.725 144.820 63.015 145.545 ;
        RECT 63.735 144.995 63.905 145.285 ;
        RECT 64.075 145.165 64.405 145.545 ;
        RECT 63.735 144.825 64.400 144.995 ;
        RECT 61.575 142.995 61.905 143.715 ;
        RECT 62.095 143.165 62.555 143.715 ;
        RECT 62.725 142.995 63.015 144.160 ;
        RECT 63.650 144.005 64.000 144.655 ;
        RECT 64.170 143.835 64.400 144.825 ;
        RECT 63.735 143.665 64.400 143.835 ;
        RECT 63.735 143.165 63.905 143.665 ;
        RECT 64.075 142.995 64.405 143.495 ;
        RECT 64.575 143.165 64.760 145.285 ;
        RECT 65.015 145.085 65.265 145.545 ;
        RECT 65.435 145.095 65.770 145.265 ;
        RECT 65.965 145.095 66.640 145.265 ;
        RECT 65.435 144.955 65.605 145.095 ;
        RECT 64.930 143.965 65.210 144.915 ;
        RECT 65.380 144.825 65.605 144.955 ;
        RECT 65.380 143.720 65.550 144.825 ;
        RECT 65.775 144.675 66.300 144.895 ;
        RECT 65.720 143.910 65.960 144.505 ;
        RECT 66.130 143.975 66.300 144.675 ;
        RECT 66.470 144.315 66.640 145.095 ;
        RECT 66.960 145.045 67.330 145.545 ;
        RECT 67.510 145.095 67.915 145.265 ;
        RECT 68.085 145.095 68.870 145.265 ;
        RECT 67.510 144.865 67.680 145.095 ;
        RECT 66.850 144.565 67.680 144.865 ;
        RECT 68.065 144.595 68.530 144.925 ;
        RECT 66.850 144.535 67.050 144.565 ;
        RECT 67.170 144.315 67.340 144.385 ;
        RECT 66.470 144.145 67.340 144.315 ;
        RECT 66.830 144.055 67.340 144.145 ;
        RECT 65.380 143.590 65.685 143.720 ;
        RECT 66.130 143.610 66.660 143.975 ;
        RECT 65.000 142.995 65.265 143.455 ;
        RECT 65.435 143.165 65.685 143.590 ;
        RECT 66.830 143.440 67.000 144.055 ;
        RECT 65.895 143.270 67.000 143.440 ;
        RECT 67.170 142.995 67.340 143.795 ;
        RECT 67.510 143.495 67.680 144.565 ;
        RECT 67.850 143.665 68.040 144.385 ;
        RECT 68.210 143.635 68.530 144.595 ;
        RECT 68.700 144.635 68.870 145.095 ;
        RECT 69.145 145.015 69.355 145.545 ;
        RECT 69.615 144.805 69.945 145.330 ;
        RECT 70.115 144.935 70.285 145.545 ;
        RECT 70.455 144.890 70.785 145.325 ;
        RECT 71.095 144.995 71.265 145.285 ;
        RECT 71.435 145.165 71.765 145.545 ;
        RECT 70.455 144.805 70.835 144.890 ;
        RECT 71.095 144.825 71.760 144.995 ;
        RECT 69.745 144.635 69.945 144.805 ;
        RECT 70.610 144.765 70.835 144.805 ;
        RECT 68.700 144.305 69.575 144.635 ;
        RECT 69.745 144.305 70.495 144.635 ;
        RECT 67.510 143.165 67.760 143.495 ;
        RECT 68.700 143.465 68.870 144.305 ;
        RECT 69.745 144.100 69.935 144.305 ;
        RECT 70.665 144.185 70.835 144.765 ;
        RECT 70.620 144.135 70.835 144.185 ;
        RECT 69.040 143.725 69.935 144.100 ;
        RECT 70.445 144.055 70.835 144.135 ;
        RECT 67.985 143.295 68.870 143.465 ;
        RECT 69.050 142.995 69.365 143.495 ;
        RECT 69.595 143.165 69.935 143.725 ;
        RECT 70.105 142.995 70.275 144.005 ;
        RECT 70.445 143.210 70.775 144.055 ;
        RECT 71.010 144.005 71.360 144.655 ;
        RECT 71.530 143.835 71.760 144.825 ;
        RECT 71.095 143.665 71.760 143.835 ;
        RECT 71.095 143.165 71.265 143.665 ;
        RECT 71.435 142.995 71.765 143.495 ;
        RECT 71.935 143.165 72.120 145.285 ;
        RECT 72.375 145.085 72.625 145.545 ;
        RECT 72.795 145.095 73.130 145.265 ;
        RECT 73.325 145.095 74.000 145.265 ;
        RECT 72.795 144.955 72.965 145.095 ;
        RECT 72.290 143.965 72.570 144.915 ;
        RECT 72.740 144.825 72.965 144.955 ;
        RECT 72.740 143.720 72.910 144.825 ;
        RECT 73.135 144.675 73.660 144.895 ;
        RECT 73.080 143.910 73.320 144.505 ;
        RECT 73.490 143.975 73.660 144.675 ;
        RECT 73.830 144.315 74.000 145.095 ;
        RECT 74.320 145.045 74.690 145.545 ;
        RECT 74.870 145.095 75.275 145.265 ;
        RECT 75.445 145.095 76.230 145.265 ;
        RECT 74.870 144.865 75.040 145.095 ;
        RECT 74.210 144.565 75.040 144.865 ;
        RECT 75.425 144.595 75.890 144.925 ;
        RECT 74.210 144.535 74.410 144.565 ;
        RECT 74.530 144.315 74.700 144.385 ;
        RECT 73.830 144.145 74.700 144.315 ;
        RECT 74.190 144.055 74.700 144.145 ;
        RECT 72.740 143.590 73.045 143.720 ;
        RECT 73.490 143.610 74.020 143.975 ;
        RECT 72.360 142.995 72.625 143.455 ;
        RECT 72.795 143.165 73.045 143.590 ;
        RECT 74.190 143.440 74.360 144.055 ;
        RECT 73.255 143.270 74.360 143.440 ;
        RECT 74.530 142.995 74.700 143.795 ;
        RECT 74.870 143.495 75.040 144.565 ;
        RECT 75.210 143.665 75.400 144.385 ;
        RECT 75.570 143.635 75.890 144.595 ;
        RECT 76.060 144.635 76.230 145.095 ;
        RECT 76.505 145.015 76.715 145.545 ;
        RECT 76.975 144.805 77.305 145.330 ;
        RECT 77.475 144.935 77.645 145.545 ;
        RECT 77.815 144.890 78.145 145.325 ;
        RECT 78.435 145.145 78.765 145.545 ;
        RECT 78.935 144.975 79.105 145.245 ;
        RECT 79.275 145.145 79.605 145.545 ;
        RECT 79.775 144.975 80.030 145.245 ;
        RECT 77.815 144.805 78.195 144.890 ;
        RECT 77.105 144.635 77.305 144.805 ;
        RECT 77.970 144.765 78.195 144.805 ;
        RECT 76.060 144.305 76.935 144.635 ;
        RECT 77.105 144.305 77.855 144.635 ;
        RECT 74.870 143.165 75.120 143.495 ;
        RECT 76.060 143.465 76.230 144.305 ;
        RECT 77.105 144.100 77.295 144.305 ;
        RECT 78.025 144.185 78.195 144.765 ;
        RECT 77.980 144.135 78.195 144.185 ;
        RECT 76.400 143.725 77.295 144.100 ;
        RECT 77.805 144.055 78.195 144.135 ;
        RECT 75.345 143.295 76.230 143.465 ;
        RECT 76.410 142.995 76.725 143.495 ;
        RECT 76.955 143.165 77.295 143.725 ;
        RECT 77.465 142.995 77.635 144.005 ;
        RECT 77.805 143.210 78.135 144.055 ;
        RECT 78.365 143.965 78.635 144.975 ;
        RECT 78.805 144.805 80.030 144.975 ;
        RECT 78.805 144.135 78.975 144.805 ;
        RECT 80.205 144.775 81.875 145.545 ;
        RECT 82.080 144.805 82.695 145.375 ;
        RECT 82.865 145.035 83.080 145.545 ;
        RECT 83.310 145.035 83.590 145.365 ;
        RECT 83.770 145.035 84.010 145.545 ;
        RECT 79.145 144.305 79.525 144.635 ;
        RECT 79.695 144.305 80.030 144.635 ;
        RECT 78.805 143.965 79.120 144.135 ;
        RECT 78.370 142.995 78.685 143.795 ;
        RECT 78.950 143.350 79.120 143.965 ;
        RECT 79.290 143.625 79.525 144.305 ;
        RECT 80.205 144.255 80.955 144.775 ;
        RECT 79.695 143.350 80.030 144.135 ;
        RECT 81.125 144.085 81.875 144.605 ;
        RECT 78.950 143.180 80.030 143.350 ;
        RECT 80.205 142.995 81.875 144.085 ;
        RECT 82.080 143.785 82.395 144.805 ;
        RECT 82.565 144.135 82.735 144.635 ;
        RECT 82.985 144.305 83.250 144.865 ;
        RECT 83.420 144.135 83.590 145.035 ;
        RECT 83.760 144.305 84.115 144.865 ;
        RECT 84.345 144.775 86.015 145.545 ;
        RECT 86.185 144.895 86.445 145.375 ;
        RECT 86.615 145.005 86.865 145.545 ;
        RECT 84.345 144.255 85.095 144.775 ;
        RECT 82.565 143.965 83.990 144.135 ;
        RECT 85.265 144.085 86.015 144.605 ;
        RECT 82.080 143.165 82.615 143.785 ;
        RECT 82.785 142.995 83.115 143.795 ;
        RECT 83.600 143.790 83.990 143.965 ;
        RECT 84.345 142.995 86.015 144.085 ;
        RECT 86.185 143.865 86.355 144.895 ;
        RECT 87.035 144.865 87.255 145.325 ;
        RECT 87.005 144.840 87.255 144.865 ;
        RECT 86.525 144.245 86.755 144.640 ;
        RECT 86.925 144.415 87.255 144.840 ;
        RECT 87.425 145.165 88.315 145.335 ;
        RECT 87.425 144.440 87.595 145.165 ;
        RECT 87.765 144.610 88.315 144.995 ;
        RECT 88.485 144.820 88.775 145.545 ;
        RECT 88.945 145.085 89.505 145.375 ;
        RECT 89.675 145.085 89.925 145.545 ;
        RECT 87.425 144.370 88.315 144.440 ;
        RECT 87.420 144.345 88.315 144.370 ;
        RECT 87.410 144.330 88.315 144.345 ;
        RECT 87.405 144.315 88.315 144.330 ;
        RECT 87.395 144.310 88.315 144.315 ;
        RECT 87.390 144.300 88.315 144.310 ;
        RECT 87.385 144.290 88.315 144.300 ;
        RECT 87.375 144.285 88.315 144.290 ;
        RECT 87.365 144.275 88.315 144.285 ;
        RECT 87.355 144.270 88.315 144.275 ;
        RECT 87.355 144.265 87.690 144.270 ;
        RECT 87.340 144.260 87.690 144.265 ;
        RECT 87.325 144.250 87.690 144.260 ;
        RECT 87.300 144.245 87.690 144.250 ;
        RECT 86.525 144.240 87.690 144.245 ;
        RECT 86.525 144.205 87.660 144.240 ;
        RECT 86.525 144.180 87.625 144.205 ;
        RECT 86.525 144.150 87.595 144.180 ;
        RECT 86.525 144.120 87.575 144.150 ;
        RECT 86.525 144.090 87.555 144.120 ;
        RECT 86.525 144.080 87.485 144.090 ;
        RECT 86.525 144.070 87.460 144.080 ;
        RECT 86.525 144.055 87.440 144.070 ;
        RECT 86.525 144.040 87.420 144.055 ;
        RECT 86.630 144.030 87.415 144.040 ;
        RECT 86.630 143.995 87.400 144.030 ;
        RECT 86.185 143.165 86.460 143.865 ;
        RECT 86.630 143.745 87.385 143.995 ;
        RECT 87.555 143.675 87.885 143.920 ;
        RECT 88.055 143.820 88.315 144.270 ;
        RECT 87.700 143.650 87.885 143.675 ;
        RECT 87.700 143.550 88.315 143.650 ;
        RECT 86.630 142.995 86.885 143.540 ;
        RECT 87.055 143.165 87.535 143.505 ;
        RECT 87.710 142.995 88.315 143.550 ;
        RECT 88.485 142.995 88.775 144.160 ;
        RECT 88.945 143.715 89.195 145.085 ;
        RECT 90.545 144.915 90.875 145.275 ;
        RECT 89.485 144.725 90.875 144.915 ;
        RECT 92.165 144.805 92.630 145.350 ;
        RECT 89.485 144.635 89.655 144.725 ;
        RECT 89.365 144.305 89.655 144.635 ;
        RECT 89.825 144.305 90.165 144.555 ;
        RECT 90.385 144.305 91.060 144.555 ;
        RECT 89.485 144.055 89.655 144.305 ;
        RECT 89.485 143.885 90.425 144.055 ;
        RECT 90.795 143.945 91.060 144.305 ;
        RECT 88.945 143.165 89.405 143.715 ;
        RECT 89.595 142.995 89.925 143.715 ;
        RECT 90.125 143.335 90.425 143.885 ;
        RECT 92.165 143.845 92.335 144.805 ;
        RECT 93.135 144.725 93.305 145.545 ;
        RECT 93.475 144.895 93.805 145.375 ;
        RECT 93.975 145.155 94.325 145.545 ;
        RECT 94.495 144.975 94.725 145.375 ;
        RECT 94.215 144.895 94.725 144.975 ;
        RECT 93.475 144.805 94.725 144.895 ;
        RECT 94.895 144.805 95.215 145.285 ;
        RECT 95.385 145.000 100.730 145.545 ;
        RECT 93.475 144.725 94.385 144.805 ;
        RECT 92.505 144.185 92.750 144.635 ;
        RECT 93.010 144.355 93.705 144.555 ;
        RECT 93.875 144.385 94.475 144.555 ;
        RECT 93.875 144.185 94.045 144.385 ;
        RECT 94.705 144.215 94.875 144.635 ;
        RECT 92.505 144.015 94.045 144.185 ;
        RECT 94.215 144.045 94.875 144.215 ;
        RECT 94.215 143.845 94.385 144.045 ;
        RECT 95.045 143.875 95.215 144.805 ;
        RECT 96.970 144.170 97.310 145.000 ;
        RECT 100.905 144.775 102.575 145.545 ;
        RECT 102.750 145.040 103.085 145.545 ;
        RECT 103.255 144.975 103.495 145.350 ;
        RECT 103.775 145.215 103.945 145.360 ;
        RECT 103.775 145.020 104.150 145.215 ;
        RECT 104.510 145.050 104.905 145.545 ;
        RECT 92.165 143.675 94.385 143.845 ;
        RECT 94.555 143.675 95.215 143.875 ;
        RECT 90.595 142.995 90.875 143.665 ;
        RECT 92.165 142.995 92.465 143.505 ;
        RECT 92.635 143.165 92.965 143.675 ;
        RECT 94.555 143.505 94.725 143.675 ;
        RECT 93.135 142.995 93.765 143.505 ;
        RECT 94.345 143.335 94.725 143.505 ;
        RECT 94.895 142.995 95.195 143.505 ;
        RECT 98.790 143.430 99.140 144.680 ;
        RECT 100.905 144.255 101.655 144.775 ;
        RECT 101.825 144.085 102.575 144.605 ;
        RECT 95.385 142.995 100.730 143.430 ;
        RECT 100.905 142.995 102.575 144.085 ;
        RECT 102.805 144.015 103.105 144.865 ;
        RECT 103.275 144.825 103.495 144.975 ;
        RECT 103.275 144.495 103.810 144.825 ;
        RECT 103.980 144.685 104.150 145.020 ;
        RECT 105.075 144.855 105.315 145.375 ;
        RECT 105.505 145.000 110.850 145.545 ;
        RECT 103.275 143.845 103.510 144.495 ;
        RECT 103.980 144.325 104.965 144.685 ;
        RECT 102.835 143.615 103.510 143.845 ;
        RECT 103.680 144.305 104.965 144.325 ;
        RECT 103.680 144.155 104.540 144.305 ;
        RECT 102.835 143.185 103.005 143.615 ;
        RECT 103.175 142.995 103.505 143.445 ;
        RECT 103.680 143.210 103.965 144.155 ;
        RECT 105.140 144.050 105.315 144.855 ;
        RECT 107.090 144.170 107.430 145.000 ;
        RECT 111.025 144.775 113.615 145.545 ;
        RECT 114.245 144.820 114.535 145.545 ;
        RECT 115.715 144.995 115.885 145.375 ;
        RECT 116.065 145.165 116.395 145.545 ;
        RECT 115.715 144.825 116.380 144.995 ;
        RECT 116.575 144.870 116.835 145.375 ;
        RECT 117.005 145.000 122.350 145.545 ;
        RECT 122.525 145.000 127.870 145.545 ;
        RECT 128.045 145.000 133.390 145.545 ;
        RECT 133.565 145.000 138.910 145.545 ;
        RECT 104.140 143.675 104.835 143.985 ;
        RECT 104.145 142.995 104.830 143.465 ;
        RECT 105.010 143.265 105.315 144.050 ;
        RECT 108.910 143.430 109.260 144.680 ;
        RECT 111.025 144.255 112.235 144.775 ;
        RECT 112.405 144.085 113.615 144.605 ;
        RECT 115.645 144.275 115.975 144.645 ;
        RECT 116.210 144.570 116.380 144.825 ;
        RECT 116.210 144.240 116.495 144.570 ;
        RECT 105.505 142.995 110.850 143.430 ;
        RECT 111.025 142.995 113.615 144.085 ;
        RECT 114.245 142.995 114.535 144.160 ;
        RECT 116.210 144.095 116.380 144.240 ;
        RECT 115.715 143.925 116.380 144.095 ;
        RECT 116.665 144.070 116.835 144.870 ;
        RECT 118.590 144.170 118.930 145.000 ;
        RECT 115.715 143.165 115.885 143.925 ;
        RECT 116.065 142.995 116.395 143.755 ;
        RECT 116.565 143.165 116.835 144.070 ;
        RECT 120.410 143.430 120.760 144.680 ;
        RECT 124.110 144.170 124.450 145.000 ;
        RECT 125.930 143.430 126.280 144.680 ;
        RECT 129.630 144.170 129.970 145.000 ;
        RECT 131.450 143.430 131.800 144.680 ;
        RECT 135.150 144.170 135.490 145.000 ;
        RECT 140.005 144.820 140.295 145.545 ;
        RECT 140.465 145.000 145.810 145.545 ;
        RECT 136.970 143.430 137.320 144.680 ;
        RECT 142.050 144.170 142.390 145.000 ;
        RECT 145.985 144.775 148.575 145.545 ;
        RECT 149.205 144.795 150.415 145.545 ;
        RECT 117.005 142.995 122.350 143.430 ;
        RECT 122.525 142.995 127.870 143.430 ;
        RECT 128.045 142.995 133.390 143.430 ;
        RECT 133.565 142.995 138.910 143.430 ;
        RECT 140.005 142.995 140.295 144.160 ;
        RECT 143.870 143.430 144.220 144.680 ;
        RECT 145.985 144.255 147.195 144.775 ;
        RECT 147.365 144.085 148.575 144.605 ;
        RECT 140.465 142.995 145.810 143.430 ;
        RECT 145.985 142.995 148.575 144.085 ;
        RECT 149.205 144.085 149.725 144.625 ;
        RECT 149.895 144.255 150.415 144.795 ;
        RECT 149.205 142.995 150.415 144.085 ;
        RECT 11.120 142.825 150.500 142.995 ;
        RECT 11.205 141.735 12.415 142.825 ;
        RECT 12.585 141.735 16.095 142.825 ;
        RECT 16.265 141.735 17.475 142.825 ;
        RECT 11.205 141.025 11.725 141.565 ;
        RECT 11.895 141.195 12.415 141.735 ;
        RECT 12.585 141.045 14.235 141.565 ;
        RECT 14.405 141.215 16.095 141.735 ;
        RECT 11.205 140.275 12.415 141.025 ;
        RECT 12.585 140.275 16.095 141.045 ;
        RECT 16.265 141.025 16.785 141.565 ;
        RECT 16.955 141.195 17.475 141.735 ;
        RECT 17.645 141.750 17.915 142.655 ;
        RECT 18.085 142.065 18.415 142.825 ;
        RECT 18.595 141.895 18.765 142.655 ;
        RECT 16.265 140.275 17.475 141.025 ;
        RECT 17.645 140.950 17.815 141.750 ;
        RECT 18.100 141.725 18.765 141.895 ;
        RECT 19.025 141.735 22.535 142.825 ;
        RECT 22.705 141.735 23.915 142.825 ;
        RECT 18.100 141.580 18.270 141.725 ;
        RECT 17.985 141.250 18.270 141.580 ;
        RECT 18.100 140.995 18.270 141.250 ;
        RECT 18.505 141.175 18.835 141.545 ;
        RECT 19.025 141.045 20.675 141.565 ;
        RECT 20.845 141.215 22.535 141.735 ;
        RECT 17.645 140.445 17.905 140.950 ;
        RECT 18.100 140.825 18.765 140.995 ;
        RECT 18.085 140.275 18.415 140.655 ;
        RECT 18.595 140.445 18.765 140.825 ;
        RECT 19.025 140.275 22.535 141.045 ;
        RECT 22.705 141.025 23.225 141.565 ;
        RECT 23.395 141.195 23.915 141.735 ;
        RECT 24.085 141.660 24.375 142.825 ;
        RECT 24.545 141.735 28.055 142.825 ;
        RECT 24.545 141.045 26.195 141.565 ;
        RECT 26.365 141.215 28.055 141.735 ;
        RECT 28.225 141.685 28.505 142.825 ;
        RECT 28.675 141.675 29.005 142.655 ;
        RECT 29.175 141.685 29.435 142.825 ;
        RECT 29.605 142.390 34.950 142.825 ;
        RECT 35.590 142.435 35.925 142.655 ;
        RECT 36.930 142.445 37.285 142.825 ;
        RECT 28.235 141.245 28.570 141.515 ;
        RECT 28.740 141.075 28.910 141.675 ;
        RECT 29.080 141.265 29.415 141.515 ;
        RECT 22.705 140.275 23.915 141.025 ;
        RECT 24.085 140.275 24.375 141.000 ;
        RECT 24.545 140.275 28.055 141.045 ;
        RECT 28.225 140.275 28.535 141.075 ;
        RECT 28.740 140.445 29.435 141.075 ;
        RECT 31.190 140.820 31.530 141.650 ;
        RECT 33.010 141.140 33.360 142.390 ;
        RECT 35.590 141.815 35.845 142.435 ;
        RECT 36.095 142.275 36.325 142.315 ;
        RECT 37.455 142.275 37.705 142.655 ;
        RECT 36.095 142.075 37.705 142.275 ;
        RECT 36.095 141.985 36.280 142.075 ;
        RECT 36.870 142.065 37.705 142.075 ;
        RECT 37.955 142.045 38.205 142.825 ;
        RECT 38.375 141.975 38.635 142.655 ;
        RECT 36.435 141.875 36.765 141.905 ;
        RECT 36.435 141.815 38.235 141.875 ;
        RECT 35.590 141.705 38.295 141.815 ;
        RECT 35.590 141.645 36.765 141.705 ;
        RECT 38.095 141.670 38.295 141.705 ;
        RECT 35.585 141.265 36.075 141.465 ;
        RECT 36.265 141.265 36.740 141.475 ;
        RECT 29.605 140.275 34.950 140.820 ;
        RECT 35.590 140.275 36.045 141.040 ;
        RECT 36.520 140.865 36.740 141.265 ;
        RECT 36.985 141.265 37.315 141.475 ;
        RECT 36.985 140.865 37.195 141.265 ;
        RECT 37.485 141.230 37.895 141.535 ;
        RECT 38.125 141.095 38.295 141.670 ;
        RECT 38.025 140.975 38.295 141.095 ;
        RECT 37.450 140.930 38.295 140.975 ;
        RECT 37.450 140.805 38.205 140.930 ;
        RECT 37.450 140.655 37.620 140.805 ;
        RECT 38.465 140.775 38.635 141.975 ;
        RECT 38.805 141.735 42.315 142.825 ;
        RECT 42.575 142.205 42.745 142.635 ;
        RECT 42.915 142.375 43.245 142.825 ;
        RECT 42.575 141.975 43.250 142.205 ;
        RECT 36.320 140.445 37.620 140.655 ;
        RECT 37.875 140.275 38.205 140.635 ;
        RECT 38.375 140.445 38.635 140.775 ;
        RECT 38.805 141.045 40.455 141.565 ;
        RECT 40.625 141.215 42.315 141.735 ;
        RECT 38.805 140.275 42.315 141.045 ;
        RECT 42.545 140.955 42.845 141.805 ;
        RECT 43.015 141.325 43.250 141.975 ;
        RECT 43.420 141.665 43.705 142.610 ;
        RECT 43.885 142.355 44.570 142.825 ;
        RECT 43.880 141.835 44.575 142.145 ;
        RECT 44.750 141.770 45.055 142.555 ;
        RECT 43.420 141.515 44.280 141.665 ;
        RECT 43.420 141.495 44.705 141.515 ;
        RECT 43.015 140.995 43.550 141.325 ;
        RECT 43.720 141.135 44.705 141.495 ;
        RECT 43.015 140.845 43.235 140.995 ;
        RECT 42.490 140.275 42.825 140.780 ;
        RECT 42.995 140.470 43.235 140.845 ;
        RECT 43.720 140.800 43.890 141.135 ;
        RECT 44.880 140.965 45.055 141.770 ;
        RECT 43.515 140.605 43.890 140.800 ;
        RECT 43.515 140.460 43.685 140.605 ;
        RECT 44.250 140.275 44.645 140.770 ;
        RECT 44.815 140.445 45.055 140.965 ;
        RECT 45.265 141.770 45.570 142.555 ;
        RECT 45.750 142.355 46.435 142.825 ;
        RECT 45.745 141.835 46.440 142.145 ;
        RECT 45.265 140.965 45.440 141.770 ;
        RECT 46.615 141.665 46.900 142.610 ;
        RECT 47.075 142.375 47.405 142.825 ;
        RECT 47.575 142.205 47.745 142.635 ;
        RECT 46.040 141.515 46.900 141.665 ;
        RECT 45.615 141.495 46.900 141.515 ;
        RECT 47.070 141.975 47.745 142.205 ;
        RECT 45.615 141.135 46.600 141.495 ;
        RECT 47.070 141.325 47.305 141.975 ;
        RECT 45.265 140.445 45.505 140.965 ;
        RECT 46.430 140.800 46.600 141.135 ;
        RECT 46.770 140.995 47.305 141.325 ;
        RECT 47.085 140.845 47.305 140.995 ;
        RECT 47.475 140.955 47.775 141.805 ;
        RECT 48.005 141.735 49.675 142.825 ;
        RECT 48.005 141.045 48.755 141.565 ;
        RECT 48.925 141.215 49.675 141.735 ;
        RECT 49.845 141.660 50.135 142.825 ;
        RECT 50.305 141.735 51.975 142.825 ;
        RECT 50.305 141.045 51.055 141.565 ;
        RECT 51.225 141.215 51.975 141.735 ;
        RECT 52.145 141.855 52.455 142.655 ;
        RECT 52.625 142.025 52.935 142.825 ;
        RECT 53.105 142.195 53.365 142.655 ;
        RECT 53.535 142.365 53.790 142.825 ;
        RECT 53.965 142.195 54.225 142.655 ;
        RECT 53.105 142.025 54.225 142.195 ;
        RECT 52.145 141.685 53.175 141.855 ;
        RECT 45.675 140.275 46.070 140.770 ;
        RECT 46.430 140.605 46.805 140.800 ;
        RECT 46.635 140.460 46.805 140.605 ;
        RECT 47.085 140.470 47.325 140.845 ;
        RECT 47.495 140.275 47.830 140.780 ;
        RECT 48.005 140.275 49.675 141.045 ;
        RECT 49.845 140.275 50.135 141.000 ;
        RECT 50.305 140.275 51.975 141.045 ;
        RECT 52.145 140.775 52.315 141.685 ;
        RECT 52.485 140.945 52.835 141.515 ;
        RECT 53.005 141.435 53.175 141.685 ;
        RECT 53.965 141.775 54.225 142.025 ;
        RECT 54.395 141.955 54.680 142.825 ;
        RECT 54.905 142.390 60.250 142.825 ;
        RECT 53.965 141.605 54.720 141.775 ;
        RECT 53.005 141.265 54.145 141.435 ;
        RECT 54.315 141.095 54.720 141.605 ;
        RECT 53.070 140.925 54.720 141.095 ;
        RECT 52.145 140.445 52.445 140.775 ;
        RECT 52.615 140.275 52.890 140.755 ;
        RECT 53.070 140.535 53.365 140.925 ;
        RECT 53.535 140.275 53.790 140.755 ;
        RECT 53.965 140.535 54.225 140.925 ;
        RECT 56.490 140.820 56.830 141.650 ;
        RECT 58.310 141.140 58.660 142.390 ;
        RECT 60.425 141.735 63.935 142.825 ;
        RECT 64.105 141.735 65.315 142.825 ;
        RECT 60.425 141.045 62.075 141.565 ;
        RECT 62.245 141.215 63.935 141.735 ;
        RECT 54.395 140.275 54.675 140.755 ;
        RECT 54.905 140.275 60.250 140.820 ;
        RECT 60.425 140.275 63.935 141.045 ;
        RECT 64.105 141.025 64.625 141.565 ;
        RECT 64.795 141.195 65.315 141.735 ;
        RECT 65.485 141.750 65.755 142.655 ;
        RECT 65.925 142.065 66.255 142.825 ;
        RECT 66.435 141.895 66.605 142.655 ;
        RECT 66.865 142.390 72.210 142.825 ;
        RECT 64.105 140.275 65.315 141.025 ;
        RECT 65.485 140.950 65.655 141.750 ;
        RECT 65.940 141.725 66.605 141.895 ;
        RECT 65.940 141.580 66.110 141.725 ;
        RECT 65.825 141.250 66.110 141.580 ;
        RECT 65.940 140.995 66.110 141.250 ;
        RECT 66.345 141.175 66.675 141.545 ;
        RECT 65.485 140.445 65.745 140.950 ;
        RECT 65.940 140.825 66.605 140.995 ;
        RECT 65.925 140.275 66.255 140.655 ;
        RECT 66.435 140.445 66.605 140.825 ;
        RECT 68.450 140.820 68.790 141.650 ;
        RECT 70.270 141.140 70.620 142.390 ;
        RECT 72.385 141.735 74.975 142.825 ;
        RECT 72.385 141.045 73.595 141.565 ;
        RECT 73.765 141.215 74.975 141.735 ;
        RECT 75.605 141.660 75.895 142.825 ;
        RECT 76.525 141.685 76.785 142.825 ;
        RECT 76.955 141.675 77.285 142.655 ;
        RECT 77.455 141.685 77.735 142.825 ;
        RECT 77.905 142.390 83.250 142.825 ;
        RECT 83.425 142.390 88.770 142.825 ;
        RECT 88.945 142.390 94.290 142.825 ;
        RECT 94.465 142.390 99.810 142.825 ;
        RECT 76.545 141.265 76.880 141.515 ;
        RECT 77.050 141.075 77.220 141.675 ;
        RECT 77.390 141.245 77.725 141.515 ;
        RECT 66.865 140.275 72.210 140.820 ;
        RECT 72.385 140.275 74.975 141.045 ;
        RECT 75.605 140.275 75.895 141.000 ;
        RECT 76.525 140.445 77.220 141.075 ;
        RECT 77.425 140.275 77.735 141.075 ;
        RECT 79.490 140.820 79.830 141.650 ;
        RECT 81.310 141.140 81.660 142.390 ;
        RECT 85.010 140.820 85.350 141.650 ;
        RECT 86.830 141.140 87.180 142.390 ;
        RECT 90.530 140.820 90.870 141.650 ;
        RECT 92.350 141.140 92.700 142.390 ;
        RECT 96.050 140.820 96.390 141.650 ;
        RECT 97.870 141.140 98.220 142.390 ;
        RECT 99.985 141.735 101.195 142.825 ;
        RECT 99.985 141.025 100.505 141.565 ;
        RECT 100.675 141.195 101.195 141.735 ;
        RECT 101.365 141.660 101.655 142.825 ;
        RECT 101.825 141.220 102.105 142.655 ;
        RECT 102.275 142.050 102.985 142.825 ;
        RECT 103.155 141.880 103.485 142.655 ;
        RECT 102.335 141.665 103.485 141.880 ;
        RECT 77.905 140.275 83.250 140.820 ;
        RECT 83.425 140.275 88.770 140.820 ;
        RECT 88.945 140.275 94.290 140.820 ;
        RECT 94.465 140.275 99.810 140.820 ;
        RECT 99.985 140.275 101.195 141.025 ;
        RECT 101.365 140.275 101.655 141.000 ;
        RECT 101.825 140.445 102.165 141.220 ;
        RECT 102.335 141.095 102.620 141.665 ;
        RECT 102.805 141.265 103.275 141.495 ;
        RECT 103.680 141.465 103.895 142.580 ;
        RECT 104.075 142.105 104.405 142.825 ;
        RECT 104.185 141.465 104.415 141.805 ;
        RECT 105.055 141.685 105.385 142.825 ;
        RECT 105.915 141.855 106.245 142.640 ;
        RECT 105.565 141.685 106.245 141.855 ;
        RECT 106.885 141.975 107.265 142.655 ;
        RECT 107.855 141.975 108.025 142.825 ;
        RECT 108.195 142.145 108.525 142.655 ;
        RECT 108.695 142.315 108.865 142.825 ;
        RECT 109.035 142.145 109.435 142.655 ;
        RECT 108.195 141.975 109.435 142.145 ;
        RECT 103.445 141.285 103.895 141.465 ;
        RECT 103.445 141.265 103.775 141.285 ;
        RECT 104.085 141.265 104.415 141.465 ;
        RECT 105.045 141.265 105.395 141.515 ;
        RECT 102.335 140.905 103.045 141.095 ;
        RECT 102.745 140.765 103.045 140.905 ;
        RECT 103.235 140.905 104.415 141.095 ;
        RECT 105.565 141.085 105.735 141.685 ;
        RECT 105.905 141.265 106.255 141.515 ;
        RECT 103.235 140.825 103.565 140.905 ;
        RECT 102.745 140.755 103.060 140.765 ;
        RECT 102.745 140.745 103.070 140.755 ;
        RECT 102.745 140.740 103.080 140.745 ;
        RECT 102.335 140.275 102.505 140.735 ;
        RECT 102.745 140.730 103.085 140.740 ;
        RECT 102.745 140.725 103.090 140.730 ;
        RECT 102.745 140.715 103.095 140.725 ;
        RECT 102.745 140.710 103.100 140.715 ;
        RECT 102.745 140.445 103.105 140.710 ;
        RECT 103.735 140.275 103.905 140.735 ;
        RECT 104.075 140.445 104.415 140.905 ;
        RECT 105.055 140.275 105.325 141.085 ;
        RECT 105.495 140.445 105.825 141.085 ;
        RECT 105.995 140.275 106.235 141.085 ;
        RECT 106.885 141.015 107.055 141.975 ;
        RECT 107.225 141.635 108.530 141.805 ;
        RECT 109.615 141.725 109.935 142.655 ;
        RECT 107.225 141.185 107.470 141.635 ;
        RECT 107.640 141.265 108.190 141.465 ;
        RECT 108.360 141.435 108.530 141.635 ;
        RECT 109.305 141.555 109.935 141.725 ;
        RECT 111.030 142.435 111.365 142.655 ;
        RECT 112.370 142.445 112.725 142.825 ;
        RECT 111.030 141.815 111.285 142.435 ;
        RECT 111.535 142.275 111.765 142.315 ;
        RECT 112.895 142.275 113.145 142.655 ;
        RECT 111.535 142.075 113.145 142.275 ;
        RECT 111.535 141.985 111.720 142.075 ;
        RECT 112.310 142.065 113.145 142.075 ;
        RECT 113.395 142.045 113.645 142.825 ;
        RECT 113.815 141.975 114.075 142.655 ;
        RECT 111.875 141.875 112.205 141.905 ;
        RECT 111.875 141.815 113.675 141.875 ;
        RECT 111.030 141.705 113.735 141.815 ;
        RECT 111.030 141.645 112.205 141.705 ;
        RECT 113.535 141.670 113.735 141.705 ;
        RECT 108.360 141.265 108.735 141.435 ;
        RECT 108.905 141.015 109.135 141.515 ;
        RECT 106.885 140.845 109.135 141.015 ;
        RECT 106.935 140.275 107.265 140.665 ;
        RECT 107.435 140.525 107.605 140.845 ;
        RECT 109.305 140.675 109.475 141.555 ;
        RECT 111.025 141.265 111.515 141.465 ;
        RECT 111.705 141.265 112.180 141.475 ;
        RECT 107.775 140.275 108.105 140.665 ;
        RECT 108.520 140.505 109.475 140.675 ;
        RECT 109.645 140.275 109.935 141.110 ;
        RECT 111.030 140.275 111.485 141.040 ;
        RECT 111.960 140.865 112.180 141.265 ;
        RECT 112.425 141.265 112.755 141.475 ;
        RECT 112.425 140.865 112.635 141.265 ;
        RECT 112.925 141.230 113.335 141.535 ;
        RECT 113.565 141.095 113.735 141.670 ;
        RECT 113.465 140.975 113.735 141.095 ;
        RECT 112.890 140.930 113.735 140.975 ;
        RECT 112.890 140.805 113.645 140.930 ;
        RECT 112.890 140.655 113.060 140.805 ;
        RECT 113.905 140.785 114.075 141.975 ;
        RECT 114.305 141.765 114.635 142.610 ;
        RECT 114.805 141.815 114.975 142.825 ;
        RECT 115.145 142.095 115.485 142.655 ;
        RECT 115.715 142.325 116.030 142.825 ;
        RECT 116.210 142.355 117.095 142.525 ;
        RECT 114.245 141.685 114.635 141.765 ;
        RECT 115.145 141.720 116.040 142.095 ;
        RECT 114.245 141.635 114.460 141.685 ;
        RECT 114.245 141.055 114.415 141.635 ;
        RECT 115.145 141.515 115.335 141.720 ;
        RECT 116.210 141.515 116.380 142.355 ;
        RECT 117.320 142.325 117.570 142.655 ;
        RECT 114.585 141.185 115.335 141.515 ;
        RECT 115.505 141.185 116.380 141.515 ;
        RECT 114.245 141.015 114.470 141.055 ;
        RECT 115.135 141.015 115.335 141.185 ;
        RECT 114.245 140.930 114.625 141.015 ;
        RECT 113.845 140.775 114.075 140.785 ;
        RECT 111.760 140.445 113.060 140.655 ;
        RECT 113.315 140.275 113.645 140.635 ;
        RECT 113.815 140.445 114.075 140.775 ;
        RECT 114.295 140.495 114.625 140.930 ;
        RECT 114.795 140.275 114.965 140.885 ;
        RECT 115.135 140.490 115.465 141.015 ;
        RECT 115.725 140.275 115.935 140.805 ;
        RECT 116.210 140.725 116.380 141.185 ;
        RECT 116.550 141.225 116.870 142.185 ;
        RECT 117.040 141.435 117.230 142.155 ;
        RECT 117.400 141.255 117.570 142.325 ;
        RECT 117.740 142.025 117.910 142.825 ;
        RECT 118.080 142.380 119.185 142.550 ;
        RECT 118.080 141.765 118.250 142.380 ;
        RECT 119.395 142.230 119.645 142.655 ;
        RECT 119.815 142.365 120.080 142.825 ;
        RECT 118.420 141.845 118.950 142.210 ;
        RECT 119.395 142.100 119.700 142.230 ;
        RECT 117.740 141.675 118.250 141.765 ;
        RECT 117.740 141.505 118.610 141.675 ;
        RECT 117.740 141.435 117.910 141.505 ;
        RECT 118.030 141.255 118.230 141.285 ;
        RECT 116.550 140.895 117.015 141.225 ;
        RECT 117.400 140.955 118.230 141.255 ;
        RECT 117.400 140.725 117.570 140.955 ;
        RECT 116.210 140.555 116.995 140.725 ;
        RECT 117.165 140.555 117.570 140.725 ;
        RECT 117.750 140.275 118.120 140.775 ;
        RECT 118.440 140.725 118.610 141.505 ;
        RECT 118.780 141.145 118.950 141.845 ;
        RECT 119.120 141.315 119.360 141.910 ;
        RECT 118.780 140.925 119.305 141.145 ;
        RECT 119.530 140.995 119.700 142.100 ;
        RECT 119.475 140.865 119.700 140.995 ;
        RECT 119.870 140.905 120.150 141.855 ;
        RECT 119.475 140.725 119.645 140.865 ;
        RECT 118.440 140.555 119.115 140.725 ;
        RECT 119.310 140.555 119.645 140.725 ;
        RECT 119.815 140.275 120.065 140.735 ;
        RECT 120.320 140.535 120.505 142.655 ;
        RECT 120.675 142.325 121.005 142.825 ;
        RECT 121.175 142.155 121.345 142.655 ;
        RECT 121.605 142.390 126.950 142.825 ;
        RECT 120.680 141.985 121.345 142.155 ;
        RECT 120.680 140.995 120.910 141.985 ;
        RECT 121.080 141.165 121.430 141.815 ;
        RECT 120.680 140.825 121.345 140.995 ;
        RECT 120.675 140.275 121.005 140.655 ;
        RECT 121.175 140.535 121.345 140.825 ;
        RECT 123.190 140.820 123.530 141.650 ;
        RECT 125.010 141.140 125.360 142.390 ;
        RECT 127.125 141.660 127.415 142.825 ;
        RECT 127.585 142.390 132.930 142.825 ;
        RECT 133.105 142.390 138.450 142.825 ;
        RECT 138.625 142.390 143.970 142.825 ;
        RECT 121.605 140.275 126.950 140.820 ;
        RECT 127.125 140.275 127.415 141.000 ;
        RECT 129.170 140.820 129.510 141.650 ;
        RECT 130.990 141.140 131.340 142.390 ;
        RECT 134.690 140.820 135.030 141.650 ;
        RECT 136.510 141.140 136.860 142.390 ;
        RECT 140.210 140.820 140.550 141.650 ;
        RECT 142.030 141.140 142.380 142.390 ;
        RECT 144.145 141.735 147.655 142.825 ;
        RECT 147.825 141.735 149.035 142.825 ;
        RECT 144.145 141.045 145.795 141.565 ;
        RECT 145.965 141.215 147.655 141.735 ;
        RECT 127.585 140.275 132.930 140.820 ;
        RECT 133.105 140.275 138.450 140.820 ;
        RECT 138.625 140.275 143.970 140.820 ;
        RECT 144.145 140.275 147.655 141.045 ;
        RECT 147.825 141.025 148.345 141.565 ;
        RECT 148.515 141.195 149.035 141.735 ;
        RECT 149.205 141.735 150.415 142.825 ;
        RECT 149.205 141.195 149.725 141.735 ;
        RECT 149.895 141.025 150.415 141.565 ;
        RECT 147.825 140.275 149.035 141.025 ;
        RECT 149.205 140.275 150.415 141.025 ;
        RECT 11.120 140.105 150.500 140.275 ;
        RECT 11.205 139.355 12.415 140.105 ;
        RECT 11.205 138.815 11.725 139.355 ;
        RECT 12.585 139.335 15.175 140.105 ;
        RECT 15.895 139.555 16.065 139.845 ;
        RECT 16.235 139.725 16.565 140.105 ;
        RECT 15.895 139.385 16.560 139.555 ;
        RECT 11.895 138.645 12.415 139.185 ;
        RECT 12.585 138.815 13.795 139.335 ;
        RECT 13.965 138.645 15.175 139.165 ;
        RECT 11.205 137.555 12.415 138.645 ;
        RECT 12.585 137.555 15.175 138.645 ;
        RECT 15.810 138.565 16.160 139.215 ;
        RECT 16.330 138.395 16.560 139.385 ;
        RECT 15.895 138.225 16.560 138.395 ;
        RECT 15.895 137.725 16.065 138.225 ;
        RECT 16.235 137.555 16.565 138.055 ;
        RECT 16.735 137.725 16.920 139.845 ;
        RECT 17.175 139.645 17.425 140.105 ;
        RECT 17.595 139.655 17.930 139.825 ;
        RECT 18.125 139.655 18.800 139.825 ;
        RECT 17.595 139.515 17.765 139.655 ;
        RECT 17.090 138.525 17.370 139.475 ;
        RECT 17.540 139.385 17.765 139.515 ;
        RECT 17.540 138.280 17.710 139.385 ;
        RECT 17.935 139.235 18.460 139.455 ;
        RECT 17.880 138.470 18.120 139.065 ;
        RECT 18.290 138.535 18.460 139.235 ;
        RECT 18.630 138.875 18.800 139.655 ;
        RECT 19.120 139.605 19.490 140.105 ;
        RECT 19.670 139.655 20.075 139.825 ;
        RECT 20.245 139.655 21.030 139.825 ;
        RECT 19.670 139.425 19.840 139.655 ;
        RECT 19.010 139.125 19.840 139.425 ;
        RECT 20.225 139.155 20.690 139.485 ;
        RECT 19.010 139.095 19.210 139.125 ;
        RECT 19.330 138.875 19.500 138.945 ;
        RECT 18.630 138.705 19.500 138.875 ;
        RECT 18.990 138.615 19.500 138.705 ;
        RECT 17.540 138.150 17.845 138.280 ;
        RECT 18.290 138.170 18.820 138.535 ;
        RECT 17.160 137.555 17.425 138.015 ;
        RECT 17.595 137.725 17.845 138.150 ;
        RECT 18.990 138.000 19.160 138.615 ;
        RECT 18.055 137.830 19.160 138.000 ;
        RECT 19.330 137.555 19.500 138.355 ;
        RECT 19.670 138.055 19.840 139.125 ;
        RECT 20.010 138.225 20.200 138.945 ;
        RECT 20.370 138.195 20.690 139.155 ;
        RECT 20.860 139.195 21.030 139.655 ;
        RECT 21.305 139.575 21.515 140.105 ;
        RECT 21.775 139.365 22.105 139.890 ;
        RECT 22.275 139.495 22.445 140.105 ;
        RECT 22.615 139.450 22.945 139.885 ;
        RECT 22.615 139.365 22.995 139.450 ;
        RECT 21.905 139.195 22.105 139.365 ;
        RECT 22.770 139.325 22.995 139.365 ;
        RECT 20.860 138.865 21.735 139.195 ;
        RECT 21.905 138.865 22.655 139.195 ;
        RECT 19.670 137.725 19.920 138.055 ;
        RECT 20.860 138.025 21.030 138.865 ;
        RECT 21.905 138.660 22.095 138.865 ;
        RECT 22.825 138.745 22.995 139.325 ;
        RECT 22.780 138.695 22.995 138.745 ;
        RECT 21.200 138.285 22.095 138.660 ;
        RECT 22.605 138.615 22.995 138.695 ;
        RECT 23.165 139.365 23.630 139.910 ;
        RECT 20.145 137.855 21.030 138.025 ;
        RECT 21.210 137.555 21.525 138.055 ;
        RECT 21.755 137.725 22.095 138.285 ;
        RECT 22.265 137.555 22.435 138.565 ;
        RECT 22.605 137.770 22.935 138.615 ;
        RECT 23.165 138.405 23.335 139.365 ;
        RECT 24.135 139.285 24.305 140.105 ;
        RECT 24.475 139.455 24.805 139.935 ;
        RECT 24.975 139.715 25.325 140.105 ;
        RECT 25.495 139.535 25.725 139.935 ;
        RECT 25.215 139.455 25.725 139.535 ;
        RECT 24.475 139.365 25.725 139.455 ;
        RECT 25.895 139.365 26.215 139.845 ;
        RECT 24.475 139.285 25.385 139.365 ;
        RECT 23.505 138.745 23.750 139.195 ;
        RECT 24.010 138.915 24.705 139.115 ;
        RECT 24.875 138.945 25.475 139.115 ;
        RECT 24.875 138.745 25.045 138.945 ;
        RECT 25.705 138.775 25.875 139.195 ;
        RECT 23.505 138.575 25.045 138.745 ;
        RECT 25.215 138.605 25.875 138.775 ;
        RECT 25.215 138.405 25.385 138.605 ;
        RECT 26.045 138.435 26.215 139.365 ;
        RECT 26.865 139.475 27.195 139.935 ;
        RECT 27.375 139.645 27.545 140.105 ;
        RECT 27.725 139.475 28.055 139.935 ;
        RECT 28.285 139.645 28.455 140.105 ;
        RECT 28.695 139.765 29.885 139.935 ;
        RECT 28.695 139.475 29.025 139.765 ;
        RECT 29.575 139.595 29.885 139.765 ;
        RECT 30.065 139.605 30.325 139.935 ;
        RECT 30.495 139.745 30.825 140.105 ;
        RECT 31.080 139.725 32.380 139.935 ;
        RECT 26.865 139.305 29.025 139.475 ;
        RECT 26.880 138.745 27.210 139.135 ;
        RECT 27.380 138.915 28.180 139.115 ;
        RECT 28.360 138.745 28.855 139.115 ;
        RECT 26.880 138.575 28.915 138.745 ;
        RECT 23.165 138.235 25.385 138.405 ;
        RECT 25.555 138.235 26.215 138.435 ;
        RECT 29.195 138.405 29.405 139.595 ;
        RECT 29.575 138.790 29.890 139.425 ;
        RECT 23.165 137.555 23.465 138.065 ;
        RECT 23.635 137.725 23.965 138.235 ;
        RECT 25.555 138.065 25.725 138.235 ;
        RECT 24.135 137.555 24.765 138.065 ;
        RECT 25.345 137.895 25.725 138.065 ;
        RECT 25.895 137.555 26.195 138.065 ;
        RECT 26.865 137.555 27.195 138.405 ;
        RECT 27.365 137.895 27.585 138.405 ;
        RECT 27.755 138.225 29.405 138.405 ;
        RECT 27.755 138.065 28.055 138.225 ;
        RECT 28.285 137.895 28.475 138.055 ;
        RECT 27.365 137.725 28.475 137.895 ;
        RECT 28.670 137.555 29.000 138.015 ;
        RECT 29.170 137.725 29.405 138.225 ;
        RECT 29.575 137.555 29.885 138.620 ;
        RECT 30.065 138.405 30.235 139.605 ;
        RECT 31.080 139.575 31.250 139.725 ;
        RECT 30.495 139.450 31.250 139.575 ;
        RECT 30.405 139.405 31.250 139.450 ;
        RECT 30.405 139.285 30.675 139.405 ;
        RECT 30.405 138.710 30.575 139.285 ;
        RECT 30.805 138.845 31.215 139.150 ;
        RECT 31.505 139.115 31.715 139.515 ;
        RECT 31.385 138.905 31.715 139.115 ;
        RECT 31.960 139.115 32.180 139.515 ;
        RECT 32.655 139.340 33.110 140.105 ;
        RECT 33.285 139.335 36.795 140.105 ;
        RECT 36.965 139.380 37.255 140.105 ;
        RECT 37.515 139.625 37.815 140.105 ;
        RECT 37.985 139.455 38.245 139.910 ;
        RECT 38.415 139.625 38.675 140.105 ;
        RECT 38.855 139.455 39.115 139.910 ;
        RECT 39.285 139.625 39.535 140.105 ;
        RECT 39.715 139.455 39.975 139.910 ;
        RECT 40.145 139.625 40.395 140.105 ;
        RECT 40.575 139.455 40.835 139.910 ;
        RECT 41.005 139.625 41.250 140.105 ;
        RECT 41.420 139.455 41.695 139.910 ;
        RECT 41.865 139.625 42.110 140.105 ;
        RECT 42.280 139.455 42.540 139.910 ;
        RECT 42.710 139.625 42.970 140.105 ;
        RECT 43.140 139.455 43.400 139.910 ;
        RECT 43.570 139.625 43.830 140.105 ;
        RECT 44.000 139.455 44.260 139.910 ;
        RECT 44.430 139.545 44.690 140.105 ;
        RECT 31.960 138.905 32.435 139.115 ;
        RECT 32.625 138.915 33.115 139.115 ;
        RECT 33.285 138.815 34.935 139.335 ;
        RECT 37.515 139.285 44.260 139.455 ;
        RECT 30.405 138.675 30.605 138.710 ;
        RECT 31.935 138.675 33.110 138.735 ;
        RECT 30.405 138.565 33.110 138.675 ;
        RECT 35.105 138.645 36.795 139.165 ;
        RECT 30.465 138.505 32.265 138.565 ;
        RECT 31.935 138.475 32.265 138.505 ;
        RECT 30.065 137.725 30.325 138.405 ;
        RECT 30.495 137.555 30.745 138.335 ;
        RECT 30.995 138.305 31.830 138.315 ;
        RECT 32.420 138.305 32.605 138.395 ;
        RECT 30.995 138.105 32.605 138.305 ;
        RECT 30.995 137.725 31.245 138.105 ;
        RECT 32.375 138.065 32.605 138.105 ;
        RECT 32.855 137.945 33.110 138.565 ;
        RECT 31.415 137.555 31.770 137.935 ;
        RECT 32.775 137.725 33.110 137.945 ;
        RECT 33.285 137.555 36.795 138.645 ;
        RECT 36.965 137.555 37.255 138.720 ;
        RECT 37.515 138.695 38.680 139.285 ;
        RECT 44.860 139.115 45.110 139.925 ;
        RECT 45.290 139.580 45.550 140.105 ;
        RECT 45.720 139.115 45.970 139.925 ;
        RECT 46.150 139.595 46.455 140.105 ;
        RECT 47.545 139.595 47.850 140.105 ;
        RECT 38.850 138.865 45.970 139.115 ;
        RECT 46.140 138.865 46.455 139.425 ;
        RECT 47.545 138.865 47.860 139.425 ;
        RECT 48.030 139.115 48.280 139.925 ;
        RECT 48.450 139.580 48.710 140.105 ;
        RECT 48.890 139.115 49.140 139.925 ;
        RECT 49.310 139.545 49.570 140.105 ;
        RECT 49.740 139.455 50.000 139.910 ;
        RECT 50.170 139.625 50.430 140.105 ;
        RECT 50.600 139.455 50.860 139.910 ;
        RECT 51.030 139.625 51.290 140.105 ;
        RECT 51.460 139.455 51.720 139.910 ;
        RECT 51.890 139.625 52.135 140.105 ;
        RECT 52.305 139.455 52.580 139.910 ;
        RECT 52.750 139.625 52.995 140.105 ;
        RECT 53.165 139.455 53.425 139.910 ;
        RECT 53.605 139.625 53.855 140.105 ;
        RECT 54.025 139.455 54.285 139.910 ;
        RECT 54.465 139.625 54.715 140.105 ;
        RECT 54.885 139.455 55.145 139.910 ;
        RECT 55.325 139.625 55.585 140.105 ;
        RECT 55.755 139.455 56.015 139.910 ;
        RECT 56.185 139.625 56.485 140.105 ;
        RECT 49.740 139.425 56.485 139.455 ;
        RECT 49.740 139.285 56.515 139.425 ;
        RECT 55.320 139.255 56.515 139.285 ;
        RECT 48.030 138.865 55.150 139.115 ;
        RECT 37.515 138.470 44.260 138.695 ;
        RECT 37.515 137.555 37.785 138.300 ;
        RECT 37.955 137.730 38.245 138.470 ;
        RECT 38.855 138.455 44.260 138.470 ;
        RECT 38.415 137.560 38.670 138.285 ;
        RECT 38.855 137.730 39.115 138.455 ;
        RECT 39.285 137.560 39.530 138.285 ;
        RECT 39.715 137.730 39.975 138.455 ;
        RECT 40.145 137.560 40.390 138.285 ;
        RECT 40.575 137.730 40.835 138.455 ;
        RECT 41.005 137.560 41.250 138.285 ;
        RECT 41.420 137.730 41.680 138.455 ;
        RECT 41.850 137.560 42.110 138.285 ;
        RECT 42.280 137.730 42.540 138.455 ;
        RECT 42.710 137.560 42.970 138.285 ;
        RECT 43.140 137.730 43.400 138.455 ;
        RECT 43.570 137.560 43.830 138.285 ;
        RECT 44.000 137.730 44.260 138.455 ;
        RECT 44.430 137.560 44.690 138.355 ;
        RECT 44.860 137.730 45.110 138.865 ;
        RECT 38.415 137.555 44.690 137.560 ;
        RECT 45.290 137.555 45.550 138.365 ;
        RECT 45.725 137.725 45.970 138.865 ;
        RECT 46.150 137.555 46.445 138.365 ;
        RECT 47.555 137.555 47.850 138.365 ;
        RECT 48.030 137.725 48.275 138.865 ;
        RECT 48.450 137.555 48.710 138.365 ;
        RECT 48.890 137.730 49.140 138.865 ;
        RECT 55.320 138.695 56.485 139.255 ;
        RECT 49.740 138.470 56.485 138.695 ;
        RECT 49.740 138.455 55.145 138.470 ;
        RECT 49.310 137.560 49.570 138.355 ;
        RECT 49.740 137.730 50.000 138.455 ;
        RECT 50.170 137.560 50.430 138.285 ;
        RECT 50.600 137.730 50.860 138.455 ;
        RECT 51.030 137.560 51.290 138.285 ;
        RECT 51.460 137.730 51.720 138.455 ;
        RECT 51.890 137.560 52.150 138.285 ;
        RECT 52.320 137.730 52.580 138.455 ;
        RECT 52.750 137.560 52.995 138.285 ;
        RECT 53.165 137.730 53.425 138.455 ;
        RECT 53.610 137.560 53.855 138.285 ;
        RECT 54.025 137.730 54.285 138.455 ;
        RECT 54.470 137.560 54.715 138.285 ;
        RECT 54.885 137.730 55.145 138.455 ;
        RECT 55.330 137.560 55.585 138.285 ;
        RECT 55.755 137.730 56.045 138.470 ;
        RECT 49.310 137.555 55.585 137.560 ;
        RECT 56.215 137.555 56.485 138.300 ;
        RECT 56.755 137.735 57.015 139.925 ;
        RECT 57.275 139.735 57.945 140.105 ;
        RECT 58.125 139.555 58.435 139.925 ;
        RECT 57.205 139.355 58.435 139.555 ;
        RECT 57.205 138.685 57.495 139.355 ;
        RECT 58.615 139.175 58.845 139.815 ;
        RECT 59.025 139.375 59.315 140.105 ;
        RECT 59.520 139.535 59.775 139.885 ;
        RECT 59.945 139.705 60.275 140.105 ;
        RECT 60.445 139.535 60.615 139.885 ;
        RECT 60.785 139.705 61.165 140.105 ;
        RECT 59.520 139.365 61.185 139.535 ;
        RECT 61.355 139.430 61.630 139.775 ;
        RECT 61.015 139.195 61.185 139.365 ;
        RECT 57.675 138.865 58.140 139.175 ;
        RECT 58.320 138.865 58.845 139.175 ;
        RECT 59.025 138.865 59.325 139.195 ;
        RECT 59.505 138.865 59.850 139.195 ;
        RECT 60.020 138.865 60.845 139.195 ;
        RECT 61.015 138.865 61.290 139.195 ;
        RECT 57.205 138.465 57.975 138.685 ;
        RECT 57.185 137.555 57.525 138.285 ;
        RECT 57.705 137.735 57.975 138.465 ;
        RECT 58.155 138.445 59.315 138.685 ;
        RECT 58.155 137.735 58.385 138.445 ;
        RECT 58.555 137.555 58.885 138.265 ;
        RECT 59.055 137.735 59.315 138.445 ;
        RECT 59.525 138.405 59.850 138.695 ;
        RECT 60.020 138.575 60.215 138.865 ;
        RECT 61.015 138.695 61.185 138.865 ;
        RECT 61.460 138.695 61.630 139.430 ;
        RECT 62.725 139.380 63.015 140.105 ;
        RECT 63.185 139.335 64.855 140.105 ;
        RECT 65.025 139.605 65.325 139.935 ;
        RECT 65.495 139.625 65.770 140.105 ;
        RECT 63.185 138.815 63.935 139.335 ;
        RECT 60.525 138.525 61.185 138.695 ;
        RECT 60.525 138.405 60.695 138.525 ;
        RECT 59.525 138.235 60.695 138.405 ;
        RECT 59.505 137.775 60.695 138.065 ;
        RECT 60.865 137.555 61.145 138.355 ;
        RECT 61.355 137.725 61.630 138.695 ;
        RECT 62.725 137.555 63.015 138.720 ;
        RECT 64.105 138.645 64.855 139.165 ;
        RECT 63.185 137.555 64.855 138.645 ;
        RECT 65.025 138.695 65.195 139.605 ;
        RECT 65.950 139.455 66.245 139.845 ;
        RECT 66.415 139.625 66.670 140.105 ;
        RECT 66.845 139.455 67.105 139.845 ;
        RECT 67.275 139.625 67.555 140.105 ;
        RECT 65.365 138.865 65.715 139.435 ;
        RECT 65.950 139.285 67.600 139.455 ;
        RECT 65.885 138.945 67.025 139.115 ;
        RECT 65.885 138.695 66.055 138.945 ;
        RECT 67.195 138.775 67.600 139.285 ;
        RECT 67.785 139.335 71.295 140.105 ;
        RECT 71.465 139.355 72.675 140.105 ;
        RECT 72.845 139.365 73.310 139.910 ;
        RECT 67.785 138.815 69.435 139.335 ;
        RECT 65.025 138.525 66.055 138.695 ;
        RECT 66.845 138.605 67.600 138.775 ;
        RECT 69.605 138.645 71.295 139.165 ;
        RECT 71.465 138.815 71.985 139.355 ;
        RECT 72.155 138.645 72.675 139.185 ;
        RECT 65.025 137.725 65.335 138.525 ;
        RECT 66.845 138.355 67.105 138.605 ;
        RECT 65.505 137.555 65.815 138.355 ;
        RECT 65.985 138.185 67.105 138.355 ;
        RECT 65.985 137.725 66.245 138.185 ;
        RECT 66.415 137.555 66.670 138.015 ;
        RECT 66.845 137.725 67.105 138.185 ;
        RECT 67.275 137.555 67.560 138.425 ;
        RECT 67.785 137.555 71.295 138.645 ;
        RECT 71.465 137.555 72.675 138.645 ;
        RECT 72.845 138.405 73.015 139.365 ;
        RECT 73.815 139.285 73.985 140.105 ;
        RECT 74.155 139.455 74.485 139.935 ;
        RECT 74.655 139.715 75.005 140.105 ;
        RECT 75.175 139.535 75.405 139.935 ;
        RECT 74.895 139.455 75.405 139.535 ;
        RECT 74.155 139.365 75.405 139.455 ;
        RECT 75.575 139.365 75.895 139.845 ;
        RECT 74.155 139.285 75.065 139.365 ;
        RECT 73.185 138.745 73.430 139.195 ;
        RECT 73.690 138.915 74.385 139.115 ;
        RECT 74.555 138.945 75.155 139.115 ;
        RECT 74.555 138.745 74.725 138.945 ;
        RECT 75.385 138.775 75.555 139.195 ;
        RECT 73.185 138.575 74.725 138.745 ;
        RECT 74.895 138.605 75.555 138.775 ;
        RECT 74.895 138.405 75.065 138.605 ;
        RECT 75.725 138.435 75.895 139.365 ;
        RECT 72.845 138.235 75.065 138.405 ;
        RECT 75.235 138.235 75.895 138.435 ;
        RECT 76.100 139.365 76.715 139.935 ;
        RECT 76.885 139.595 77.100 140.105 ;
        RECT 77.330 139.595 77.610 139.925 ;
        RECT 77.790 139.595 78.030 140.105 ;
        RECT 78.830 139.630 79.165 139.890 ;
        RECT 79.335 139.705 79.665 140.105 ;
        RECT 79.835 139.705 81.450 139.875 ;
        RECT 76.100 138.345 76.415 139.365 ;
        RECT 76.585 138.695 76.755 139.195 ;
        RECT 77.005 138.865 77.270 139.425 ;
        RECT 77.440 138.695 77.610 139.595 ;
        RECT 77.780 138.865 78.135 139.425 ;
        RECT 76.585 138.525 78.010 138.695 ;
        RECT 72.845 137.555 73.145 138.065 ;
        RECT 73.315 137.725 73.645 138.235 ;
        RECT 75.235 138.065 75.405 138.235 ;
        RECT 73.815 137.555 74.445 138.065 ;
        RECT 75.025 137.895 75.405 138.065 ;
        RECT 75.575 137.555 75.875 138.065 ;
        RECT 76.100 137.725 76.635 138.345 ;
        RECT 76.805 137.555 77.135 138.355 ;
        RECT 77.620 138.350 78.010 138.525 ;
        RECT 78.830 138.275 79.085 139.630 ;
        RECT 79.835 139.535 80.005 139.705 ;
        RECT 79.445 139.365 80.005 139.535 ;
        RECT 79.445 139.195 79.615 139.365 ;
        RECT 79.310 138.865 79.615 139.195 ;
        RECT 79.810 139.085 80.060 139.195 ;
        RECT 80.270 139.085 80.540 139.525 ;
        RECT 80.730 139.085 81.020 139.525 ;
        RECT 79.805 138.915 80.060 139.085 ;
        RECT 80.265 138.915 80.540 139.085 ;
        RECT 80.725 138.915 81.020 139.085 ;
        RECT 79.810 138.865 80.060 138.915 ;
        RECT 80.270 138.865 80.540 138.915 ;
        RECT 80.730 138.865 81.020 138.915 ;
        RECT 81.190 138.865 81.610 139.530 ;
        RECT 81.995 139.385 82.325 140.105 ;
        RECT 82.505 139.335 84.175 140.105 ;
        RECT 84.545 139.475 84.875 139.835 ;
        RECT 85.495 139.645 85.745 140.105 ;
        RECT 85.915 139.645 86.475 139.935 ;
        RECT 81.920 138.865 82.270 139.195 ;
        RECT 79.445 138.695 79.615 138.865 ;
        RECT 82.065 138.745 82.270 138.865 ;
        RECT 82.505 138.815 83.255 139.335 ;
        RECT 84.545 139.285 85.935 139.475 ;
        RECT 85.765 139.195 85.935 139.285 ;
        RECT 79.445 138.525 81.815 138.695 ;
        RECT 82.065 138.575 82.275 138.745 ;
        RECT 83.425 138.645 84.175 139.165 ;
        RECT 78.830 137.765 79.165 138.275 ;
        RECT 79.415 137.555 79.745 138.355 ;
        RECT 79.990 138.145 81.415 138.315 ;
        RECT 79.990 137.725 80.275 138.145 ;
        RECT 80.530 137.555 80.860 137.975 ;
        RECT 81.085 137.895 81.415 138.145 ;
        RECT 81.645 138.065 81.815 138.525 ;
        RECT 82.075 137.895 82.245 138.395 ;
        RECT 81.085 137.725 82.245 137.895 ;
        RECT 82.505 137.555 84.175 138.645 ;
        RECT 84.360 138.865 85.035 139.115 ;
        RECT 85.255 138.865 85.595 139.115 ;
        RECT 85.765 138.865 86.055 139.195 ;
        RECT 84.360 138.505 84.625 138.865 ;
        RECT 85.765 138.615 85.935 138.865 ;
        RECT 84.995 138.445 85.935 138.615 ;
        RECT 84.545 137.555 84.825 138.225 ;
        RECT 84.995 137.895 85.295 138.445 ;
        RECT 86.225 138.275 86.475 139.645 ;
        RECT 86.655 139.295 86.925 140.105 ;
        RECT 87.095 139.295 87.425 139.935 ;
        RECT 87.595 139.295 87.835 140.105 ;
        RECT 88.485 139.380 88.775 140.105 ;
        RECT 88.965 139.295 89.205 140.105 ;
        RECT 89.375 139.295 89.705 139.935 ;
        RECT 89.875 139.295 90.145 140.105 ;
        RECT 90.325 139.355 91.535 140.105 ;
        RECT 91.755 139.450 92.085 139.885 ;
        RECT 92.255 139.495 92.425 140.105 ;
        RECT 91.705 139.365 92.085 139.450 ;
        RECT 92.595 139.365 92.925 139.890 ;
        RECT 93.185 139.575 93.395 140.105 ;
        RECT 93.670 139.655 94.455 139.825 ;
        RECT 94.625 139.655 95.030 139.825 ;
        RECT 86.645 138.865 86.995 139.115 ;
        RECT 87.165 138.695 87.335 139.295 ;
        RECT 87.505 138.865 87.855 139.115 ;
        RECT 88.945 138.865 89.295 139.115 ;
        RECT 85.495 137.555 85.825 138.275 ;
        RECT 86.015 137.725 86.475 138.275 ;
        RECT 86.655 137.555 86.985 138.695 ;
        RECT 87.165 138.525 87.845 138.695 ;
        RECT 87.515 137.740 87.845 138.525 ;
        RECT 88.485 137.555 88.775 138.720 ;
        RECT 89.465 138.695 89.635 139.295 ;
        RECT 89.805 138.865 90.155 139.115 ;
        RECT 90.325 138.815 90.845 139.355 ;
        RECT 91.705 139.325 91.930 139.365 ;
        RECT 88.955 138.525 89.635 138.695 ;
        RECT 88.955 137.740 89.285 138.525 ;
        RECT 89.815 137.555 90.145 138.695 ;
        RECT 91.015 138.645 91.535 139.185 ;
        RECT 90.325 137.555 91.535 138.645 ;
        RECT 91.705 138.745 91.875 139.325 ;
        RECT 92.595 139.195 92.795 139.365 ;
        RECT 93.670 139.195 93.840 139.655 ;
        RECT 92.045 138.865 92.795 139.195 ;
        RECT 92.965 138.865 93.840 139.195 ;
        RECT 91.705 138.695 91.920 138.745 ;
        RECT 91.705 138.615 92.095 138.695 ;
        RECT 91.765 137.770 92.095 138.615 ;
        RECT 92.605 138.660 92.795 138.865 ;
        RECT 92.265 137.555 92.435 138.565 ;
        RECT 92.605 138.285 93.500 138.660 ;
        RECT 92.605 137.725 92.945 138.285 ;
        RECT 93.175 137.555 93.490 138.055 ;
        RECT 93.670 138.025 93.840 138.865 ;
        RECT 94.010 139.155 94.475 139.485 ;
        RECT 94.860 139.425 95.030 139.655 ;
        RECT 95.210 139.605 95.580 140.105 ;
        RECT 95.900 139.655 96.575 139.825 ;
        RECT 96.770 139.655 97.105 139.825 ;
        RECT 94.010 138.195 94.330 139.155 ;
        RECT 94.860 139.125 95.690 139.425 ;
        RECT 94.500 138.225 94.690 138.945 ;
        RECT 94.860 138.055 95.030 139.125 ;
        RECT 95.490 139.095 95.690 139.125 ;
        RECT 95.200 138.875 95.370 138.945 ;
        RECT 95.900 138.875 96.070 139.655 ;
        RECT 96.935 139.515 97.105 139.655 ;
        RECT 97.275 139.645 97.525 140.105 ;
        RECT 95.200 138.705 96.070 138.875 ;
        RECT 96.240 139.235 96.765 139.455 ;
        RECT 96.935 139.385 97.160 139.515 ;
        RECT 95.200 138.615 95.710 138.705 ;
        RECT 93.670 137.855 94.555 138.025 ;
        RECT 94.780 137.725 95.030 138.055 ;
        RECT 95.200 137.555 95.370 138.355 ;
        RECT 95.540 138.000 95.710 138.615 ;
        RECT 96.240 138.535 96.410 139.235 ;
        RECT 95.880 138.170 96.410 138.535 ;
        RECT 96.580 138.470 96.820 139.065 ;
        RECT 96.990 138.280 97.160 139.385 ;
        RECT 97.330 138.525 97.610 139.475 ;
        RECT 96.855 138.150 97.160 138.280 ;
        RECT 95.540 137.830 96.645 138.000 ;
        RECT 96.855 137.725 97.105 138.150 ;
        RECT 97.275 137.555 97.540 138.015 ;
        RECT 97.780 137.725 97.965 139.845 ;
        RECT 98.135 139.725 98.465 140.105 ;
        RECT 98.635 139.555 98.805 139.845 ;
        RECT 98.140 139.385 98.805 139.555 ;
        RECT 98.140 138.395 98.370 139.385 ;
        RECT 99.065 139.355 100.275 140.105 ;
        RECT 100.455 139.380 100.785 139.890 ;
        RECT 100.955 139.705 101.285 140.105 ;
        RECT 102.335 139.535 102.665 139.875 ;
        RECT 102.835 139.705 103.165 140.105 ;
        RECT 103.670 139.600 104.005 140.105 ;
        RECT 104.175 139.535 104.415 139.910 ;
        RECT 104.695 139.775 104.865 139.920 ;
        RECT 104.695 139.580 105.070 139.775 ;
        RECT 105.430 139.610 105.825 140.105 ;
        RECT 98.540 138.565 98.890 139.215 ;
        RECT 99.065 138.815 99.585 139.355 ;
        RECT 99.755 138.645 100.275 139.185 ;
        RECT 98.140 138.225 98.805 138.395 ;
        RECT 98.135 137.555 98.465 138.055 ;
        RECT 98.635 137.725 98.805 138.225 ;
        RECT 99.065 137.555 100.275 138.645 ;
        RECT 100.455 138.615 100.645 139.380 ;
        RECT 100.955 139.365 103.320 139.535 ;
        RECT 100.955 139.195 101.125 139.365 ;
        RECT 100.815 138.865 101.125 139.195 ;
        RECT 101.295 138.865 101.600 139.195 ;
        RECT 100.455 137.765 100.785 138.615 ;
        RECT 100.955 137.555 101.205 138.695 ;
        RECT 101.385 138.535 101.600 138.865 ;
        RECT 101.775 138.535 102.060 139.195 ;
        RECT 102.255 138.535 102.520 139.195 ;
        RECT 102.735 138.535 102.980 139.195 ;
        RECT 103.150 138.365 103.320 139.365 ;
        RECT 103.725 138.575 104.025 139.425 ;
        RECT 104.195 139.385 104.415 139.535 ;
        RECT 104.195 139.055 104.730 139.385 ;
        RECT 104.900 139.245 105.070 139.580 ;
        RECT 105.995 139.415 106.235 139.935 ;
        RECT 106.450 139.715 106.780 140.105 ;
        RECT 106.950 139.545 107.175 139.925 ;
        RECT 104.195 138.405 104.430 139.055 ;
        RECT 104.900 138.885 105.885 139.245 ;
        RECT 101.395 138.195 102.685 138.365 ;
        RECT 101.395 137.775 101.645 138.195 ;
        RECT 101.875 137.555 102.205 138.025 ;
        RECT 102.435 137.775 102.685 138.195 ;
        RECT 102.865 138.195 103.320 138.365 ;
        RECT 102.865 137.765 103.195 138.195 ;
        RECT 103.755 138.175 104.430 138.405 ;
        RECT 104.600 138.865 105.885 138.885 ;
        RECT 104.600 138.715 105.460 138.865 ;
        RECT 103.755 137.745 103.925 138.175 ;
        RECT 104.095 137.555 104.425 138.005 ;
        RECT 104.600 137.770 104.885 138.715 ;
        RECT 106.060 138.610 106.235 139.415 ;
        RECT 106.435 138.865 106.675 139.515 ;
        RECT 106.845 139.365 107.175 139.545 ;
        RECT 106.845 138.695 107.020 139.365 ;
        RECT 107.375 139.195 107.605 139.815 ;
        RECT 107.785 139.375 108.085 140.105 ;
        RECT 108.265 139.560 113.610 140.105 ;
        RECT 107.190 138.865 107.605 139.195 ;
        RECT 107.785 138.865 108.080 139.195 ;
        RECT 109.850 138.730 110.190 139.560 ;
        RECT 114.245 139.380 114.535 140.105 ;
        RECT 114.905 139.475 115.235 139.835 ;
        RECT 115.855 139.645 116.105 140.105 ;
        RECT 116.275 139.645 116.835 139.935 ;
        RECT 114.905 139.285 116.295 139.475 ;
        RECT 105.060 138.235 105.755 138.545 ;
        RECT 105.065 137.555 105.750 138.025 ;
        RECT 105.930 137.825 106.235 138.610 ;
        RECT 106.435 138.505 107.020 138.695 ;
        RECT 106.435 137.735 106.710 138.505 ;
        RECT 107.190 138.335 108.085 138.665 ;
        RECT 106.880 138.165 108.085 138.335 ;
        RECT 106.880 137.735 107.210 138.165 ;
        RECT 107.380 137.555 107.575 137.995 ;
        RECT 107.755 137.735 108.085 138.165 ;
        RECT 111.670 137.990 112.020 139.240 ;
        RECT 116.125 139.195 116.295 139.285 ;
        RECT 114.720 138.865 115.395 139.115 ;
        RECT 115.615 138.865 115.955 139.115 ;
        RECT 116.125 138.865 116.415 139.195 ;
        RECT 108.265 137.555 113.610 137.990 ;
        RECT 114.245 137.555 114.535 138.720 ;
        RECT 114.720 138.505 114.985 138.865 ;
        RECT 116.125 138.615 116.295 138.865 ;
        RECT 115.355 138.445 116.295 138.615 ;
        RECT 114.905 137.555 115.185 138.225 ;
        RECT 115.355 137.895 115.655 138.445 ;
        RECT 116.585 138.275 116.835 139.645 ;
        RECT 117.005 139.560 122.350 140.105 ;
        RECT 122.525 139.560 127.870 140.105 ;
        RECT 128.045 139.560 133.390 140.105 ;
        RECT 133.565 139.560 138.910 140.105 ;
        RECT 118.590 138.730 118.930 139.560 ;
        RECT 115.855 137.555 116.185 138.275 ;
        RECT 116.375 137.725 116.835 138.275 ;
        RECT 120.410 137.990 120.760 139.240 ;
        RECT 124.110 138.730 124.450 139.560 ;
        RECT 125.930 137.990 126.280 139.240 ;
        RECT 129.630 138.730 129.970 139.560 ;
        RECT 131.450 137.990 131.800 139.240 ;
        RECT 135.150 138.730 135.490 139.560 ;
        RECT 140.005 139.380 140.295 140.105 ;
        RECT 140.465 139.560 145.810 140.105 ;
        RECT 136.970 137.990 137.320 139.240 ;
        RECT 142.050 138.730 142.390 139.560 ;
        RECT 145.985 139.335 148.575 140.105 ;
        RECT 149.205 139.355 150.415 140.105 ;
        RECT 117.005 137.555 122.350 137.990 ;
        RECT 122.525 137.555 127.870 137.990 ;
        RECT 128.045 137.555 133.390 137.990 ;
        RECT 133.565 137.555 138.910 137.990 ;
        RECT 140.005 137.555 140.295 138.720 ;
        RECT 143.870 137.990 144.220 139.240 ;
        RECT 145.985 138.815 147.195 139.335 ;
        RECT 147.365 138.645 148.575 139.165 ;
        RECT 140.465 137.555 145.810 137.990 ;
        RECT 145.985 137.555 148.575 138.645 ;
        RECT 149.205 138.645 149.725 139.185 ;
        RECT 149.895 138.815 150.415 139.355 ;
        RECT 149.205 137.555 150.415 138.645 ;
        RECT 11.120 137.385 150.500 137.555 ;
        RECT 11.205 136.295 12.415 137.385 ;
        RECT 12.585 136.950 17.930 137.385 ;
        RECT 11.205 135.585 11.725 136.125 ;
        RECT 11.895 135.755 12.415 136.295 ;
        RECT 11.205 134.835 12.415 135.585 ;
        RECT 14.170 135.380 14.510 136.210 ;
        RECT 15.990 135.700 16.340 136.950 ;
        RECT 18.565 136.665 19.025 137.215 ;
        RECT 19.215 136.665 19.545 137.385 ;
        RECT 12.585 134.835 17.930 135.380 ;
        RECT 18.565 135.295 18.815 136.665 ;
        RECT 19.745 136.495 20.045 137.045 ;
        RECT 20.215 136.715 20.495 137.385 ;
        RECT 19.105 136.325 20.045 136.495 ;
        RECT 19.105 136.075 19.275 136.325 ;
        RECT 20.415 136.075 20.680 136.435 ;
        RECT 20.865 136.295 23.455 137.385 ;
        RECT 18.985 135.745 19.275 136.075 ;
        RECT 19.445 135.825 19.785 136.075 ;
        RECT 20.005 135.825 20.680 136.075 ;
        RECT 19.105 135.655 19.275 135.745 ;
        RECT 19.105 135.465 20.495 135.655 ;
        RECT 18.565 135.005 19.125 135.295 ;
        RECT 19.295 134.835 19.545 135.295 ;
        RECT 20.165 135.105 20.495 135.465 ;
        RECT 20.865 135.605 22.075 136.125 ;
        RECT 22.245 135.775 23.455 136.295 ;
        RECT 24.085 136.220 24.375 137.385 ;
        RECT 24.545 136.295 26.215 137.385 ;
        RECT 26.385 136.875 26.685 137.385 ;
        RECT 26.855 136.705 27.185 137.215 ;
        RECT 27.355 136.875 27.985 137.385 ;
        RECT 28.565 136.875 28.945 137.045 ;
        RECT 29.115 136.875 29.415 137.385 ;
        RECT 29.605 136.950 34.950 137.385 ;
        RECT 28.775 136.705 28.945 136.875 ;
        RECT 24.545 135.605 25.295 136.125 ;
        RECT 25.465 135.775 26.215 136.295 ;
        RECT 26.385 136.535 28.605 136.705 ;
        RECT 20.865 134.835 23.455 135.605 ;
        RECT 24.085 134.835 24.375 135.560 ;
        RECT 24.545 134.835 26.215 135.605 ;
        RECT 26.385 135.575 26.555 136.535 ;
        RECT 26.725 136.195 28.265 136.365 ;
        RECT 26.725 135.745 26.970 136.195 ;
        RECT 27.230 135.825 27.925 136.025 ;
        RECT 28.095 135.995 28.265 136.195 ;
        RECT 28.435 136.335 28.605 136.535 ;
        RECT 28.775 136.505 29.435 136.705 ;
        RECT 28.435 136.165 29.095 136.335 ;
        RECT 28.095 135.825 28.695 135.995 ;
        RECT 28.925 135.745 29.095 136.165 ;
        RECT 26.385 135.030 26.850 135.575 ;
        RECT 27.355 134.835 27.525 135.655 ;
        RECT 27.695 135.575 28.605 135.655 ;
        RECT 29.265 135.575 29.435 136.505 ;
        RECT 27.695 135.485 28.945 135.575 ;
        RECT 27.695 135.005 28.025 135.485 ;
        RECT 28.435 135.405 28.945 135.485 ;
        RECT 28.195 134.835 28.545 135.225 ;
        RECT 28.715 135.005 28.945 135.405 ;
        RECT 29.115 135.095 29.435 135.575 ;
        RECT 31.190 135.380 31.530 136.210 ;
        RECT 33.010 135.700 33.360 136.950 ;
        RECT 35.125 136.295 36.795 137.385 ;
        RECT 35.125 135.605 35.875 136.125 ;
        RECT 36.045 135.775 36.795 136.295 ;
        RECT 37.425 136.285 37.745 137.215 ;
        RECT 37.925 136.705 38.325 137.215 ;
        RECT 38.495 136.875 38.665 137.385 ;
        RECT 38.835 136.705 39.165 137.215 ;
        RECT 37.925 136.535 39.165 136.705 ;
        RECT 39.335 136.535 39.505 137.385 ;
        RECT 40.095 136.535 40.475 137.215 ;
        RECT 37.425 136.115 38.055 136.285 ;
        RECT 29.605 134.835 34.950 135.380 ;
        RECT 35.125 134.835 36.795 135.605 ;
        RECT 37.425 134.835 37.715 135.670 ;
        RECT 37.885 135.235 38.055 136.115 ;
        RECT 38.830 136.195 40.135 136.365 ;
        RECT 38.225 135.575 38.455 136.075 ;
        RECT 38.830 135.995 39.000 136.195 ;
        RECT 38.625 135.825 39.000 135.995 ;
        RECT 39.170 135.825 39.720 136.025 ;
        RECT 39.890 135.745 40.135 136.195 ;
        RECT 40.305 135.575 40.475 136.535 ;
        RECT 41.585 136.495 41.845 137.205 ;
        RECT 42.015 136.675 42.345 137.385 ;
        RECT 42.515 136.495 42.745 137.205 ;
        RECT 41.585 136.255 42.745 136.495 ;
        RECT 42.925 136.475 43.195 137.205 ;
        RECT 43.375 136.655 43.715 137.385 ;
        RECT 42.925 136.255 43.695 136.475 ;
        RECT 41.575 135.745 41.875 136.075 ;
        RECT 42.055 135.765 42.580 136.075 ;
        RECT 42.760 135.765 43.225 136.075 ;
        RECT 38.225 135.405 40.475 135.575 ;
        RECT 37.885 135.065 38.840 135.235 ;
        RECT 39.255 134.835 39.585 135.225 ;
        RECT 39.755 135.085 39.925 135.405 ;
        RECT 40.095 134.835 40.425 135.225 ;
        RECT 41.585 134.835 41.875 135.565 ;
        RECT 42.055 135.125 42.285 135.765 ;
        RECT 43.405 135.585 43.695 136.255 ;
        RECT 42.465 135.385 43.695 135.585 ;
        RECT 42.465 135.015 42.775 135.385 ;
        RECT 42.955 134.835 43.625 135.205 ;
        RECT 43.885 135.015 44.145 137.205 ;
        RECT 44.325 136.310 44.665 137.385 ;
        RECT 44.850 136.875 46.900 137.165 ;
        RECT 44.835 136.075 45.075 136.670 ;
        RECT 45.270 136.535 46.900 136.705 ;
        RECT 47.070 136.585 47.350 137.385 ;
        RECT 45.270 136.245 45.590 136.535 ;
        RECT 46.730 136.415 46.900 136.535 ;
        RECT 44.325 135.505 44.665 136.075 ;
        RECT 44.835 135.745 45.490 136.075 ;
        RECT 45.760 135.745 46.500 136.365 ;
        RECT 46.730 136.245 47.390 136.415 ;
        RECT 47.560 136.245 47.835 137.215 ;
        RECT 48.015 136.415 48.345 137.200 ;
        RECT 48.015 136.245 48.695 136.415 ;
        RECT 48.875 136.245 49.205 137.385 ;
        RECT 47.220 136.075 47.390 136.245 ;
        RECT 46.670 135.745 47.050 136.075 ;
        RECT 47.220 135.745 47.495 136.075 ;
        RECT 44.325 134.835 44.665 135.335 ;
        RECT 44.835 135.055 45.080 135.745 ;
        RECT 47.220 135.575 47.390 135.745 ;
        RECT 45.805 135.405 47.390 135.575 ;
        RECT 47.665 135.510 47.835 136.245 ;
        RECT 48.005 135.825 48.355 136.075 ;
        RECT 48.525 135.645 48.695 136.245 ;
        RECT 49.845 136.220 50.135 137.385 ;
        RECT 50.765 136.535 51.145 137.215 ;
        RECT 51.735 136.535 51.905 137.385 ;
        RECT 52.075 136.705 52.405 137.215 ;
        RECT 52.575 136.875 52.745 137.385 ;
        RECT 52.915 136.705 53.315 137.215 ;
        RECT 52.075 136.535 53.315 136.705 ;
        RECT 48.865 135.825 49.215 136.075 ;
        RECT 45.275 134.835 45.605 135.335 ;
        RECT 45.805 135.055 45.975 135.405 ;
        RECT 46.150 134.835 46.480 135.235 ;
        RECT 46.650 135.055 46.820 135.405 ;
        RECT 46.990 134.835 47.370 135.235 ;
        RECT 47.560 135.165 47.835 135.510 ;
        RECT 48.025 134.835 48.265 135.645 ;
        RECT 48.435 135.005 48.765 135.645 ;
        RECT 48.935 134.835 49.205 135.645 ;
        RECT 50.765 135.575 50.935 136.535 ;
        RECT 51.105 136.195 52.410 136.365 ;
        RECT 53.495 136.285 53.815 137.215 ;
        RECT 53.985 136.295 56.575 137.385 ;
        RECT 51.105 135.745 51.350 136.195 ;
        RECT 51.520 135.825 52.070 136.025 ;
        RECT 52.240 135.995 52.410 136.195 ;
        RECT 53.185 136.115 53.815 136.285 ;
        RECT 52.240 135.825 52.615 135.995 ;
        RECT 52.785 135.575 53.015 136.075 ;
        RECT 49.845 134.835 50.135 135.560 ;
        RECT 50.765 135.405 53.015 135.575 ;
        RECT 50.815 134.835 51.145 135.225 ;
        RECT 51.315 135.085 51.485 135.405 ;
        RECT 53.185 135.235 53.355 136.115 ;
        RECT 51.655 134.835 51.985 135.225 ;
        RECT 52.400 135.065 53.355 135.235 ;
        RECT 53.525 134.835 53.815 135.670 ;
        RECT 53.985 135.605 55.195 136.125 ;
        RECT 55.365 135.775 56.575 136.295 ;
        RECT 57.205 136.245 57.485 137.385 ;
        RECT 57.655 136.235 57.985 137.215 ;
        RECT 58.155 136.245 58.415 137.385 ;
        RECT 58.585 136.245 58.855 137.215 ;
        RECT 59.065 136.585 59.345 137.385 ;
        RECT 59.525 136.835 60.720 137.165 ;
        RECT 59.850 136.415 60.270 136.665 ;
        RECT 59.025 136.245 60.270 136.415 ;
        RECT 57.215 135.805 57.550 136.075 ;
        RECT 57.720 135.685 57.890 136.235 ;
        RECT 58.585 136.195 58.815 136.245 ;
        RECT 58.060 135.825 58.395 136.075 ;
        RECT 57.720 135.635 57.895 135.685 ;
        RECT 53.985 134.835 56.575 135.605 ;
        RECT 57.205 134.835 57.515 135.635 ;
        RECT 57.720 135.005 58.415 135.635 ;
        RECT 58.585 135.510 58.755 136.195 ;
        RECT 59.025 136.075 59.195 136.245 ;
        RECT 60.495 136.075 60.665 136.635 ;
        RECT 60.915 136.245 61.170 137.385 ;
        RECT 61.345 136.515 61.620 137.215 ;
        RECT 61.790 136.840 62.045 137.385 ;
        RECT 62.215 136.875 62.695 137.215 ;
        RECT 62.870 136.830 63.475 137.385 ;
        RECT 62.860 136.730 63.475 136.830 ;
        RECT 62.860 136.705 63.045 136.730 ;
        RECT 58.965 135.745 59.195 136.075 ;
        RECT 59.925 135.745 60.665 136.075 ;
        RECT 60.835 135.825 61.170 136.075 ;
        RECT 59.025 135.575 59.195 135.745 ;
        RECT 60.415 135.655 60.665 135.745 ;
        RECT 58.585 135.165 58.855 135.510 ;
        RECT 59.025 135.405 59.765 135.575 ;
        RECT 60.415 135.485 61.150 135.655 ;
        RECT 59.045 134.835 59.425 135.235 ;
        RECT 59.595 135.055 59.765 135.405 ;
        RECT 59.935 134.835 60.670 135.315 ;
        RECT 60.840 135.015 61.150 135.485 ;
        RECT 61.345 135.485 61.515 136.515 ;
        RECT 61.790 136.385 62.545 136.635 ;
        RECT 62.715 136.460 63.045 136.705 ;
        RECT 64.655 136.715 64.825 137.215 ;
        RECT 64.995 136.885 65.325 137.385 ;
        RECT 61.790 136.350 62.560 136.385 ;
        RECT 61.790 136.340 62.575 136.350 ;
        RECT 61.685 136.325 62.580 136.340 ;
        RECT 61.685 136.310 62.600 136.325 ;
        RECT 61.685 136.300 62.620 136.310 ;
        RECT 61.685 136.290 62.645 136.300 ;
        RECT 61.685 136.260 62.715 136.290 ;
        RECT 61.685 136.230 62.735 136.260 ;
        RECT 61.685 136.200 62.755 136.230 ;
        RECT 61.685 136.175 62.785 136.200 ;
        RECT 61.685 136.140 62.820 136.175 ;
        RECT 61.685 136.135 62.850 136.140 ;
        RECT 61.685 135.740 61.915 136.135 ;
        RECT 62.460 136.130 62.850 136.135 ;
        RECT 62.485 136.120 62.850 136.130 ;
        RECT 62.500 136.115 62.850 136.120 ;
        RECT 62.515 136.110 62.850 136.115 ;
        RECT 63.215 136.110 63.475 136.560 ;
        RECT 64.655 136.545 65.320 136.715 ;
        RECT 62.515 136.105 63.475 136.110 ;
        RECT 62.525 136.095 63.475 136.105 ;
        RECT 62.535 136.090 63.475 136.095 ;
        RECT 62.545 136.080 63.475 136.090 ;
        RECT 62.550 136.070 63.475 136.080 ;
        RECT 62.555 136.065 63.475 136.070 ;
        RECT 62.565 136.050 63.475 136.065 ;
        RECT 62.570 136.035 63.475 136.050 ;
        RECT 62.580 136.010 63.475 136.035 ;
        RECT 62.085 135.540 62.415 135.965 ;
        RECT 61.345 135.005 61.605 135.485 ;
        RECT 61.775 134.835 62.025 135.375 ;
        RECT 62.195 135.055 62.415 135.540 ;
        RECT 62.585 135.940 63.475 136.010 ;
        RECT 62.585 135.215 62.755 135.940 ;
        RECT 62.925 135.385 63.475 135.770 ;
        RECT 64.570 135.725 64.920 136.375 ;
        RECT 65.090 135.555 65.320 136.545 ;
        RECT 64.655 135.385 65.320 135.555 ;
        RECT 62.585 135.045 63.475 135.215 ;
        RECT 64.655 135.095 64.825 135.385 ;
        RECT 64.995 134.835 65.325 135.215 ;
        RECT 65.495 135.095 65.680 137.215 ;
        RECT 65.920 136.925 66.185 137.385 ;
        RECT 66.355 136.790 66.605 137.215 ;
        RECT 66.815 136.940 67.920 137.110 ;
        RECT 66.300 136.660 66.605 136.790 ;
        RECT 65.850 135.465 66.130 136.415 ;
        RECT 66.300 135.555 66.470 136.660 ;
        RECT 66.640 135.875 66.880 136.470 ;
        RECT 67.050 136.405 67.580 136.770 ;
        RECT 67.050 135.705 67.220 136.405 ;
        RECT 67.750 136.325 67.920 136.940 ;
        RECT 68.090 136.585 68.260 137.385 ;
        RECT 68.430 136.885 68.680 137.215 ;
        RECT 68.905 136.915 69.790 137.085 ;
        RECT 67.750 136.235 68.260 136.325 ;
        RECT 66.300 135.425 66.525 135.555 ;
        RECT 66.695 135.485 67.220 135.705 ;
        RECT 67.390 136.065 68.260 136.235 ;
        RECT 65.935 134.835 66.185 135.295 ;
        RECT 66.355 135.285 66.525 135.425 ;
        RECT 67.390 135.285 67.560 136.065 ;
        RECT 68.090 135.995 68.260 136.065 ;
        RECT 67.770 135.815 67.970 135.845 ;
        RECT 68.430 135.815 68.600 136.885 ;
        RECT 68.770 135.995 68.960 136.715 ;
        RECT 67.770 135.515 68.600 135.815 ;
        RECT 69.130 135.785 69.450 136.745 ;
        RECT 66.355 135.115 66.690 135.285 ;
        RECT 66.885 135.115 67.560 135.285 ;
        RECT 67.880 134.835 68.250 135.335 ;
        RECT 68.430 135.285 68.600 135.515 ;
        RECT 68.985 135.455 69.450 135.785 ;
        RECT 69.620 136.075 69.790 136.915 ;
        RECT 69.970 136.885 70.285 137.385 ;
        RECT 70.515 136.655 70.855 137.215 ;
        RECT 69.960 136.280 70.855 136.655 ;
        RECT 71.025 136.375 71.195 137.385 ;
        RECT 70.665 136.075 70.855 136.280 ;
        RECT 71.365 136.325 71.695 137.170 ;
        RECT 71.865 136.470 72.035 137.385 ;
        RECT 72.385 136.515 72.660 137.215 ;
        RECT 72.830 136.840 73.085 137.385 ;
        RECT 73.255 136.875 73.735 137.215 ;
        RECT 73.910 136.830 74.515 137.385 ;
        RECT 73.900 136.730 74.515 136.830 ;
        RECT 73.900 136.705 74.085 136.730 ;
        RECT 71.365 136.245 71.755 136.325 ;
        RECT 71.540 136.195 71.755 136.245 ;
        RECT 69.620 135.745 70.495 136.075 ;
        RECT 70.665 135.745 71.415 136.075 ;
        RECT 69.620 135.285 69.790 135.745 ;
        RECT 70.665 135.575 70.865 135.745 ;
        RECT 71.585 135.615 71.755 136.195 ;
        RECT 71.530 135.575 71.755 135.615 ;
        RECT 68.430 135.115 68.835 135.285 ;
        RECT 69.005 135.115 69.790 135.285 ;
        RECT 70.065 134.835 70.275 135.365 ;
        RECT 70.535 135.050 70.865 135.575 ;
        RECT 71.375 135.490 71.755 135.575 ;
        RECT 71.035 134.835 71.205 135.445 ;
        RECT 71.375 135.055 71.705 135.490 ;
        RECT 72.385 135.485 72.555 136.515 ;
        RECT 72.830 136.385 73.585 136.635 ;
        RECT 73.755 136.460 74.085 136.705 ;
        RECT 72.830 136.350 73.600 136.385 ;
        RECT 72.830 136.340 73.615 136.350 ;
        RECT 72.725 136.325 73.620 136.340 ;
        RECT 72.725 136.310 73.640 136.325 ;
        RECT 72.725 136.300 73.660 136.310 ;
        RECT 72.725 136.290 73.685 136.300 ;
        RECT 72.725 136.260 73.755 136.290 ;
        RECT 72.725 136.230 73.775 136.260 ;
        RECT 72.725 136.200 73.795 136.230 ;
        RECT 72.725 136.175 73.825 136.200 ;
        RECT 72.725 136.140 73.860 136.175 ;
        RECT 72.725 136.135 73.890 136.140 ;
        RECT 72.725 135.740 72.955 136.135 ;
        RECT 73.500 136.130 73.890 136.135 ;
        RECT 73.525 136.120 73.890 136.130 ;
        RECT 73.540 136.115 73.890 136.120 ;
        RECT 73.555 136.110 73.890 136.115 ;
        RECT 74.255 136.110 74.515 136.560 ;
        RECT 75.605 136.220 75.895 137.385 ;
        RECT 76.065 136.515 76.340 137.215 ;
        RECT 76.510 136.840 76.765 137.385 ;
        RECT 76.935 136.875 77.415 137.215 ;
        RECT 77.590 136.830 78.195 137.385 ;
        RECT 77.580 136.730 78.195 136.830 ;
        RECT 77.580 136.705 77.765 136.730 ;
        RECT 73.555 136.105 74.515 136.110 ;
        RECT 73.565 136.095 74.515 136.105 ;
        RECT 73.575 136.090 74.515 136.095 ;
        RECT 73.585 136.080 74.515 136.090 ;
        RECT 73.590 136.070 74.515 136.080 ;
        RECT 73.595 136.065 74.515 136.070 ;
        RECT 73.605 136.050 74.515 136.065 ;
        RECT 73.610 136.035 74.515 136.050 ;
        RECT 73.620 136.010 74.515 136.035 ;
        RECT 73.125 135.540 73.455 135.965 ;
        RECT 71.875 134.835 72.045 135.350 ;
        RECT 72.385 135.005 72.645 135.485 ;
        RECT 72.815 134.835 73.065 135.375 ;
        RECT 73.235 135.055 73.455 135.540 ;
        RECT 73.625 135.940 74.515 136.010 ;
        RECT 73.625 135.215 73.795 135.940 ;
        RECT 73.965 135.385 74.515 135.770 ;
        RECT 73.625 135.045 74.515 135.215 ;
        RECT 75.605 134.835 75.895 135.560 ;
        RECT 76.065 135.485 76.235 136.515 ;
        RECT 76.510 136.385 77.265 136.635 ;
        RECT 77.435 136.460 77.765 136.705 ;
        RECT 76.510 136.350 77.280 136.385 ;
        RECT 76.510 136.340 77.295 136.350 ;
        RECT 76.405 136.325 77.300 136.340 ;
        RECT 76.405 136.310 77.320 136.325 ;
        RECT 76.405 136.300 77.340 136.310 ;
        RECT 76.405 136.290 77.365 136.300 ;
        RECT 76.405 136.260 77.435 136.290 ;
        RECT 76.405 136.230 77.455 136.260 ;
        RECT 76.405 136.200 77.475 136.230 ;
        RECT 76.405 136.175 77.505 136.200 ;
        RECT 76.405 136.140 77.540 136.175 ;
        RECT 76.405 136.135 77.570 136.140 ;
        RECT 76.405 135.740 76.635 136.135 ;
        RECT 77.180 136.130 77.570 136.135 ;
        RECT 77.205 136.120 77.570 136.130 ;
        RECT 77.220 136.115 77.570 136.120 ;
        RECT 77.235 136.110 77.570 136.115 ;
        RECT 77.935 136.110 78.195 136.560 ;
        RECT 78.365 136.295 81.875 137.385 ;
        RECT 77.235 136.105 78.195 136.110 ;
        RECT 77.245 136.095 78.195 136.105 ;
        RECT 77.255 136.090 78.195 136.095 ;
        RECT 77.265 136.080 78.195 136.090 ;
        RECT 77.270 136.070 78.195 136.080 ;
        RECT 77.275 136.065 78.195 136.070 ;
        RECT 77.285 136.050 78.195 136.065 ;
        RECT 77.290 136.035 78.195 136.050 ;
        RECT 77.300 136.010 78.195 136.035 ;
        RECT 76.805 135.540 77.135 135.965 ;
        RECT 76.065 135.005 76.325 135.485 ;
        RECT 76.495 134.835 76.745 135.375 ;
        RECT 76.915 135.055 77.135 135.540 ;
        RECT 77.305 135.940 78.195 136.010 ;
        RECT 77.305 135.215 77.475 135.940 ;
        RECT 77.645 135.385 78.195 135.770 ;
        RECT 78.365 135.605 80.015 136.125 ;
        RECT 80.185 135.775 81.875 136.295 ;
        RECT 82.055 136.775 82.385 137.205 ;
        RECT 82.565 136.945 82.760 137.385 ;
        RECT 82.930 136.775 83.260 137.205 ;
        RECT 82.055 136.605 83.260 136.775 ;
        RECT 82.055 136.275 82.950 136.605 ;
        RECT 83.430 136.435 83.705 137.205 ;
        RECT 83.120 136.245 83.705 136.435 ;
        RECT 83.885 136.245 84.145 137.385 ;
        RECT 82.060 135.745 82.355 136.075 ;
        RECT 82.535 135.745 82.950 136.075 ;
        RECT 77.305 135.045 78.195 135.215 ;
        RECT 78.365 134.835 81.875 135.605 ;
        RECT 82.055 134.835 82.355 135.565 ;
        RECT 82.535 135.125 82.765 135.745 ;
        RECT 83.120 135.575 83.295 136.245 ;
        RECT 84.315 136.235 84.645 137.215 ;
        RECT 84.815 136.245 85.095 137.385 ;
        RECT 85.265 136.295 86.935 137.385 ;
        RECT 82.965 135.395 83.295 135.575 ;
        RECT 83.465 135.425 83.705 136.075 ;
        RECT 83.905 135.825 84.240 136.075 ;
        RECT 84.410 135.635 84.580 136.235 ;
        RECT 84.750 135.805 85.085 136.075 ;
        RECT 82.965 135.015 83.190 135.395 ;
        RECT 83.360 134.835 83.690 135.225 ;
        RECT 83.885 135.005 84.580 135.635 ;
        RECT 84.785 134.835 85.095 135.635 ;
        RECT 85.265 135.605 86.015 136.125 ;
        RECT 86.185 135.775 86.935 136.295 ;
        RECT 87.565 136.535 87.945 137.215 ;
        RECT 88.535 136.535 88.705 137.385 ;
        RECT 88.875 136.705 89.205 137.215 ;
        RECT 89.375 136.875 89.545 137.385 ;
        RECT 89.715 136.705 90.115 137.215 ;
        RECT 88.875 136.535 90.115 136.705 ;
        RECT 85.265 134.835 86.935 135.605 ;
        RECT 87.565 135.575 87.735 136.535 ;
        RECT 87.905 136.195 89.210 136.365 ;
        RECT 90.295 136.285 90.615 137.215 ;
        RECT 90.785 136.295 91.995 137.385 ;
        RECT 87.905 135.745 88.150 136.195 ;
        RECT 88.320 135.825 88.870 136.025 ;
        RECT 89.040 135.995 89.210 136.195 ;
        RECT 89.985 136.115 90.615 136.285 ;
        RECT 89.040 135.825 89.415 135.995 ;
        RECT 89.585 135.575 89.815 136.075 ;
        RECT 87.565 135.405 89.815 135.575 ;
        RECT 87.615 134.835 87.945 135.225 ;
        RECT 88.115 135.085 88.285 135.405 ;
        RECT 89.985 135.235 90.155 136.115 ;
        RECT 88.455 134.835 88.785 135.225 ;
        RECT 89.200 135.065 90.155 135.235 ;
        RECT 90.325 134.835 90.615 135.670 ;
        RECT 90.785 135.585 91.305 136.125 ;
        RECT 91.475 135.755 91.995 136.295 ;
        RECT 92.170 136.995 92.505 137.215 ;
        RECT 93.510 137.005 93.865 137.385 ;
        RECT 92.170 136.375 92.425 136.995 ;
        RECT 92.675 136.835 92.905 136.875 ;
        RECT 94.035 136.835 94.285 137.215 ;
        RECT 92.675 136.635 94.285 136.835 ;
        RECT 92.675 136.545 92.860 136.635 ;
        RECT 93.450 136.625 94.285 136.635 ;
        RECT 94.535 136.605 94.785 137.385 ;
        RECT 94.955 136.535 95.215 137.215 ;
        RECT 95.585 136.715 95.865 137.385 ;
        RECT 93.015 136.435 93.345 136.465 ;
        RECT 93.015 136.375 94.815 136.435 ;
        RECT 92.170 136.265 94.875 136.375 ;
        RECT 92.170 136.205 93.345 136.265 ;
        RECT 94.675 136.230 94.875 136.265 ;
        RECT 92.165 135.825 92.655 136.025 ;
        RECT 92.845 135.825 93.320 136.035 ;
        RECT 90.785 134.835 91.995 135.585 ;
        RECT 92.170 134.835 92.625 135.600 ;
        RECT 93.100 135.425 93.320 135.825 ;
        RECT 93.565 135.825 93.895 136.035 ;
        RECT 93.565 135.425 93.775 135.825 ;
        RECT 94.065 135.790 94.475 136.095 ;
        RECT 94.705 135.655 94.875 136.230 ;
        RECT 94.605 135.535 94.875 135.655 ;
        RECT 94.030 135.490 94.875 135.535 ;
        RECT 94.030 135.365 94.785 135.490 ;
        RECT 94.030 135.215 94.200 135.365 ;
        RECT 95.045 135.335 95.215 136.535 ;
        RECT 96.035 136.495 96.335 137.045 ;
        RECT 96.535 136.665 96.865 137.385 ;
        RECT 97.055 136.665 97.515 137.215 ;
        RECT 95.400 136.075 95.665 136.435 ;
        RECT 96.035 136.325 96.975 136.495 ;
        RECT 96.805 136.075 96.975 136.325 ;
        RECT 95.400 135.825 96.075 136.075 ;
        RECT 96.295 135.825 96.635 136.075 ;
        RECT 96.805 135.745 97.095 136.075 ;
        RECT 96.805 135.655 96.975 135.745 ;
        RECT 92.900 135.005 94.200 135.215 ;
        RECT 94.455 134.835 94.785 135.195 ;
        RECT 94.955 135.005 95.215 135.335 ;
        RECT 95.585 135.465 96.975 135.655 ;
        RECT 95.585 135.105 95.915 135.465 ;
        RECT 97.265 135.295 97.515 136.665 ;
        RECT 96.535 134.835 96.785 135.295 ;
        RECT 96.955 135.005 97.515 135.295 ;
        RECT 97.685 136.310 97.955 137.215 ;
        RECT 98.125 136.625 98.455 137.385 ;
        RECT 98.635 136.455 98.805 137.215 ;
        RECT 97.685 135.510 97.855 136.310 ;
        RECT 98.140 136.285 98.805 136.455 ;
        RECT 99.065 136.295 100.735 137.385 ;
        RECT 98.140 136.140 98.310 136.285 ;
        RECT 98.025 135.810 98.310 136.140 ;
        RECT 98.140 135.555 98.310 135.810 ;
        RECT 98.545 135.735 98.875 136.105 ;
        RECT 99.065 135.605 99.815 136.125 ;
        RECT 99.985 135.775 100.735 136.295 ;
        RECT 101.365 136.220 101.655 137.385 ;
        RECT 101.825 136.950 107.170 137.385 ;
        RECT 107.345 136.950 112.690 137.385 ;
        RECT 112.865 136.950 118.210 137.385 ;
        RECT 118.385 136.950 123.730 137.385 ;
        RECT 97.685 135.005 97.945 135.510 ;
        RECT 98.140 135.385 98.805 135.555 ;
        RECT 98.125 134.835 98.455 135.215 ;
        RECT 98.635 135.005 98.805 135.385 ;
        RECT 99.065 134.835 100.735 135.605 ;
        RECT 101.365 134.835 101.655 135.560 ;
        RECT 103.410 135.380 103.750 136.210 ;
        RECT 105.230 135.700 105.580 136.950 ;
        RECT 108.930 135.380 109.270 136.210 ;
        RECT 110.750 135.700 111.100 136.950 ;
        RECT 114.450 135.380 114.790 136.210 ;
        RECT 116.270 135.700 116.620 136.950 ;
        RECT 119.970 135.380 120.310 136.210 ;
        RECT 121.790 135.700 122.140 136.950 ;
        RECT 123.905 136.295 126.495 137.385 ;
        RECT 123.905 135.605 125.115 136.125 ;
        RECT 125.285 135.775 126.495 136.295 ;
        RECT 127.125 136.220 127.415 137.385 ;
        RECT 127.585 136.950 132.930 137.385 ;
        RECT 133.105 136.950 138.450 137.385 ;
        RECT 138.625 136.950 143.970 137.385 ;
        RECT 101.825 134.835 107.170 135.380 ;
        RECT 107.345 134.835 112.690 135.380 ;
        RECT 112.865 134.835 118.210 135.380 ;
        RECT 118.385 134.835 123.730 135.380 ;
        RECT 123.905 134.835 126.495 135.605 ;
        RECT 127.125 134.835 127.415 135.560 ;
        RECT 129.170 135.380 129.510 136.210 ;
        RECT 130.990 135.700 131.340 136.950 ;
        RECT 134.690 135.380 135.030 136.210 ;
        RECT 136.510 135.700 136.860 136.950 ;
        RECT 140.210 135.380 140.550 136.210 ;
        RECT 142.030 135.700 142.380 136.950 ;
        RECT 144.145 136.295 147.655 137.385 ;
        RECT 147.825 136.295 149.035 137.385 ;
        RECT 144.145 135.605 145.795 136.125 ;
        RECT 145.965 135.775 147.655 136.295 ;
        RECT 127.585 134.835 132.930 135.380 ;
        RECT 133.105 134.835 138.450 135.380 ;
        RECT 138.625 134.835 143.970 135.380 ;
        RECT 144.145 134.835 147.655 135.605 ;
        RECT 147.825 135.585 148.345 136.125 ;
        RECT 148.515 135.755 149.035 136.295 ;
        RECT 149.205 136.295 150.415 137.385 ;
        RECT 149.205 135.755 149.725 136.295 ;
        RECT 149.895 135.585 150.415 136.125 ;
        RECT 147.825 134.835 149.035 135.585 ;
        RECT 149.205 134.835 150.415 135.585 ;
        RECT 11.120 134.665 150.500 134.835 ;
        RECT 11.205 133.915 12.415 134.665 ;
        RECT 12.585 134.120 17.930 134.665 ;
        RECT 18.105 134.120 23.450 134.665 ;
        RECT 23.625 134.120 28.970 134.665 ;
        RECT 11.205 133.375 11.725 133.915 ;
        RECT 11.895 133.205 12.415 133.745 ;
        RECT 14.170 133.290 14.510 134.120 ;
        RECT 11.205 132.115 12.415 133.205 ;
        RECT 15.990 132.550 16.340 133.800 ;
        RECT 19.690 133.290 20.030 134.120 ;
        RECT 21.510 132.550 21.860 133.800 ;
        RECT 25.210 133.290 25.550 134.120 ;
        RECT 29.145 133.895 30.815 134.665 ;
        RECT 27.030 132.550 27.380 133.800 ;
        RECT 29.145 133.375 29.895 133.895 ;
        RECT 31.505 133.845 31.715 134.665 ;
        RECT 31.885 133.865 32.215 134.495 ;
        RECT 30.065 133.205 30.815 133.725 ;
        RECT 31.885 133.265 32.135 133.865 ;
        RECT 32.385 133.845 32.615 134.665 ;
        RECT 32.825 133.895 35.415 134.665 ;
        RECT 32.305 133.425 32.635 133.675 ;
        RECT 32.825 133.375 34.035 133.895 ;
        RECT 35.585 133.865 36.280 134.495 ;
        RECT 36.485 133.865 36.795 134.665 ;
        RECT 36.965 133.940 37.255 134.665 ;
        RECT 37.425 133.865 37.765 134.495 ;
        RECT 37.935 133.865 38.185 134.665 ;
        RECT 38.375 134.015 38.705 134.495 ;
        RECT 38.875 134.205 39.100 134.665 ;
        RECT 39.270 134.015 39.600 134.495 ;
        RECT 12.585 132.115 17.930 132.550 ;
        RECT 18.105 132.115 23.450 132.550 ;
        RECT 23.625 132.115 28.970 132.550 ;
        RECT 29.145 132.115 30.815 133.205 ;
        RECT 31.505 132.115 31.715 133.255 ;
        RECT 31.885 132.285 32.215 133.265 ;
        RECT 32.385 132.115 32.615 133.255 ;
        RECT 34.205 133.205 35.415 133.725 ;
        RECT 35.605 133.425 35.940 133.675 ;
        RECT 36.110 133.265 36.280 133.865 ;
        RECT 36.450 133.425 36.785 133.695 ;
        RECT 32.825 132.115 35.415 133.205 ;
        RECT 35.585 132.115 35.845 133.255 ;
        RECT 36.015 132.285 36.345 133.265 ;
        RECT 36.515 132.115 36.795 133.255 ;
        RECT 36.965 132.115 37.255 133.280 ;
        RECT 37.425 133.255 37.600 133.865 ;
        RECT 38.375 133.845 39.600 134.015 ;
        RECT 40.230 133.885 40.730 134.495 ;
        RECT 37.770 133.505 38.465 133.675 ;
        RECT 38.295 133.255 38.465 133.505 ;
        RECT 38.640 133.475 39.060 133.675 ;
        RECT 39.230 133.475 39.560 133.675 ;
        RECT 39.730 133.475 40.060 133.675 ;
        RECT 40.230 133.255 40.400 133.885 ;
        RECT 41.575 133.855 41.845 134.665 ;
        RECT 42.015 133.855 42.345 134.495 ;
        RECT 42.515 133.855 42.755 134.665 ;
        RECT 40.585 133.425 40.935 133.675 ;
        RECT 41.565 133.425 41.915 133.675 ;
        RECT 42.085 133.255 42.255 133.855 ;
        RECT 42.945 133.830 43.235 134.665 ;
        RECT 43.405 134.265 44.360 134.435 ;
        RECT 44.775 134.275 45.105 134.665 ;
        RECT 42.425 133.425 42.775 133.675 ;
        RECT 43.405 133.385 43.575 134.265 ;
        RECT 45.275 134.095 45.445 134.415 ;
        RECT 45.615 134.275 45.945 134.665 ;
        RECT 43.745 133.925 45.995 134.095 ;
        RECT 46.185 133.935 46.475 134.665 ;
        RECT 43.745 133.425 43.975 133.925 ;
        RECT 44.145 133.505 44.520 133.675 ;
        RECT 37.425 132.285 37.765 133.255 ;
        RECT 37.935 132.115 38.105 133.255 ;
        RECT 38.295 133.085 40.730 133.255 ;
        RECT 38.375 132.115 38.625 132.915 ;
        RECT 39.270 132.285 39.600 133.085 ;
        RECT 39.900 132.115 40.230 132.915 ;
        RECT 40.400 132.285 40.730 133.085 ;
        RECT 41.575 132.115 41.905 133.255 ;
        RECT 42.085 133.085 42.765 133.255 ;
        RECT 42.435 132.300 42.765 133.085 ;
        RECT 42.945 133.215 43.575 133.385 ;
        RECT 44.350 133.305 44.520 133.505 ;
        RECT 44.690 133.475 45.240 133.675 ;
        RECT 45.410 133.305 45.655 133.755 ;
        RECT 42.945 132.285 43.265 133.215 ;
        RECT 44.350 133.135 45.655 133.305 ;
        RECT 45.825 132.965 45.995 133.925 ;
        RECT 46.175 133.425 46.475 133.755 ;
        RECT 46.655 133.735 46.885 134.375 ;
        RECT 47.065 134.115 47.375 134.485 ;
        RECT 47.555 134.295 48.225 134.665 ;
        RECT 47.065 133.915 48.295 134.115 ;
        RECT 46.655 133.425 47.180 133.735 ;
        RECT 47.360 133.425 47.825 133.735 ;
        RECT 48.005 133.245 48.295 133.915 ;
        RECT 43.445 132.795 44.685 132.965 ;
        RECT 43.445 132.285 43.845 132.795 ;
        RECT 44.015 132.115 44.185 132.625 ;
        RECT 44.355 132.285 44.685 132.795 ;
        RECT 44.855 132.115 45.025 132.965 ;
        RECT 45.615 132.285 45.995 132.965 ;
        RECT 46.185 133.005 47.345 133.245 ;
        RECT 46.185 132.295 46.445 133.005 ;
        RECT 46.615 132.115 46.945 132.825 ;
        RECT 47.115 132.295 47.345 133.005 ;
        RECT 47.525 133.025 48.295 133.245 ;
        RECT 47.525 132.295 47.795 133.025 ;
        RECT 47.975 132.115 48.315 132.845 ;
        RECT 48.485 132.295 48.745 134.485 ;
        RECT 48.925 133.895 51.515 134.665 ;
        RECT 52.170 134.015 52.480 134.485 ;
        RECT 52.650 134.185 53.385 134.665 ;
        RECT 53.555 134.095 53.725 134.445 ;
        RECT 53.895 134.265 54.275 134.665 ;
        RECT 48.925 133.375 50.135 133.895 ;
        RECT 52.170 133.845 52.905 134.015 ;
        RECT 53.555 133.925 54.295 134.095 ;
        RECT 54.465 133.990 54.735 134.335 ;
        RECT 54.905 134.120 60.250 134.665 ;
        RECT 52.655 133.755 52.905 133.845 ;
        RECT 54.125 133.755 54.295 133.925 ;
        RECT 50.305 133.205 51.515 133.725 ;
        RECT 52.150 133.425 52.485 133.675 ;
        RECT 52.655 133.425 53.395 133.755 ;
        RECT 54.125 133.425 54.355 133.755 ;
        RECT 48.925 132.115 51.515 133.205 ;
        RECT 52.150 132.115 52.405 133.255 ;
        RECT 52.655 132.865 52.825 133.425 ;
        RECT 54.125 133.255 54.295 133.425 ;
        RECT 54.565 133.255 54.735 133.990 ;
        RECT 56.490 133.290 56.830 134.120 ;
        RECT 60.425 133.895 62.095 134.665 ;
        RECT 62.725 133.940 63.015 134.665 ;
        RECT 63.185 133.895 64.855 134.665 ;
        RECT 53.050 133.085 54.295 133.255 ;
        RECT 53.050 132.835 53.470 133.085 ;
        RECT 52.600 132.335 53.795 132.665 ;
        RECT 53.975 132.115 54.255 132.915 ;
        RECT 54.465 132.285 54.735 133.255 ;
        RECT 58.310 132.550 58.660 133.800 ;
        RECT 60.425 133.375 61.175 133.895 ;
        RECT 61.345 133.205 62.095 133.725 ;
        RECT 63.185 133.375 63.935 133.895 ;
        RECT 65.485 133.865 66.180 134.495 ;
        RECT 66.385 133.865 66.695 134.665 ;
        RECT 54.905 132.115 60.250 132.550 ;
        RECT 60.425 132.115 62.095 133.205 ;
        RECT 62.725 132.115 63.015 133.280 ;
        RECT 64.105 133.205 64.855 133.725 ;
        RECT 65.505 133.425 65.840 133.675 ;
        RECT 66.010 133.265 66.180 133.865 ;
        RECT 67.785 133.720 68.125 134.495 ;
        RECT 68.295 134.205 68.465 134.665 ;
        RECT 68.705 134.230 69.065 134.495 ;
        RECT 68.705 134.225 69.060 134.230 ;
        RECT 68.705 134.215 69.055 134.225 ;
        RECT 68.705 134.210 69.050 134.215 ;
        RECT 68.705 134.200 69.045 134.210 ;
        RECT 69.695 134.205 69.865 134.665 ;
        RECT 68.705 134.195 69.040 134.200 ;
        RECT 68.705 134.185 69.030 134.195 ;
        RECT 68.705 134.175 69.020 134.185 ;
        RECT 68.705 134.035 69.005 134.175 ;
        RECT 68.295 133.845 69.005 134.035 ;
        RECT 69.195 134.035 69.525 134.115 ;
        RECT 70.035 134.035 70.375 134.495 ;
        RECT 70.545 134.120 75.890 134.665 ;
        RECT 76.065 134.120 81.410 134.665 ;
        RECT 81.585 134.120 86.930 134.665 ;
        RECT 69.195 133.845 70.375 134.035 ;
        RECT 66.350 133.425 66.685 133.695 ;
        RECT 63.185 132.115 64.855 133.205 ;
        RECT 65.485 132.115 65.745 133.255 ;
        RECT 65.915 132.285 66.245 133.265 ;
        RECT 66.415 132.115 66.695 133.255 ;
        RECT 67.785 132.285 68.065 133.720 ;
        RECT 68.295 133.275 68.580 133.845 ;
        RECT 68.765 133.445 69.235 133.675 ;
        RECT 69.405 133.655 69.735 133.675 ;
        RECT 69.405 133.475 69.855 133.655 ;
        RECT 70.045 133.475 70.375 133.675 ;
        RECT 68.295 133.060 69.445 133.275 ;
        RECT 68.235 132.115 68.945 132.890 ;
        RECT 69.115 132.285 69.445 133.060 ;
        RECT 69.640 132.360 69.855 133.475 ;
        RECT 70.145 133.135 70.375 133.475 ;
        RECT 72.130 133.290 72.470 134.120 ;
        RECT 70.035 132.115 70.365 132.835 ;
        RECT 73.950 132.550 74.300 133.800 ;
        RECT 77.650 133.290 77.990 134.120 ;
        RECT 79.470 132.550 79.820 133.800 ;
        RECT 83.170 133.290 83.510 134.120 ;
        RECT 87.105 133.915 88.315 134.665 ;
        RECT 88.485 133.940 88.775 134.665 ;
        RECT 88.945 134.120 94.290 134.665 ;
        RECT 94.465 134.120 99.810 134.665 ;
        RECT 84.990 132.550 85.340 133.800 ;
        RECT 87.105 133.375 87.625 133.915 ;
        RECT 87.795 133.205 88.315 133.745 ;
        RECT 90.530 133.290 90.870 134.120 ;
        RECT 70.545 132.115 75.890 132.550 ;
        RECT 76.065 132.115 81.410 132.550 ;
        RECT 81.585 132.115 86.930 132.550 ;
        RECT 87.105 132.115 88.315 133.205 ;
        RECT 88.485 132.115 88.775 133.280 ;
        RECT 92.350 132.550 92.700 133.800 ;
        RECT 96.050 133.290 96.390 134.120 ;
        RECT 99.985 133.915 101.195 134.665 ;
        RECT 101.365 133.925 101.830 134.470 ;
        RECT 97.870 132.550 98.220 133.800 ;
        RECT 99.985 133.375 100.505 133.915 ;
        RECT 100.675 133.205 101.195 133.745 ;
        RECT 88.945 132.115 94.290 132.550 ;
        RECT 94.465 132.115 99.810 132.550 ;
        RECT 99.985 132.115 101.195 133.205 ;
        RECT 101.365 132.965 101.535 133.925 ;
        RECT 102.335 133.845 102.505 134.665 ;
        RECT 102.675 134.015 103.005 134.495 ;
        RECT 103.175 134.275 103.525 134.665 ;
        RECT 103.695 134.095 103.925 134.495 ;
        RECT 103.415 134.015 103.925 134.095 ;
        RECT 102.675 133.925 103.925 134.015 ;
        RECT 104.095 133.925 104.415 134.405 ;
        RECT 102.675 133.845 103.585 133.925 ;
        RECT 101.705 133.305 101.950 133.755 ;
        RECT 102.210 133.475 102.905 133.675 ;
        RECT 103.075 133.505 103.675 133.675 ;
        RECT 103.075 133.305 103.245 133.505 ;
        RECT 103.905 133.335 104.075 133.755 ;
        RECT 101.705 133.135 103.245 133.305 ;
        RECT 103.415 133.165 104.075 133.335 ;
        RECT 103.415 132.965 103.585 133.165 ;
        RECT 104.245 132.995 104.415 133.925 ;
        RECT 104.625 133.845 104.855 134.665 ;
        RECT 105.025 133.865 105.355 134.495 ;
        RECT 104.605 133.425 104.935 133.675 ;
        RECT 105.105 133.265 105.355 133.865 ;
        RECT 105.525 133.845 105.735 134.665 ;
        RECT 106.430 133.900 106.885 134.665 ;
        RECT 107.160 134.285 108.460 134.495 ;
        RECT 108.715 134.305 109.045 134.665 ;
        RECT 108.290 134.135 108.460 134.285 ;
        RECT 109.215 134.165 109.475 134.495 ;
        RECT 107.360 133.675 107.580 134.075 ;
        RECT 106.425 133.475 106.915 133.675 ;
        RECT 107.105 133.465 107.580 133.675 ;
        RECT 107.825 133.675 108.035 134.075 ;
        RECT 108.290 134.010 109.045 134.135 ;
        RECT 108.290 133.965 109.135 134.010 ;
        RECT 108.865 133.845 109.135 133.965 ;
        RECT 107.825 133.465 108.155 133.675 ;
        RECT 108.325 133.405 108.735 133.710 ;
        RECT 101.365 132.795 103.585 132.965 ;
        RECT 103.755 132.795 104.415 132.995 ;
        RECT 101.365 132.115 101.665 132.625 ;
        RECT 101.835 132.285 102.165 132.795 ;
        RECT 103.755 132.625 103.925 132.795 ;
        RECT 102.335 132.115 102.965 132.625 ;
        RECT 103.545 132.455 103.925 132.625 ;
        RECT 104.095 132.115 104.395 132.625 ;
        RECT 104.625 132.115 104.855 133.255 ;
        RECT 105.025 132.285 105.355 133.265 ;
        RECT 105.525 132.115 105.735 133.255 ;
        RECT 106.430 133.235 107.605 133.295 ;
        RECT 108.965 133.270 109.135 133.845 ;
        RECT 108.935 133.235 109.135 133.270 ;
        RECT 106.430 133.125 109.135 133.235 ;
        RECT 106.430 132.505 106.685 133.125 ;
        RECT 107.275 133.065 109.075 133.125 ;
        RECT 107.275 133.035 107.605 133.065 ;
        RECT 109.305 132.965 109.475 134.165 ;
        RECT 109.845 134.035 110.175 134.395 ;
        RECT 110.795 134.205 111.045 134.665 ;
        RECT 111.215 134.205 111.775 134.495 ;
        RECT 109.845 133.845 111.235 134.035 ;
        RECT 111.065 133.755 111.235 133.845 ;
        RECT 109.660 133.425 110.335 133.675 ;
        RECT 110.555 133.425 110.895 133.675 ;
        RECT 111.065 133.425 111.355 133.755 ;
        RECT 109.660 133.065 109.925 133.425 ;
        RECT 111.065 133.175 111.235 133.425 ;
        RECT 106.935 132.865 107.120 132.955 ;
        RECT 107.710 132.865 108.545 132.875 ;
        RECT 106.935 132.665 108.545 132.865 ;
        RECT 106.935 132.625 107.165 132.665 ;
        RECT 106.430 132.285 106.765 132.505 ;
        RECT 107.770 132.115 108.125 132.495 ;
        RECT 108.295 132.285 108.545 132.665 ;
        RECT 108.795 132.115 109.045 132.895 ;
        RECT 109.215 132.285 109.475 132.965 ;
        RECT 110.295 133.005 111.235 133.175 ;
        RECT 109.845 132.115 110.125 132.785 ;
        RECT 110.295 132.455 110.595 133.005 ;
        RECT 111.525 132.835 111.775 134.205 ;
        RECT 112.035 134.115 112.205 134.495 ;
        RECT 112.385 134.285 112.715 134.665 ;
        RECT 112.035 133.945 112.700 134.115 ;
        RECT 112.895 133.990 113.155 134.495 ;
        RECT 111.965 133.395 112.295 133.765 ;
        RECT 112.530 133.690 112.700 133.945 ;
        RECT 112.530 133.360 112.815 133.690 ;
        RECT 112.530 133.215 112.700 133.360 ;
        RECT 110.795 132.115 111.125 132.835 ;
        RECT 111.315 132.285 111.775 132.835 ;
        RECT 112.035 133.045 112.700 133.215 ;
        RECT 112.985 133.190 113.155 133.990 ;
        RECT 114.245 133.940 114.535 134.665 ;
        RECT 114.705 134.120 120.050 134.665 ;
        RECT 120.225 134.120 125.570 134.665 ;
        RECT 125.745 134.120 131.090 134.665 ;
        RECT 131.265 134.120 136.610 134.665 ;
        RECT 116.290 133.290 116.630 134.120 ;
        RECT 112.035 132.285 112.205 133.045 ;
        RECT 112.385 132.115 112.715 132.875 ;
        RECT 112.885 132.285 113.155 133.190 ;
        RECT 114.245 132.115 114.535 133.280 ;
        RECT 118.110 132.550 118.460 133.800 ;
        RECT 121.810 133.290 122.150 134.120 ;
        RECT 123.630 132.550 123.980 133.800 ;
        RECT 127.330 133.290 127.670 134.120 ;
        RECT 129.150 132.550 129.500 133.800 ;
        RECT 132.850 133.290 133.190 134.120 ;
        RECT 136.785 133.895 139.375 134.665 ;
        RECT 140.005 133.940 140.295 134.665 ;
        RECT 140.465 134.120 145.810 134.665 ;
        RECT 134.670 132.550 135.020 133.800 ;
        RECT 136.785 133.375 137.995 133.895 ;
        RECT 138.165 133.205 139.375 133.725 ;
        RECT 142.050 133.290 142.390 134.120 ;
        RECT 145.985 133.895 148.575 134.665 ;
        RECT 149.205 133.915 150.415 134.665 ;
        RECT 114.705 132.115 120.050 132.550 ;
        RECT 120.225 132.115 125.570 132.550 ;
        RECT 125.745 132.115 131.090 132.550 ;
        RECT 131.265 132.115 136.610 132.550 ;
        RECT 136.785 132.115 139.375 133.205 ;
        RECT 140.005 132.115 140.295 133.280 ;
        RECT 143.870 132.550 144.220 133.800 ;
        RECT 145.985 133.375 147.195 133.895 ;
        RECT 147.365 133.205 148.575 133.725 ;
        RECT 140.465 132.115 145.810 132.550 ;
        RECT 145.985 132.115 148.575 133.205 ;
        RECT 149.205 133.205 149.725 133.745 ;
        RECT 149.895 133.375 150.415 133.915 ;
        RECT 149.205 132.115 150.415 133.205 ;
        RECT 11.120 131.945 150.500 132.115 ;
        RECT 11.205 130.855 12.415 131.945 ;
        RECT 12.585 131.510 17.930 131.945 ;
        RECT 18.105 131.510 23.450 131.945 ;
        RECT 11.205 130.145 11.725 130.685 ;
        RECT 11.895 130.315 12.415 130.855 ;
        RECT 11.205 129.395 12.415 130.145 ;
        RECT 14.170 129.940 14.510 130.770 ;
        RECT 15.990 130.260 16.340 131.510 ;
        RECT 19.690 129.940 20.030 130.770 ;
        RECT 21.510 130.260 21.860 131.510 ;
        RECT 24.085 130.780 24.375 131.945 ;
        RECT 24.545 130.855 27.135 131.945 ;
        RECT 27.365 130.885 27.695 131.730 ;
        RECT 27.865 130.935 28.035 131.945 ;
        RECT 28.205 131.215 28.545 131.775 ;
        RECT 28.775 131.445 29.090 131.945 ;
        RECT 29.270 131.475 30.155 131.645 ;
        RECT 24.545 130.165 25.755 130.685 ;
        RECT 25.925 130.335 27.135 130.855 ;
        RECT 27.305 130.805 27.695 130.885 ;
        RECT 28.205 130.840 29.100 131.215 ;
        RECT 27.305 130.755 27.520 130.805 ;
        RECT 27.305 130.175 27.475 130.755 ;
        RECT 28.205 130.635 28.395 130.840 ;
        RECT 29.270 130.635 29.440 131.475 ;
        RECT 30.380 131.445 30.630 131.775 ;
        RECT 27.645 130.305 28.395 130.635 ;
        RECT 28.565 130.305 29.440 130.635 ;
        RECT 12.585 129.395 17.930 129.940 ;
        RECT 18.105 129.395 23.450 129.940 ;
        RECT 24.085 129.395 24.375 130.120 ;
        RECT 24.545 129.395 27.135 130.165 ;
        RECT 27.305 130.135 27.530 130.175 ;
        RECT 28.195 130.135 28.395 130.305 ;
        RECT 27.305 130.050 27.685 130.135 ;
        RECT 27.355 129.615 27.685 130.050 ;
        RECT 27.855 129.395 28.025 130.005 ;
        RECT 28.195 129.610 28.525 130.135 ;
        RECT 28.785 129.395 28.995 129.925 ;
        RECT 29.270 129.845 29.440 130.305 ;
        RECT 29.610 130.345 29.930 131.305 ;
        RECT 30.100 130.555 30.290 131.275 ;
        RECT 30.460 130.375 30.630 131.445 ;
        RECT 30.800 131.145 30.970 131.945 ;
        RECT 31.140 131.500 32.245 131.670 ;
        RECT 31.140 130.885 31.310 131.500 ;
        RECT 32.455 131.350 32.705 131.775 ;
        RECT 32.875 131.485 33.140 131.945 ;
        RECT 31.480 130.965 32.010 131.330 ;
        RECT 32.455 131.220 32.760 131.350 ;
        RECT 30.800 130.795 31.310 130.885 ;
        RECT 30.800 130.625 31.670 130.795 ;
        RECT 30.800 130.555 30.970 130.625 ;
        RECT 31.090 130.375 31.290 130.405 ;
        RECT 29.610 130.015 30.075 130.345 ;
        RECT 30.460 130.075 31.290 130.375 ;
        RECT 30.460 129.845 30.630 130.075 ;
        RECT 29.270 129.675 30.055 129.845 ;
        RECT 30.225 129.675 30.630 129.845 ;
        RECT 30.810 129.395 31.180 129.895 ;
        RECT 31.500 129.845 31.670 130.625 ;
        RECT 31.840 130.265 32.010 130.965 ;
        RECT 32.180 130.435 32.420 131.030 ;
        RECT 31.840 130.045 32.365 130.265 ;
        RECT 32.590 130.115 32.760 131.220 ;
        RECT 32.535 129.985 32.760 130.115 ;
        RECT 32.930 130.025 33.210 130.975 ;
        RECT 32.535 129.845 32.705 129.985 ;
        RECT 31.500 129.675 32.175 129.845 ;
        RECT 32.370 129.675 32.705 129.845 ;
        RECT 32.875 129.395 33.125 129.855 ;
        RECT 33.380 129.655 33.565 131.775 ;
        RECT 33.735 131.445 34.065 131.945 ;
        RECT 34.235 131.275 34.405 131.775 ;
        RECT 34.665 131.510 40.010 131.945 ;
        RECT 33.740 131.105 34.405 131.275 ;
        RECT 33.740 130.115 33.970 131.105 ;
        RECT 34.140 130.285 34.490 130.935 ;
        RECT 33.740 129.945 34.405 130.115 ;
        RECT 33.735 129.395 34.065 129.775 ;
        RECT 34.235 129.655 34.405 129.945 ;
        RECT 36.250 129.940 36.590 130.770 ;
        RECT 38.070 130.260 38.420 131.510 ;
        RECT 40.185 130.855 41.855 131.945 ;
        RECT 40.185 130.165 40.935 130.685 ;
        RECT 41.105 130.335 41.855 130.855 ;
        RECT 34.665 129.395 40.010 129.940 ;
        RECT 40.185 129.395 41.855 130.165 ;
        RECT 42.025 129.675 42.305 131.775 ;
        RECT 42.495 131.185 43.280 131.945 ;
        RECT 43.675 131.115 44.060 131.775 ;
        RECT 43.675 131.015 44.085 131.115 ;
        RECT 42.475 130.805 44.085 131.015 ;
        RECT 44.385 130.925 44.585 131.715 ;
        RECT 42.475 130.205 42.750 130.805 ;
        RECT 44.255 130.755 44.585 130.925 ;
        RECT 44.755 130.765 45.075 131.945 ;
        RECT 45.245 130.855 48.755 131.945 ;
        RECT 44.255 130.635 44.435 130.755 ;
        RECT 42.920 130.385 43.275 130.635 ;
        RECT 43.470 130.585 43.935 130.635 ;
        RECT 43.465 130.415 43.935 130.585 ;
        RECT 43.470 130.385 43.935 130.415 ;
        RECT 44.105 130.385 44.435 130.635 ;
        RECT 44.610 130.385 45.075 130.585 ;
        RECT 42.475 130.025 43.725 130.205 ;
        RECT 43.360 129.955 43.725 130.025 ;
        RECT 43.895 130.005 45.075 130.175 ;
        RECT 42.535 129.395 42.705 129.855 ;
        RECT 43.895 129.785 44.225 130.005 ;
        RECT 42.975 129.605 44.225 129.785 ;
        RECT 44.395 129.395 44.565 129.835 ;
        RECT 44.735 129.590 45.075 130.005 ;
        RECT 45.245 130.165 46.895 130.685 ;
        RECT 47.065 130.335 48.755 130.855 ;
        RECT 49.845 130.780 50.135 131.945 ;
        RECT 50.305 130.855 51.975 131.945 ;
        RECT 50.305 130.165 51.055 130.685 ;
        RECT 51.225 130.335 51.975 130.855 ;
        RECT 52.615 130.995 52.890 131.765 ;
        RECT 53.060 131.335 53.390 131.765 ;
        RECT 53.560 131.505 53.755 131.945 ;
        RECT 53.935 131.335 54.265 131.765 ;
        RECT 53.060 131.165 54.265 131.335 ;
        RECT 52.615 130.805 53.200 130.995 ;
        RECT 53.370 130.835 54.265 131.165 ;
        RECT 54.455 130.885 54.785 131.735 ;
        RECT 45.245 129.395 48.755 130.165 ;
        RECT 49.845 129.395 50.135 130.120 ;
        RECT 50.305 129.395 51.975 130.165 ;
        RECT 52.615 129.985 52.855 130.635 ;
        RECT 53.025 130.135 53.200 130.805 ;
        RECT 53.370 130.305 53.785 130.635 ;
        RECT 53.965 130.305 54.260 130.635 ;
        RECT 53.025 129.955 53.355 130.135 ;
        RECT 52.630 129.395 52.960 129.785 ;
        RECT 53.130 129.575 53.355 129.955 ;
        RECT 53.555 129.685 53.785 130.305 ;
        RECT 53.965 129.395 54.265 130.125 ;
        RECT 54.455 130.120 54.645 130.885 ;
        RECT 54.955 130.805 55.205 131.945 ;
        RECT 55.395 131.305 55.645 131.725 ;
        RECT 55.875 131.475 56.205 131.945 ;
        RECT 56.435 131.305 56.685 131.725 ;
        RECT 55.395 131.135 56.685 131.305 ;
        RECT 56.865 131.305 57.195 131.735 ;
        RECT 56.865 131.135 57.320 131.305 ;
        RECT 55.385 130.635 55.600 130.965 ;
        RECT 54.815 130.305 55.125 130.635 ;
        RECT 55.295 130.305 55.600 130.635 ;
        RECT 55.775 130.305 56.060 130.965 ;
        RECT 56.255 130.305 56.520 130.965 ;
        RECT 56.735 130.305 56.980 130.965 ;
        RECT 54.955 130.135 55.125 130.305 ;
        RECT 57.150 130.135 57.320 131.135 ;
        RECT 58.585 130.805 58.845 131.945 ;
        RECT 59.085 131.435 60.700 131.765 ;
        RECT 59.095 130.635 59.265 131.195 ;
        RECT 59.525 131.095 60.700 131.265 ;
        RECT 60.870 131.145 61.150 131.945 ;
        RECT 59.525 130.805 59.855 131.095 ;
        RECT 60.530 130.975 60.700 131.095 ;
        RECT 60.025 130.635 60.270 130.925 ;
        RECT 60.530 130.805 61.190 130.975 ;
        RECT 61.360 130.805 61.635 131.775 ;
        RECT 61.805 131.510 67.150 131.945 ;
        RECT 61.020 130.635 61.190 130.805 ;
        RECT 58.590 130.385 58.925 130.635 ;
        RECT 59.095 130.305 59.810 130.635 ;
        RECT 60.025 130.305 60.850 130.635 ;
        RECT 61.020 130.305 61.295 130.635 ;
        RECT 59.095 130.215 59.345 130.305 ;
        RECT 54.455 129.610 54.785 130.120 ;
        RECT 54.955 129.965 57.320 130.135 ;
        RECT 54.955 129.395 55.285 129.795 ;
        RECT 56.335 129.625 56.665 129.965 ;
        RECT 56.835 129.395 57.165 129.795 ;
        RECT 58.585 129.395 58.845 130.215 ;
        RECT 59.015 129.795 59.345 130.215 ;
        RECT 61.020 130.135 61.190 130.305 ;
        RECT 59.525 129.965 61.190 130.135 ;
        RECT 61.465 130.070 61.635 130.805 ;
        RECT 59.525 129.565 59.785 129.965 ;
        RECT 59.955 129.395 60.285 129.795 ;
        RECT 60.455 129.615 60.625 129.965 ;
        RECT 60.795 129.395 61.170 129.795 ;
        RECT 61.360 129.725 61.635 130.070 ;
        RECT 63.390 129.940 63.730 130.770 ;
        RECT 65.210 130.260 65.560 131.510 ;
        RECT 67.360 131.155 67.895 131.775 ;
        RECT 67.360 130.135 67.675 131.155 ;
        RECT 68.065 131.145 68.395 131.945 ;
        RECT 68.880 130.975 69.270 131.150 ;
        RECT 67.845 130.805 69.270 130.975 ;
        RECT 69.625 130.855 73.135 131.945 ;
        RECT 67.845 130.305 68.015 130.805 ;
        RECT 61.805 129.395 67.150 129.940 ;
        RECT 67.360 129.565 67.975 130.135 ;
        RECT 68.265 130.075 68.530 130.635 ;
        RECT 68.700 129.905 68.870 130.805 ;
        RECT 69.040 130.075 69.395 130.635 ;
        RECT 69.625 130.165 71.275 130.685 ;
        RECT 71.445 130.335 73.135 130.855 ;
        RECT 73.775 130.995 74.050 131.765 ;
        RECT 74.220 131.335 74.550 131.765 ;
        RECT 74.720 131.505 74.915 131.945 ;
        RECT 75.095 131.335 75.425 131.765 ;
        RECT 74.220 131.165 75.425 131.335 ;
        RECT 73.775 130.805 74.360 130.995 ;
        RECT 74.530 130.835 75.425 131.165 ;
        RECT 68.145 129.395 68.360 129.905 ;
        RECT 68.590 129.575 68.870 129.905 ;
        RECT 69.050 129.395 69.290 129.905 ;
        RECT 69.625 129.395 73.135 130.165 ;
        RECT 73.775 129.985 74.015 130.635 ;
        RECT 74.185 130.135 74.360 130.805 ;
        RECT 75.605 130.780 75.895 131.945 ;
        RECT 76.065 131.105 76.325 131.775 ;
        RECT 76.495 131.545 76.825 131.945 ;
        RECT 77.695 131.545 78.095 131.945 ;
        RECT 78.385 131.365 78.715 131.600 ;
        RECT 76.635 131.195 78.715 131.365 ;
        RECT 74.530 130.305 74.945 130.635 ;
        RECT 75.125 130.305 75.420 130.635 ;
        RECT 74.185 129.955 74.515 130.135 ;
        RECT 73.790 129.395 74.120 129.785 ;
        RECT 74.290 129.575 74.515 129.955 ;
        RECT 74.715 129.685 74.945 130.305 ;
        RECT 76.065 130.135 76.240 131.105 ;
        RECT 76.635 130.925 76.805 131.195 ;
        RECT 76.410 130.755 76.805 130.925 ;
        RECT 76.975 130.805 77.990 131.025 ;
        RECT 76.410 130.305 76.580 130.755 ;
        RECT 77.715 130.665 77.990 130.805 ;
        RECT 78.160 130.805 78.715 131.195 ;
        RECT 76.750 130.385 77.200 130.585 ;
        RECT 77.370 130.215 77.545 130.410 ;
        RECT 75.125 129.395 75.425 130.125 ;
        RECT 75.605 129.395 75.895 130.120 ;
        RECT 76.065 129.565 76.405 130.135 ;
        RECT 76.600 129.395 76.770 130.060 ;
        RECT 77.050 130.045 77.545 130.215 ;
        RECT 77.050 129.905 77.270 130.045 ;
        RECT 77.045 129.735 77.270 129.905 ;
        RECT 77.715 129.875 77.885 130.665 ;
        RECT 78.160 130.555 78.330 130.805 ;
        RECT 78.885 130.635 79.060 131.735 ;
        RECT 79.230 131.125 79.575 131.945 ;
        RECT 79.930 130.975 80.320 131.150 ;
        RECT 80.805 131.145 81.135 131.945 ;
        RECT 81.305 131.155 81.840 131.775 ;
        RECT 78.135 130.385 78.330 130.555 ;
        RECT 78.500 130.385 79.060 130.635 ;
        RECT 79.230 130.385 79.575 130.955 ;
        RECT 79.930 130.805 81.355 130.975 ;
        RECT 78.135 130.000 78.305 130.385 ;
        RECT 77.050 129.690 77.270 129.735 ;
        RECT 77.440 129.705 77.885 129.875 ;
        RECT 78.055 129.630 78.305 130.000 ;
        RECT 78.475 130.035 79.575 130.215 ;
        RECT 79.805 130.075 80.160 130.635 ;
        RECT 78.475 129.630 78.725 130.035 ;
        RECT 78.895 129.395 79.065 129.865 ;
        RECT 79.235 129.630 79.575 130.035 ;
        RECT 80.330 129.905 80.500 130.805 ;
        RECT 80.670 130.075 80.935 130.635 ;
        RECT 81.185 130.305 81.355 130.805 ;
        RECT 81.525 130.135 81.840 131.155 ;
        RECT 82.045 130.855 83.255 131.945 ;
        RECT 83.430 131.565 83.765 131.945 ;
        RECT 79.910 129.395 80.150 129.905 ;
        RECT 80.330 129.575 80.610 129.905 ;
        RECT 80.840 129.395 81.055 129.905 ;
        RECT 81.225 129.565 81.840 130.135 ;
        RECT 82.045 130.145 82.565 130.685 ;
        RECT 82.735 130.315 83.255 130.855 ;
        RECT 82.045 129.395 83.255 130.145 ;
        RECT 83.425 130.075 83.665 131.385 ;
        RECT 83.935 130.975 84.185 131.775 ;
        RECT 84.405 131.225 84.735 131.945 ;
        RECT 84.920 130.975 85.170 131.775 ;
        RECT 85.635 131.145 85.965 131.945 ;
        RECT 86.135 131.515 86.475 131.775 ;
        RECT 83.835 130.805 86.025 130.975 ;
        RECT 83.835 129.895 84.005 130.805 ;
        RECT 85.710 130.635 86.025 130.805 ;
        RECT 83.510 129.565 84.005 129.895 ;
        RECT 84.225 129.670 84.575 130.635 ;
        RECT 84.755 129.665 85.055 130.635 ;
        RECT 85.235 129.665 85.515 130.635 ;
        RECT 85.710 130.385 86.040 130.635 ;
        RECT 85.695 129.395 85.965 130.195 ;
        RECT 86.215 130.115 86.475 131.515 ;
        RECT 86.650 131.555 86.985 131.775 ;
        RECT 87.990 131.565 88.345 131.945 ;
        RECT 86.650 130.935 86.905 131.555 ;
        RECT 87.155 131.395 87.385 131.435 ;
        RECT 88.515 131.395 88.765 131.775 ;
        RECT 87.155 131.195 88.765 131.395 ;
        RECT 87.155 131.105 87.340 131.195 ;
        RECT 87.930 131.185 88.765 131.195 ;
        RECT 89.015 131.165 89.265 131.945 ;
        RECT 89.435 131.095 89.695 131.775 ;
        RECT 89.865 131.510 95.210 131.945 ;
        RECT 87.495 130.995 87.825 131.025 ;
        RECT 87.495 130.935 89.295 130.995 ;
        RECT 86.650 130.825 89.355 130.935 ;
        RECT 86.650 130.765 87.825 130.825 ;
        RECT 89.155 130.790 89.355 130.825 ;
        RECT 86.645 130.385 87.135 130.585 ;
        RECT 87.325 130.385 87.800 130.595 ;
        RECT 86.135 129.605 86.475 130.115 ;
        RECT 86.650 129.395 87.105 130.160 ;
        RECT 87.580 129.985 87.800 130.385 ;
        RECT 88.045 130.385 88.375 130.595 ;
        RECT 88.045 129.985 88.255 130.385 ;
        RECT 88.545 130.350 88.955 130.655 ;
        RECT 89.185 130.215 89.355 130.790 ;
        RECT 89.085 130.095 89.355 130.215 ;
        RECT 88.510 130.050 89.355 130.095 ;
        RECT 88.510 129.925 89.265 130.050 ;
        RECT 88.510 129.775 88.680 129.925 ;
        RECT 89.525 129.905 89.695 131.095 ;
        RECT 91.450 129.940 91.790 130.770 ;
        RECT 93.270 130.260 93.620 131.510 ;
        RECT 95.385 130.855 97.055 131.945 ;
        RECT 95.385 130.165 96.135 130.685 ;
        RECT 96.305 130.335 97.055 130.855 ;
        RECT 97.685 131.095 98.065 131.775 ;
        RECT 98.655 131.095 98.825 131.945 ;
        RECT 98.995 131.265 99.325 131.775 ;
        RECT 99.495 131.435 99.665 131.945 ;
        RECT 99.835 131.265 100.235 131.775 ;
        RECT 98.995 131.095 100.235 131.265 ;
        RECT 89.465 129.895 89.695 129.905 ;
        RECT 87.380 129.565 88.680 129.775 ;
        RECT 88.935 129.395 89.265 129.755 ;
        RECT 89.435 129.565 89.695 129.895 ;
        RECT 89.865 129.395 95.210 129.940 ;
        RECT 95.385 129.395 97.055 130.165 ;
        RECT 97.685 130.135 97.855 131.095 ;
        RECT 98.025 130.755 99.330 130.925 ;
        RECT 100.415 130.845 100.735 131.775 ;
        RECT 98.025 130.305 98.270 130.755 ;
        RECT 98.440 130.385 98.990 130.585 ;
        RECT 99.160 130.555 99.330 130.755 ;
        RECT 100.105 130.675 100.735 130.845 ;
        RECT 101.365 130.780 101.655 131.945 ;
        RECT 101.825 130.855 105.335 131.945 ;
        RECT 105.505 130.855 106.715 131.945 ;
        RECT 107.065 131.030 107.235 131.945 ;
        RECT 107.405 130.885 107.735 131.730 ;
        RECT 107.905 130.935 108.075 131.945 ;
        RECT 108.245 131.215 108.585 131.775 ;
        RECT 108.815 131.445 109.130 131.945 ;
        RECT 109.310 131.475 110.195 131.645 ;
        RECT 99.160 130.385 99.535 130.555 ;
        RECT 99.705 130.135 99.935 130.635 ;
        RECT 97.685 129.965 99.935 130.135 ;
        RECT 97.735 129.395 98.065 129.785 ;
        RECT 98.235 129.645 98.405 129.965 ;
        RECT 100.105 129.795 100.275 130.675 ;
        RECT 98.575 129.395 98.905 129.785 ;
        RECT 99.320 129.625 100.275 129.795 ;
        RECT 100.445 129.395 100.735 130.230 ;
        RECT 101.825 130.165 103.475 130.685 ;
        RECT 103.645 130.335 105.335 130.855 ;
        RECT 101.365 129.395 101.655 130.120 ;
        RECT 101.825 129.395 105.335 130.165 ;
        RECT 105.505 130.145 106.025 130.685 ;
        RECT 106.195 130.315 106.715 130.855 ;
        RECT 107.345 130.805 107.735 130.885 ;
        RECT 108.245 130.840 109.140 131.215 ;
        RECT 107.345 130.755 107.560 130.805 ;
        RECT 107.345 130.175 107.515 130.755 ;
        RECT 108.245 130.635 108.435 130.840 ;
        RECT 109.310 130.635 109.480 131.475 ;
        RECT 110.420 131.445 110.670 131.775 ;
        RECT 107.685 130.305 108.435 130.635 ;
        RECT 108.605 130.305 109.480 130.635 ;
        RECT 105.505 129.395 106.715 130.145 ;
        RECT 107.345 130.135 107.570 130.175 ;
        RECT 108.235 130.135 108.435 130.305 ;
        RECT 107.345 130.050 107.725 130.135 ;
        RECT 107.055 129.395 107.225 129.910 ;
        RECT 107.395 129.615 107.725 130.050 ;
        RECT 107.895 129.395 108.065 130.005 ;
        RECT 108.235 129.610 108.565 130.135 ;
        RECT 108.825 129.395 109.035 129.925 ;
        RECT 109.310 129.845 109.480 130.305 ;
        RECT 109.650 130.345 109.970 131.305 ;
        RECT 110.140 130.555 110.330 131.275 ;
        RECT 110.500 130.375 110.670 131.445 ;
        RECT 110.840 131.145 111.010 131.945 ;
        RECT 111.180 131.500 112.285 131.670 ;
        RECT 111.180 130.885 111.350 131.500 ;
        RECT 112.495 131.350 112.745 131.775 ;
        RECT 112.915 131.485 113.180 131.945 ;
        RECT 111.520 130.965 112.050 131.330 ;
        RECT 112.495 131.220 112.800 131.350 ;
        RECT 110.840 130.795 111.350 130.885 ;
        RECT 110.840 130.625 111.710 130.795 ;
        RECT 110.840 130.555 111.010 130.625 ;
        RECT 111.130 130.375 111.330 130.405 ;
        RECT 109.650 130.015 110.115 130.345 ;
        RECT 110.500 130.075 111.330 130.375 ;
        RECT 110.500 129.845 110.670 130.075 ;
        RECT 109.310 129.675 110.095 129.845 ;
        RECT 110.265 129.675 110.670 129.845 ;
        RECT 110.850 129.395 111.220 129.895 ;
        RECT 111.540 129.845 111.710 130.625 ;
        RECT 111.880 130.265 112.050 130.965 ;
        RECT 112.220 130.435 112.460 131.030 ;
        RECT 111.880 130.045 112.405 130.265 ;
        RECT 112.630 130.115 112.800 131.220 ;
        RECT 112.575 129.985 112.800 130.115 ;
        RECT 112.970 130.025 113.250 130.975 ;
        RECT 112.575 129.845 112.745 129.985 ;
        RECT 111.540 129.675 112.215 129.845 ;
        RECT 112.410 129.675 112.745 129.845 ;
        RECT 112.915 129.395 113.165 129.855 ;
        RECT 113.420 129.655 113.605 131.775 ;
        RECT 113.775 131.445 114.105 131.945 ;
        RECT 114.275 131.275 114.445 131.775 ;
        RECT 114.705 131.510 120.050 131.945 ;
        RECT 120.225 131.510 125.570 131.945 ;
        RECT 113.780 131.105 114.445 131.275 ;
        RECT 113.780 130.115 114.010 131.105 ;
        RECT 114.180 130.285 114.530 130.935 ;
        RECT 113.780 129.945 114.445 130.115 ;
        RECT 113.775 129.395 114.105 129.775 ;
        RECT 114.275 129.655 114.445 129.945 ;
        RECT 116.290 129.940 116.630 130.770 ;
        RECT 118.110 130.260 118.460 131.510 ;
        RECT 121.810 129.940 122.150 130.770 ;
        RECT 123.630 130.260 123.980 131.510 ;
        RECT 125.745 130.855 126.955 131.945 ;
        RECT 125.745 130.145 126.265 130.685 ;
        RECT 126.435 130.315 126.955 130.855 ;
        RECT 127.125 130.780 127.415 131.945 ;
        RECT 127.585 131.510 132.930 131.945 ;
        RECT 133.105 131.510 138.450 131.945 ;
        RECT 138.625 131.510 143.970 131.945 ;
        RECT 114.705 129.395 120.050 129.940 ;
        RECT 120.225 129.395 125.570 129.940 ;
        RECT 125.745 129.395 126.955 130.145 ;
        RECT 127.125 129.395 127.415 130.120 ;
        RECT 129.170 129.940 129.510 130.770 ;
        RECT 130.990 130.260 131.340 131.510 ;
        RECT 134.690 129.940 135.030 130.770 ;
        RECT 136.510 130.260 136.860 131.510 ;
        RECT 140.210 129.940 140.550 130.770 ;
        RECT 142.030 130.260 142.380 131.510 ;
        RECT 144.145 130.855 147.655 131.945 ;
        RECT 147.825 130.855 149.035 131.945 ;
        RECT 144.145 130.165 145.795 130.685 ;
        RECT 145.965 130.335 147.655 130.855 ;
        RECT 127.585 129.395 132.930 129.940 ;
        RECT 133.105 129.395 138.450 129.940 ;
        RECT 138.625 129.395 143.970 129.940 ;
        RECT 144.145 129.395 147.655 130.165 ;
        RECT 147.825 130.145 148.345 130.685 ;
        RECT 148.515 130.315 149.035 130.855 ;
        RECT 149.205 130.855 150.415 131.945 ;
        RECT 149.205 130.315 149.725 130.855 ;
        RECT 149.895 130.145 150.415 130.685 ;
        RECT 147.825 129.395 149.035 130.145 ;
        RECT 149.205 129.395 150.415 130.145 ;
        RECT 11.120 129.225 150.500 129.395 ;
        RECT 11.205 128.475 12.415 129.225 ;
        RECT 12.585 128.680 17.930 129.225 ;
        RECT 18.105 128.680 23.450 129.225 ;
        RECT 23.625 128.680 28.970 129.225 ;
        RECT 29.145 128.680 34.490 129.225 ;
        RECT 11.205 127.935 11.725 128.475 ;
        RECT 11.895 127.765 12.415 128.305 ;
        RECT 14.170 127.850 14.510 128.680 ;
        RECT 11.205 126.675 12.415 127.765 ;
        RECT 15.990 127.110 16.340 128.360 ;
        RECT 19.690 127.850 20.030 128.680 ;
        RECT 21.510 127.110 21.860 128.360 ;
        RECT 25.210 127.850 25.550 128.680 ;
        RECT 27.030 127.110 27.380 128.360 ;
        RECT 30.730 127.850 31.070 128.680 ;
        RECT 34.665 128.455 36.335 129.225 ;
        RECT 36.965 128.500 37.255 129.225 ;
        RECT 37.425 128.455 40.935 129.225 ;
        RECT 42.190 128.715 42.430 129.225 ;
        RECT 42.610 128.715 42.890 129.045 ;
        RECT 43.120 128.715 43.335 129.225 ;
        RECT 32.550 127.110 32.900 128.360 ;
        RECT 34.665 127.935 35.415 128.455 ;
        RECT 35.585 127.765 36.335 128.285 ;
        RECT 37.425 127.935 39.075 128.455 ;
        RECT 12.585 126.675 17.930 127.110 ;
        RECT 18.105 126.675 23.450 127.110 ;
        RECT 23.625 126.675 28.970 127.110 ;
        RECT 29.145 126.675 34.490 127.110 ;
        RECT 34.665 126.675 36.335 127.765 ;
        RECT 36.965 126.675 37.255 127.840 ;
        RECT 39.245 127.765 40.935 128.285 ;
        RECT 42.085 127.985 42.440 128.545 ;
        RECT 42.610 127.815 42.780 128.715 ;
        RECT 42.950 127.985 43.215 128.545 ;
        RECT 43.505 128.485 44.120 129.055 ;
        RECT 44.415 128.675 44.585 129.055 ;
        RECT 44.765 128.845 45.095 129.225 ;
        RECT 44.415 128.505 45.080 128.675 ;
        RECT 45.275 128.550 45.535 129.055 ;
        RECT 43.465 127.815 43.635 128.315 ;
        RECT 37.425 126.675 40.935 127.765 ;
        RECT 42.210 127.645 43.635 127.815 ;
        RECT 42.210 127.470 42.600 127.645 ;
        RECT 43.085 126.675 43.415 127.475 ;
        RECT 43.805 127.465 44.120 128.485 ;
        RECT 44.345 127.955 44.675 128.325 ;
        RECT 44.910 128.250 45.080 128.505 ;
        RECT 44.910 127.920 45.195 128.250 ;
        RECT 44.910 127.775 45.080 127.920 ;
        RECT 43.585 126.845 44.120 127.465 ;
        RECT 44.415 127.605 45.080 127.775 ;
        RECT 45.365 127.750 45.535 128.550 ;
        RECT 45.705 128.455 48.295 129.225 ;
        RECT 45.705 127.935 46.915 128.455 ;
        RECT 48.935 128.415 49.205 129.225 ;
        RECT 49.375 128.415 49.705 129.055 ;
        RECT 49.875 128.415 50.115 129.225 ;
        RECT 50.765 128.485 51.105 129.055 ;
        RECT 51.300 128.560 51.470 129.225 ;
        RECT 51.750 128.885 51.970 128.930 ;
        RECT 51.745 128.715 51.970 128.885 ;
        RECT 52.140 128.745 52.585 128.915 ;
        RECT 51.750 128.575 51.970 128.715 ;
        RECT 47.085 127.765 48.295 128.285 ;
        RECT 48.925 127.985 49.275 128.235 ;
        RECT 49.445 127.815 49.615 128.415 ;
        RECT 49.785 127.985 50.135 128.235 ;
        RECT 44.415 126.845 44.585 127.605 ;
        RECT 44.765 126.675 45.095 127.435 ;
        RECT 45.265 126.845 45.535 127.750 ;
        RECT 45.705 126.675 48.295 127.765 ;
        RECT 48.935 126.675 49.265 127.815 ;
        RECT 49.445 127.645 50.125 127.815 ;
        RECT 49.795 126.860 50.125 127.645 ;
        RECT 50.765 127.525 50.940 128.485 ;
        RECT 51.750 128.405 52.245 128.575 ;
        RECT 51.110 127.865 51.280 128.315 ;
        RECT 51.450 128.035 51.900 128.235 ;
        RECT 52.070 128.210 52.245 128.405 ;
        RECT 52.415 127.955 52.585 128.745 ;
        RECT 52.755 128.620 53.005 128.990 ;
        RECT 52.835 128.235 53.005 128.620 ;
        RECT 53.175 128.585 53.425 128.990 ;
        RECT 53.595 128.755 53.765 129.225 ;
        RECT 53.935 128.585 54.275 128.990 ;
        RECT 53.175 128.405 54.275 128.585 ;
        RECT 54.445 128.455 57.955 129.225 ;
        RECT 59.070 128.835 59.400 129.225 ;
        RECT 59.570 128.665 59.795 129.045 ;
        RECT 52.835 128.065 53.030 128.235 ;
        RECT 51.110 127.695 51.505 127.865 ;
        RECT 52.415 127.815 52.690 127.955 ;
        RECT 50.765 127.515 50.995 127.525 ;
        RECT 50.765 126.845 51.025 127.515 ;
        RECT 51.335 127.425 51.505 127.695 ;
        RECT 51.675 127.595 52.690 127.815 ;
        RECT 52.860 127.815 53.030 128.065 ;
        RECT 53.200 127.985 53.760 128.235 ;
        RECT 52.860 127.425 53.415 127.815 ;
        RECT 51.335 127.255 53.415 127.425 ;
        RECT 51.195 126.675 51.525 127.075 ;
        RECT 52.395 126.675 52.795 127.075 ;
        RECT 53.085 127.020 53.415 127.255 ;
        RECT 53.585 126.885 53.760 127.985 ;
        RECT 53.930 127.665 54.275 128.235 ;
        RECT 54.445 127.935 56.095 128.455 ;
        RECT 56.265 127.765 57.955 128.285 ;
        RECT 59.055 127.985 59.295 128.635 ;
        RECT 59.465 128.485 59.795 128.665 ;
        RECT 59.465 127.815 59.640 128.485 ;
        RECT 59.995 128.315 60.225 128.935 ;
        RECT 60.405 128.495 60.705 129.225 ;
        RECT 60.885 128.425 61.195 129.225 ;
        RECT 61.400 128.425 62.095 129.055 ;
        RECT 62.725 128.500 63.015 129.225 ;
        RECT 63.185 128.485 63.570 129.055 ;
        RECT 63.740 128.765 64.065 129.225 ;
        RECT 64.585 128.595 64.865 129.055 ;
        RECT 59.810 127.985 60.225 128.315 ;
        RECT 60.405 127.985 60.700 128.315 ;
        RECT 60.895 127.985 61.230 128.255 ;
        RECT 61.400 127.825 61.570 128.425 ;
        RECT 61.740 127.985 62.075 128.235 ;
        RECT 53.930 126.675 54.275 127.495 ;
        RECT 54.445 126.675 57.955 127.765 ;
        RECT 59.055 127.625 59.640 127.815 ;
        RECT 59.055 126.855 59.330 127.625 ;
        RECT 59.810 127.455 60.705 127.785 ;
        RECT 59.500 127.285 60.705 127.455 ;
        RECT 59.500 126.855 59.830 127.285 ;
        RECT 60.000 126.675 60.195 127.115 ;
        RECT 60.375 126.855 60.705 127.285 ;
        RECT 60.885 126.675 61.165 127.815 ;
        RECT 61.335 126.845 61.665 127.825 ;
        RECT 61.835 126.675 62.095 127.815 ;
        RECT 62.725 126.675 63.015 127.840 ;
        RECT 63.185 127.815 63.465 128.485 ;
        RECT 63.740 128.425 64.865 128.595 ;
        RECT 63.740 128.315 64.190 128.425 ;
        RECT 63.635 127.985 64.190 128.315 ;
        RECT 65.055 128.255 65.455 129.055 ;
        RECT 65.855 128.765 66.125 129.225 ;
        RECT 66.295 128.595 66.580 129.055 ;
        RECT 63.185 126.845 63.570 127.815 ;
        RECT 63.740 127.525 64.190 127.985 ;
        RECT 64.360 127.695 65.455 128.255 ;
        RECT 63.740 127.305 64.865 127.525 ;
        RECT 63.740 126.675 64.065 127.135 ;
        RECT 64.585 126.845 64.865 127.305 ;
        RECT 65.055 126.845 65.455 127.695 ;
        RECT 65.625 128.425 66.580 128.595 ;
        RECT 66.955 128.675 67.125 128.965 ;
        RECT 67.295 128.845 67.625 129.225 ;
        RECT 66.955 128.505 67.620 128.675 ;
        RECT 65.625 127.525 65.835 128.425 ;
        RECT 66.005 127.695 66.695 128.255 ;
        RECT 66.870 127.685 67.220 128.335 ;
        RECT 65.625 127.305 66.580 127.525 ;
        RECT 67.390 127.515 67.620 128.505 ;
        RECT 65.855 126.675 66.125 127.135 ;
        RECT 66.295 126.845 66.580 127.305 ;
        RECT 66.955 127.345 67.620 127.515 ;
        RECT 66.955 126.845 67.125 127.345 ;
        RECT 67.295 126.675 67.625 127.175 ;
        RECT 67.795 126.845 67.980 128.965 ;
        RECT 68.235 128.765 68.485 129.225 ;
        RECT 68.655 128.775 68.990 128.945 ;
        RECT 69.185 128.775 69.860 128.945 ;
        RECT 68.655 128.635 68.825 128.775 ;
        RECT 68.150 127.645 68.430 128.595 ;
        RECT 68.600 128.505 68.825 128.635 ;
        RECT 68.600 127.400 68.770 128.505 ;
        RECT 68.995 128.355 69.520 128.575 ;
        RECT 68.940 127.590 69.180 128.185 ;
        RECT 69.350 127.655 69.520 128.355 ;
        RECT 69.690 127.995 69.860 128.775 ;
        RECT 70.180 128.725 70.550 129.225 ;
        RECT 70.730 128.775 71.135 128.945 ;
        RECT 71.305 128.775 72.090 128.945 ;
        RECT 70.730 128.545 70.900 128.775 ;
        RECT 70.070 128.245 70.900 128.545 ;
        RECT 71.285 128.275 71.750 128.605 ;
        RECT 70.070 128.215 70.270 128.245 ;
        RECT 70.390 127.995 70.560 128.065 ;
        RECT 69.690 127.825 70.560 127.995 ;
        RECT 70.050 127.735 70.560 127.825 ;
        RECT 68.600 127.270 68.905 127.400 ;
        RECT 69.350 127.290 69.880 127.655 ;
        RECT 68.220 126.675 68.485 127.135 ;
        RECT 68.655 126.845 68.905 127.270 ;
        RECT 70.050 127.120 70.220 127.735 ;
        RECT 69.115 126.950 70.220 127.120 ;
        RECT 70.390 126.675 70.560 127.475 ;
        RECT 70.730 127.175 70.900 128.245 ;
        RECT 71.070 127.345 71.260 128.065 ;
        RECT 71.430 127.315 71.750 128.275 ;
        RECT 71.920 128.315 72.090 128.775 ;
        RECT 72.365 128.695 72.575 129.225 ;
        RECT 72.835 128.485 73.165 129.010 ;
        RECT 73.335 128.615 73.505 129.225 ;
        RECT 73.675 128.570 74.005 129.005 ;
        RECT 73.675 128.485 74.055 128.570 ;
        RECT 72.965 128.315 73.165 128.485 ;
        RECT 73.830 128.445 74.055 128.485 ;
        RECT 71.920 127.985 72.795 128.315 ;
        RECT 72.965 127.985 73.715 128.315 ;
        RECT 70.730 126.845 70.980 127.175 ;
        RECT 71.920 127.145 72.090 127.985 ;
        RECT 72.965 127.780 73.155 127.985 ;
        RECT 73.885 127.865 74.055 128.445 ;
        RECT 74.225 128.475 75.435 129.225 ;
        RECT 75.605 128.485 75.925 128.965 ;
        RECT 76.095 128.655 76.325 129.055 ;
        RECT 76.495 128.835 76.845 129.225 ;
        RECT 76.095 128.575 76.605 128.655 ;
        RECT 77.015 128.575 77.345 129.055 ;
        RECT 76.095 128.485 77.345 128.575 ;
        RECT 74.225 127.935 74.745 128.475 ;
        RECT 73.840 127.815 74.055 127.865 ;
        RECT 72.260 127.405 73.155 127.780 ;
        RECT 73.665 127.735 74.055 127.815 ;
        RECT 74.915 127.765 75.435 128.305 ;
        RECT 71.205 126.975 72.090 127.145 ;
        RECT 72.270 126.675 72.585 127.175 ;
        RECT 72.815 126.845 73.155 127.405 ;
        RECT 73.325 126.675 73.495 127.685 ;
        RECT 73.665 126.890 73.995 127.735 ;
        RECT 74.225 126.675 75.435 127.765 ;
        RECT 75.605 127.555 75.775 128.485 ;
        RECT 76.435 128.405 77.345 128.485 ;
        RECT 77.515 128.405 77.685 129.225 ;
        RECT 78.190 128.485 78.655 129.030 ;
        RECT 75.945 127.895 76.115 128.315 ;
        RECT 76.345 128.065 76.945 128.235 ;
        RECT 75.945 127.725 76.605 127.895 ;
        RECT 75.605 127.355 76.265 127.555 ;
        RECT 76.435 127.525 76.605 127.725 ;
        RECT 76.775 127.865 76.945 128.065 ;
        RECT 77.115 128.035 77.810 128.235 ;
        RECT 78.070 127.865 78.315 128.315 ;
        RECT 76.775 127.695 78.315 127.865 ;
        RECT 78.485 127.525 78.655 128.485 ;
        RECT 78.825 128.455 80.495 129.225 ;
        RECT 78.825 127.935 79.575 128.455 ;
        RECT 81.125 128.425 81.435 129.225 ;
        RECT 81.640 128.425 82.335 129.055 ;
        RECT 82.670 128.715 82.910 129.225 ;
        RECT 83.090 128.715 83.370 129.045 ;
        RECT 83.600 128.715 83.815 129.225 ;
        RECT 81.640 128.375 81.815 128.425 ;
        RECT 79.745 127.765 80.495 128.285 ;
        RECT 81.135 127.985 81.470 128.255 ;
        RECT 81.640 127.825 81.810 128.375 ;
        RECT 81.980 127.985 82.315 128.235 ;
        RECT 82.565 127.985 82.920 128.545 ;
        RECT 76.435 127.355 78.655 127.525 ;
        RECT 76.095 127.185 76.265 127.355 ;
        RECT 75.625 126.675 75.925 127.185 ;
        RECT 76.095 127.015 76.475 127.185 ;
        RECT 77.055 126.675 77.685 127.185 ;
        RECT 77.855 126.845 78.185 127.355 ;
        RECT 78.355 126.675 78.655 127.185 ;
        RECT 78.825 126.675 80.495 127.765 ;
        RECT 81.125 126.675 81.405 127.815 ;
        RECT 81.575 126.845 81.905 127.825 ;
        RECT 83.090 127.815 83.260 128.715 ;
        RECT 83.430 127.985 83.695 128.545 ;
        RECT 83.985 128.485 84.600 129.055 ;
        RECT 83.945 127.815 84.115 128.315 ;
        RECT 82.075 126.675 82.335 127.815 ;
        RECT 82.690 127.645 84.115 127.815 ;
        RECT 82.690 127.470 83.080 127.645 ;
        RECT 83.565 126.675 83.895 127.475 ;
        RECT 84.285 127.465 84.600 128.485 ;
        RECT 84.065 126.845 84.600 127.465 ;
        RECT 85.265 128.550 85.540 128.895 ;
        RECT 85.730 128.825 86.105 129.225 ;
        RECT 86.275 128.655 86.445 129.005 ;
        RECT 86.615 128.825 86.945 129.225 ;
        RECT 87.115 128.655 87.375 129.055 ;
        RECT 85.265 127.815 85.435 128.550 ;
        RECT 85.710 128.485 87.375 128.655 ;
        RECT 85.710 128.315 85.880 128.485 ;
        RECT 87.555 128.405 87.885 128.825 ;
        RECT 88.055 128.405 88.315 129.225 ;
        RECT 88.485 128.500 88.775 129.225 ;
        RECT 88.955 128.495 89.255 129.225 ;
        RECT 87.555 128.315 87.805 128.405 ;
        RECT 89.435 128.315 89.665 128.935 ;
        RECT 89.865 128.665 90.090 129.045 ;
        RECT 90.260 128.835 90.590 129.225 ;
        RECT 90.955 128.710 91.125 129.225 ;
        RECT 89.865 128.485 90.195 128.665 ;
        RECT 85.605 127.985 85.880 128.315 ;
        RECT 86.050 127.985 86.875 128.315 ;
        RECT 87.090 127.985 87.805 128.315 ;
        RECT 87.975 127.985 88.310 128.235 ;
        RECT 88.960 127.985 89.255 128.315 ;
        RECT 89.435 127.985 89.850 128.315 ;
        RECT 85.710 127.815 85.880 127.985 ;
        RECT 85.265 126.845 85.540 127.815 ;
        RECT 85.710 127.645 86.370 127.815 ;
        RECT 86.630 127.695 86.875 127.985 ;
        RECT 86.200 127.525 86.370 127.645 ;
        RECT 87.045 127.525 87.375 127.815 ;
        RECT 85.750 126.675 86.030 127.475 ;
        RECT 86.200 127.355 87.375 127.525 ;
        RECT 87.635 127.425 87.805 127.985 ;
        RECT 86.200 126.855 87.815 127.185 ;
        RECT 88.055 126.675 88.315 127.815 ;
        RECT 88.485 126.675 88.775 127.840 ;
        RECT 90.020 127.815 90.195 128.485 ;
        RECT 90.365 127.985 90.605 128.635 ;
        RECT 91.295 128.570 91.625 129.005 ;
        RECT 91.795 128.615 91.965 129.225 ;
        RECT 91.245 128.485 91.625 128.570 ;
        RECT 92.135 128.485 92.465 129.010 ;
        RECT 92.725 128.695 92.935 129.225 ;
        RECT 93.210 128.775 93.995 128.945 ;
        RECT 94.165 128.775 94.570 128.945 ;
        RECT 91.245 128.445 91.470 128.485 ;
        RECT 91.245 127.865 91.415 128.445 ;
        RECT 92.135 128.315 92.335 128.485 ;
        RECT 93.210 128.315 93.380 128.775 ;
        RECT 91.585 127.985 92.335 128.315 ;
        RECT 92.505 127.985 93.380 128.315 ;
        RECT 91.245 127.815 91.460 127.865 ;
        RECT 88.955 127.455 89.850 127.785 ;
        RECT 90.020 127.625 90.605 127.815 ;
        RECT 91.245 127.735 91.635 127.815 ;
        RECT 88.955 127.285 90.160 127.455 ;
        RECT 88.955 126.855 89.285 127.285 ;
        RECT 89.465 126.675 89.660 127.115 ;
        RECT 89.830 126.855 90.160 127.285 ;
        RECT 90.330 126.855 90.605 127.625 ;
        RECT 90.965 126.675 91.135 127.590 ;
        RECT 91.305 126.890 91.635 127.735 ;
        RECT 92.145 127.780 92.335 127.985 ;
        RECT 91.805 126.675 91.975 127.685 ;
        RECT 92.145 127.405 93.040 127.780 ;
        RECT 92.145 126.845 92.485 127.405 ;
        RECT 92.715 126.675 93.030 127.175 ;
        RECT 93.210 127.145 93.380 127.985 ;
        RECT 93.550 128.275 94.015 128.605 ;
        RECT 94.400 128.545 94.570 128.775 ;
        RECT 94.750 128.725 95.120 129.225 ;
        RECT 95.440 128.775 96.115 128.945 ;
        RECT 96.310 128.775 96.645 128.945 ;
        RECT 93.550 127.315 93.870 128.275 ;
        RECT 94.400 128.245 95.230 128.545 ;
        RECT 94.040 127.345 94.230 128.065 ;
        RECT 94.400 127.175 94.570 128.245 ;
        RECT 95.030 128.215 95.230 128.245 ;
        RECT 94.740 127.995 94.910 128.065 ;
        RECT 95.440 127.995 95.610 128.775 ;
        RECT 96.475 128.635 96.645 128.775 ;
        RECT 96.815 128.765 97.065 129.225 ;
        RECT 94.740 127.825 95.610 127.995 ;
        RECT 95.780 128.355 96.305 128.575 ;
        RECT 96.475 128.505 96.700 128.635 ;
        RECT 94.740 127.735 95.250 127.825 ;
        RECT 93.210 126.975 94.095 127.145 ;
        RECT 94.320 126.845 94.570 127.175 ;
        RECT 94.740 126.675 94.910 127.475 ;
        RECT 95.080 127.120 95.250 127.735 ;
        RECT 95.780 127.655 95.950 128.355 ;
        RECT 95.420 127.290 95.950 127.655 ;
        RECT 96.120 127.590 96.360 128.185 ;
        RECT 96.530 127.400 96.700 128.505 ;
        RECT 96.870 127.645 97.150 128.595 ;
        RECT 96.395 127.270 96.700 127.400 ;
        RECT 95.080 126.950 96.185 127.120 ;
        RECT 96.395 126.845 96.645 127.270 ;
        RECT 96.815 126.675 97.080 127.135 ;
        RECT 97.320 126.845 97.505 128.965 ;
        RECT 97.675 128.845 98.005 129.225 ;
        RECT 98.175 128.675 98.345 128.965 ;
        RECT 98.605 128.680 103.950 129.225 ;
        RECT 104.125 128.680 109.470 129.225 ;
        RECT 97.680 128.505 98.345 128.675 ;
        RECT 97.680 127.515 97.910 128.505 ;
        RECT 98.080 127.685 98.430 128.335 ;
        RECT 100.190 127.850 100.530 128.680 ;
        RECT 97.680 127.345 98.345 127.515 ;
        RECT 97.675 126.675 98.005 127.175 ;
        RECT 98.175 126.845 98.345 127.345 ;
        RECT 102.010 127.110 102.360 128.360 ;
        RECT 105.710 127.850 106.050 128.680 ;
        RECT 109.645 128.455 113.155 129.225 ;
        RECT 114.245 128.500 114.535 129.225 ;
        RECT 114.705 128.680 120.050 129.225 ;
        RECT 120.225 128.680 125.570 129.225 ;
        RECT 125.745 128.680 131.090 129.225 ;
        RECT 131.265 128.680 136.610 129.225 ;
        RECT 107.530 127.110 107.880 128.360 ;
        RECT 109.645 127.935 111.295 128.455 ;
        RECT 111.465 127.765 113.155 128.285 ;
        RECT 116.290 127.850 116.630 128.680 ;
        RECT 98.605 126.675 103.950 127.110 ;
        RECT 104.125 126.675 109.470 127.110 ;
        RECT 109.645 126.675 113.155 127.765 ;
        RECT 114.245 126.675 114.535 127.840 ;
        RECT 118.110 127.110 118.460 128.360 ;
        RECT 121.810 127.850 122.150 128.680 ;
        RECT 123.630 127.110 123.980 128.360 ;
        RECT 127.330 127.850 127.670 128.680 ;
        RECT 129.150 127.110 129.500 128.360 ;
        RECT 132.850 127.850 133.190 128.680 ;
        RECT 136.785 128.455 139.375 129.225 ;
        RECT 140.005 128.500 140.295 129.225 ;
        RECT 140.465 128.680 145.810 129.225 ;
        RECT 134.670 127.110 135.020 128.360 ;
        RECT 136.785 127.935 137.995 128.455 ;
        RECT 138.165 127.765 139.375 128.285 ;
        RECT 142.050 127.850 142.390 128.680 ;
        RECT 145.985 128.455 148.575 129.225 ;
        RECT 149.205 128.475 150.415 129.225 ;
        RECT 114.705 126.675 120.050 127.110 ;
        RECT 120.225 126.675 125.570 127.110 ;
        RECT 125.745 126.675 131.090 127.110 ;
        RECT 131.265 126.675 136.610 127.110 ;
        RECT 136.785 126.675 139.375 127.765 ;
        RECT 140.005 126.675 140.295 127.840 ;
        RECT 143.870 127.110 144.220 128.360 ;
        RECT 145.985 127.935 147.195 128.455 ;
        RECT 147.365 127.765 148.575 128.285 ;
        RECT 140.465 126.675 145.810 127.110 ;
        RECT 145.985 126.675 148.575 127.765 ;
        RECT 149.205 127.765 149.725 128.305 ;
        RECT 149.895 127.935 150.415 128.475 ;
        RECT 149.205 126.675 150.415 127.765 ;
        RECT 11.120 126.505 150.500 126.675 ;
        RECT 11.205 125.415 12.415 126.505 ;
        RECT 12.585 126.070 17.930 126.505 ;
        RECT 18.105 126.070 23.450 126.505 ;
        RECT 11.205 124.705 11.725 125.245 ;
        RECT 11.895 124.875 12.415 125.415 ;
        RECT 11.205 123.955 12.415 124.705 ;
        RECT 14.170 124.500 14.510 125.330 ;
        RECT 15.990 124.820 16.340 126.070 ;
        RECT 19.690 124.500 20.030 125.330 ;
        RECT 21.510 124.820 21.860 126.070 ;
        RECT 24.085 125.340 24.375 126.505 ;
        RECT 24.545 126.070 29.890 126.505 ;
        RECT 30.065 126.070 35.410 126.505 ;
        RECT 12.585 123.955 17.930 124.500 ;
        RECT 18.105 123.955 23.450 124.500 ;
        RECT 24.085 123.955 24.375 124.680 ;
        RECT 26.130 124.500 26.470 125.330 ;
        RECT 27.950 124.820 28.300 126.070 ;
        RECT 31.650 124.500 31.990 125.330 ;
        RECT 33.470 124.820 33.820 126.070 ;
        RECT 35.585 125.415 39.095 126.505 ;
        RECT 39.445 125.590 39.615 126.505 ;
        RECT 39.785 125.445 40.115 126.290 ;
        RECT 40.285 125.495 40.455 126.505 ;
        RECT 40.625 125.775 40.965 126.335 ;
        RECT 41.195 126.005 41.510 126.505 ;
        RECT 41.690 126.035 42.575 126.205 ;
        RECT 35.585 124.725 37.235 125.245 ;
        RECT 37.405 124.895 39.095 125.415 ;
        RECT 39.725 125.365 40.115 125.445 ;
        RECT 40.625 125.400 41.520 125.775 ;
        RECT 39.725 125.315 39.940 125.365 ;
        RECT 39.725 124.735 39.895 125.315 ;
        RECT 40.625 125.195 40.815 125.400 ;
        RECT 41.690 125.195 41.860 126.035 ;
        RECT 42.800 126.005 43.050 126.335 ;
        RECT 40.065 124.865 40.815 125.195 ;
        RECT 40.985 124.865 41.860 125.195 ;
        RECT 24.545 123.955 29.890 124.500 ;
        RECT 30.065 123.955 35.410 124.500 ;
        RECT 35.585 123.955 39.095 124.725 ;
        RECT 39.725 124.695 39.950 124.735 ;
        RECT 40.615 124.695 40.815 124.865 ;
        RECT 39.725 124.610 40.105 124.695 ;
        RECT 39.435 123.955 39.605 124.470 ;
        RECT 39.775 124.175 40.105 124.610 ;
        RECT 40.275 123.955 40.445 124.565 ;
        RECT 40.615 124.170 40.945 124.695 ;
        RECT 41.205 123.955 41.415 124.485 ;
        RECT 41.690 124.405 41.860 124.865 ;
        RECT 42.030 124.905 42.350 125.865 ;
        RECT 42.520 125.115 42.710 125.835 ;
        RECT 42.880 124.935 43.050 126.005 ;
        RECT 43.220 125.705 43.390 126.505 ;
        RECT 43.560 126.060 44.665 126.230 ;
        RECT 43.560 125.445 43.730 126.060 ;
        RECT 44.875 125.910 45.125 126.335 ;
        RECT 45.295 126.045 45.560 126.505 ;
        RECT 43.900 125.525 44.430 125.890 ;
        RECT 44.875 125.780 45.180 125.910 ;
        RECT 43.220 125.355 43.730 125.445 ;
        RECT 43.220 125.185 44.090 125.355 ;
        RECT 43.220 125.115 43.390 125.185 ;
        RECT 43.510 124.935 43.710 124.965 ;
        RECT 42.030 124.575 42.495 124.905 ;
        RECT 42.880 124.635 43.710 124.935 ;
        RECT 42.880 124.405 43.050 124.635 ;
        RECT 41.690 124.235 42.475 124.405 ;
        RECT 42.645 124.235 43.050 124.405 ;
        RECT 43.230 123.955 43.600 124.455 ;
        RECT 43.920 124.405 44.090 125.185 ;
        RECT 44.260 124.825 44.430 125.525 ;
        RECT 44.600 124.995 44.840 125.590 ;
        RECT 44.260 124.605 44.785 124.825 ;
        RECT 45.010 124.675 45.180 125.780 ;
        RECT 44.955 124.545 45.180 124.675 ;
        RECT 45.350 124.585 45.630 125.535 ;
        RECT 44.955 124.405 45.125 124.545 ;
        RECT 43.920 124.235 44.595 124.405 ;
        RECT 44.790 124.235 45.125 124.405 ;
        RECT 45.295 123.955 45.545 124.415 ;
        RECT 45.800 124.215 45.985 126.335 ;
        RECT 46.155 126.005 46.485 126.505 ;
        RECT 46.655 125.835 46.825 126.335 ;
        RECT 46.160 125.665 46.825 125.835 ;
        RECT 46.160 124.675 46.390 125.665 ;
        RECT 46.560 124.845 46.910 125.495 ;
        RECT 47.085 125.415 49.675 126.505 ;
        RECT 47.085 124.725 48.295 125.245 ;
        RECT 48.465 124.895 49.675 125.415 ;
        RECT 49.845 125.340 50.135 126.505 ;
        RECT 50.305 126.070 55.650 126.505 ;
        RECT 46.160 124.505 46.825 124.675 ;
        RECT 46.155 123.955 46.485 124.335 ;
        RECT 46.655 124.215 46.825 124.505 ;
        RECT 47.085 123.955 49.675 124.725 ;
        RECT 49.845 123.955 50.135 124.680 ;
        RECT 51.890 124.500 52.230 125.330 ;
        RECT 53.710 124.820 54.060 126.070 ;
        RECT 55.825 125.415 57.495 126.505 ;
        RECT 57.755 125.835 57.925 126.335 ;
        RECT 58.095 126.005 58.425 126.505 ;
        RECT 57.755 125.665 58.420 125.835 ;
        RECT 55.825 124.725 56.575 125.245 ;
        RECT 56.745 124.895 57.495 125.415 ;
        RECT 57.670 124.845 58.020 125.495 ;
        RECT 50.305 123.955 55.650 124.500 ;
        RECT 55.825 123.955 57.495 124.725 ;
        RECT 58.190 124.675 58.420 125.665 ;
        RECT 57.755 124.505 58.420 124.675 ;
        RECT 57.755 124.215 57.925 124.505 ;
        RECT 58.095 123.955 58.425 124.335 ;
        RECT 58.595 124.215 58.780 126.335 ;
        RECT 59.020 126.045 59.285 126.505 ;
        RECT 59.455 125.910 59.705 126.335 ;
        RECT 59.915 126.060 61.020 126.230 ;
        RECT 59.400 125.780 59.705 125.910 ;
        RECT 58.950 124.585 59.230 125.535 ;
        RECT 59.400 124.675 59.570 125.780 ;
        RECT 59.740 124.995 59.980 125.590 ;
        RECT 60.150 125.525 60.680 125.890 ;
        RECT 60.150 124.825 60.320 125.525 ;
        RECT 60.850 125.445 61.020 126.060 ;
        RECT 61.190 125.705 61.360 126.505 ;
        RECT 61.530 126.005 61.780 126.335 ;
        RECT 62.005 126.035 62.890 126.205 ;
        RECT 60.850 125.355 61.360 125.445 ;
        RECT 59.400 124.545 59.625 124.675 ;
        RECT 59.795 124.605 60.320 124.825 ;
        RECT 60.490 125.185 61.360 125.355 ;
        RECT 59.035 123.955 59.285 124.415 ;
        RECT 59.455 124.405 59.625 124.545 ;
        RECT 60.490 124.405 60.660 125.185 ;
        RECT 61.190 125.115 61.360 125.185 ;
        RECT 60.870 124.935 61.070 124.965 ;
        RECT 61.530 124.935 61.700 126.005 ;
        RECT 61.870 125.115 62.060 125.835 ;
        RECT 60.870 124.635 61.700 124.935 ;
        RECT 62.230 124.905 62.550 125.865 ;
        RECT 59.455 124.235 59.790 124.405 ;
        RECT 59.985 124.235 60.660 124.405 ;
        RECT 60.980 123.955 61.350 124.455 ;
        RECT 61.530 124.405 61.700 124.635 ;
        RECT 62.085 124.575 62.550 124.905 ;
        RECT 62.720 125.195 62.890 126.035 ;
        RECT 63.070 126.005 63.385 126.505 ;
        RECT 63.615 125.775 63.955 126.335 ;
        RECT 63.060 125.400 63.955 125.775 ;
        RECT 64.125 125.495 64.295 126.505 ;
        RECT 63.765 125.195 63.955 125.400 ;
        RECT 64.465 125.445 64.795 126.290 ;
        RECT 64.965 125.590 65.135 126.505 ;
        RECT 65.575 125.575 65.745 126.335 ;
        RECT 65.925 125.745 66.255 126.505 ;
        RECT 64.465 125.365 64.855 125.445 ;
        RECT 65.575 125.405 66.240 125.575 ;
        RECT 66.425 125.430 66.695 126.335 ;
        RECT 66.865 126.070 72.210 126.505 ;
        RECT 64.640 125.315 64.855 125.365 ;
        RECT 62.720 124.865 63.595 125.195 ;
        RECT 63.765 124.865 64.515 125.195 ;
        RECT 62.720 124.405 62.890 124.865 ;
        RECT 63.765 124.695 63.965 124.865 ;
        RECT 64.685 124.735 64.855 125.315 ;
        RECT 66.070 125.260 66.240 125.405 ;
        RECT 65.505 124.855 65.835 125.225 ;
        RECT 66.070 124.930 66.355 125.260 ;
        RECT 64.630 124.695 64.855 124.735 ;
        RECT 61.530 124.235 61.935 124.405 ;
        RECT 62.105 124.235 62.890 124.405 ;
        RECT 63.165 123.955 63.375 124.485 ;
        RECT 63.635 124.170 63.965 124.695 ;
        RECT 64.475 124.610 64.855 124.695 ;
        RECT 66.070 124.675 66.240 124.930 ;
        RECT 64.135 123.955 64.305 124.565 ;
        RECT 64.475 124.175 64.805 124.610 ;
        RECT 65.575 124.505 66.240 124.675 ;
        RECT 66.525 124.630 66.695 125.430 ;
        RECT 64.975 123.955 65.145 124.470 ;
        RECT 65.575 124.125 65.745 124.505 ;
        RECT 65.925 123.955 66.255 124.335 ;
        RECT 66.435 124.125 66.695 124.630 ;
        RECT 68.450 124.500 68.790 125.330 ;
        RECT 70.270 124.820 70.620 126.070 ;
        RECT 72.385 125.415 74.975 126.505 ;
        RECT 72.385 124.725 73.595 125.245 ;
        RECT 73.765 124.895 74.975 125.415 ;
        RECT 75.605 125.340 75.895 126.505 ;
        RECT 76.065 126.070 81.410 126.505 ;
        RECT 81.585 126.070 86.930 126.505 ;
        RECT 66.865 123.955 72.210 124.500 ;
        RECT 72.385 123.955 74.975 124.725 ;
        RECT 75.605 123.955 75.895 124.680 ;
        RECT 77.650 124.500 77.990 125.330 ;
        RECT 79.470 124.820 79.820 126.070 ;
        RECT 83.170 124.500 83.510 125.330 ;
        RECT 84.990 124.820 85.340 126.070 ;
        RECT 87.105 125.415 90.615 126.505 ;
        RECT 91.820 125.875 92.105 126.335 ;
        RECT 92.275 126.045 92.545 126.505 ;
        RECT 91.820 125.655 92.775 125.875 ;
        RECT 87.105 124.725 88.755 125.245 ;
        RECT 88.925 124.895 90.615 125.415 ;
        RECT 91.705 124.925 92.395 125.485 ;
        RECT 92.565 124.755 92.775 125.655 ;
        RECT 76.065 123.955 81.410 124.500 ;
        RECT 81.585 123.955 86.930 124.500 ;
        RECT 87.105 123.955 90.615 124.725 ;
        RECT 91.820 124.585 92.775 124.755 ;
        RECT 92.945 125.485 93.345 126.335 ;
        RECT 93.535 125.875 93.815 126.335 ;
        RECT 94.335 126.045 94.660 126.505 ;
        RECT 93.535 125.655 94.660 125.875 ;
        RECT 92.945 124.925 94.040 125.485 ;
        RECT 94.210 125.195 94.660 125.655 ;
        RECT 94.830 125.365 95.215 126.335 ;
        RECT 95.385 125.365 95.645 126.505 ;
        RECT 91.820 124.125 92.105 124.585 ;
        RECT 92.275 123.955 92.545 124.415 ;
        RECT 92.945 124.125 93.345 124.925 ;
        RECT 94.210 124.865 94.765 125.195 ;
        RECT 94.210 124.755 94.660 124.865 ;
        RECT 93.535 124.585 94.660 124.755 ;
        RECT 94.935 124.695 95.215 125.365 ;
        RECT 95.815 125.355 96.145 126.335 ;
        RECT 96.315 125.365 96.595 126.505 ;
        RECT 96.765 125.415 100.275 126.505 ;
        RECT 95.405 124.945 95.740 125.195 ;
        RECT 95.910 124.755 96.080 125.355 ;
        RECT 96.250 124.925 96.585 125.195 ;
        RECT 93.535 124.125 93.815 124.585 ;
        RECT 94.335 123.955 94.660 124.415 ;
        RECT 94.830 124.125 95.215 124.695 ;
        RECT 95.385 124.125 96.080 124.755 ;
        RECT 96.285 123.955 96.595 124.755 ;
        RECT 96.765 124.725 98.415 125.245 ;
        RECT 98.585 124.895 100.275 125.415 ;
        RECT 101.365 125.340 101.655 126.505 ;
        RECT 101.825 126.070 107.170 126.505 ;
        RECT 107.345 126.070 112.690 126.505 ;
        RECT 112.865 126.070 118.210 126.505 ;
        RECT 118.385 126.070 123.730 126.505 ;
        RECT 96.765 123.955 100.275 124.725 ;
        RECT 101.365 123.955 101.655 124.680 ;
        RECT 103.410 124.500 103.750 125.330 ;
        RECT 105.230 124.820 105.580 126.070 ;
        RECT 108.930 124.500 109.270 125.330 ;
        RECT 110.750 124.820 111.100 126.070 ;
        RECT 114.450 124.500 114.790 125.330 ;
        RECT 116.270 124.820 116.620 126.070 ;
        RECT 119.970 124.500 120.310 125.330 ;
        RECT 121.790 124.820 122.140 126.070 ;
        RECT 123.905 125.415 126.495 126.505 ;
        RECT 123.905 124.725 125.115 125.245 ;
        RECT 125.285 124.895 126.495 125.415 ;
        RECT 127.125 125.340 127.415 126.505 ;
        RECT 127.585 126.070 132.930 126.505 ;
        RECT 133.105 126.070 138.450 126.505 ;
        RECT 138.625 126.070 143.970 126.505 ;
        RECT 101.825 123.955 107.170 124.500 ;
        RECT 107.345 123.955 112.690 124.500 ;
        RECT 112.865 123.955 118.210 124.500 ;
        RECT 118.385 123.955 123.730 124.500 ;
        RECT 123.905 123.955 126.495 124.725 ;
        RECT 127.125 123.955 127.415 124.680 ;
        RECT 129.170 124.500 129.510 125.330 ;
        RECT 130.990 124.820 131.340 126.070 ;
        RECT 134.690 124.500 135.030 125.330 ;
        RECT 136.510 124.820 136.860 126.070 ;
        RECT 140.210 124.500 140.550 125.330 ;
        RECT 142.030 124.820 142.380 126.070 ;
        RECT 144.145 125.415 147.655 126.505 ;
        RECT 147.825 125.415 149.035 126.505 ;
        RECT 144.145 124.725 145.795 125.245 ;
        RECT 145.965 124.895 147.655 125.415 ;
        RECT 127.585 123.955 132.930 124.500 ;
        RECT 133.105 123.955 138.450 124.500 ;
        RECT 138.625 123.955 143.970 124.500 ;
        RECT 144.145 123.955 147.655 124.725 ;
        RECT 147.825 124.705 148.345 125.245 ;
        RECT 148.515 124.875 149.035 125.415 ;
        RECT 149.205 125.415 150.415 126.505 ;
        RECT 149.205 124.875 149.725 125.415 ;
        RECT 149.895 124.705 150.415 125.245 ;
        RECT 147.825 123.955 149.035 124.705 ;
        RECT 149.205 123.955 150.415 124.705 ;
        RECT 11.120 123.785 150.500 123.955 ;
        RECT 11.205 123.035 12.415 123.785 ;
        RECT 12.585 123.240 17.930 123.785 ;
        RECT 18.105 123.240 23.450 123.785 ;
        RECT 23.625 123.240 28.970 123.785 ;
        RECT 29.145 123.240 34.490 123.785 ;
        RECT 11.205 122.495 11.725 123.035 ;
        RECT 11.895 122.325 12.415 122.865 ;
        RECT 14.170 122.410 14.510 123.240 ;
        RECT 11.205 121.235 12.415 122.325 ;
        RECT 15.990 121.670 16.340 122.920 ;
        RECT 19.690 122.410 20.030 123.240 ;
        RECT 21.510 121.670 21.860 122.920 ;
        RECT 25.210 122.410 25.550 123.240 ;
        RECT 27.030 121.670 27.380 122.920 ;
        RECT 30.730 122.410 31.070 123.240 ;
        RECT 34.665 123.015 36.335 123.785 ;
        RECT 36.965 123.060 37.255 123.785 ;
        RECT 37.425 123.240 42.770 123.785 ;
        RECT 32.550 121.670 32.900 122.920 ;
        RECT 34.665 122.495 35.415 123.015 ;
        RECT 35.585 122.325 36.335 122.845 ;
        RECT 39.010 122.410 39.350 123.240 ;
        RECT 42.945 123.015 46.455 123.785 ;
        RECT 47.635 123.235 47.805 123.525 ;
        RECT 47.975 123.405 48.305 123.785 ;
        RECT 47.635 123.065 48.300 123.235 ;
        RECT 12.585 121.235 17.930 121.670 ;
        RECT 18.105 121.235 23.450 121.670 ;
        RECT 23.625 121.235 28.970 121.670 ;
        RECT 29.145 121.235 34.490 121.670 ;
        RECT 34.665 121.235 36.335 122.325 ;
        RECT 36.965 121.235 37.255 122.400 ;
        RECT 40.830 121.670 41.180 122.920 ;
        RECT 42.945 122.495 44.595 123.015 ;
        RECT 44.765 122.325 46.455 122.845 ;
        RECT 37.425 121.235 42.770 121.670 ;
        RECT 42.945 121.235 46.455 122.325 ;
        RECT 47.550 122.245 47.900 122.895 ;
        RECT 48.070 122.075 48.300 123.065 ;
        RECT 47.635 121.905 48.300 122.075 ;
        RECT 47.635 121.405 47.805 121.905 ;
        RECT 47.975 121.235 48.305 121.735 ;
        RECT 48.475 121.405 48.660 123.525 ;
        RECT 48.915 123.325 49.165 123.785 ;
        RECT 49.335 123.335 49.670 123.505 ;
        RECT 49.865 123.335 50.540 123.505 ;
        RECT 49.335 123.195 49.505 123.335 ;
        RECT 48.830 122.205 49.110 123.155 ;
        RECT 49.280 123.065 49.505 123.195 ;
        RECT 49.280 121.960 49.450 123.065 ;
        RECT 49.675 122.915 50.200 123.135 ;
        RECT 49.620 122.150 49.860 122.745 ;
        RECT 50.030 122.215 50.200 122.915 ;
        RECT 50.370 122.555 50.540 123.335 ;
        RECT 50.860 123.285 51.230 123.785 ;
        RECT 51.410 123.335 51.815 123.505 ;
        RECT 51.985 123.335 52.770 123.505 ;
        RECT 51.410 123.105 51.580 123.335 ;
        RECT 50.750 122.805 51.580 123.105 ;
        RECT 51.965 122.835 52.430 123.165 ;
        RECT 50.750 122.775 50.950 122.805 ;
        RECT 51.070 122.555 51.240 122.625 ;
        RECT 50.370 122.385 51.240 122.555 ;
        RECT 50.730 122.295 51.240 122.385 ;
        RECT 49.280 121.830 49.585 121.960 ;
        RECT 50.030 121.850 50.560 122.215 ;
        RECT 48.900 121.235 49.165 121.695 ;
        RECT 49.335 121.405 49.585 121.830 ;
        RECT 50.730 121.680 50.900 122.295 ;
        RECT 49.795 121.510 50.900 121.680 ;
        RECT 51.070 121.235 51.240 122.035 ;
        RECT 51.410 121.735 51.580 122.805 ;
        RECT 51.750 121.905 51.940 122.625 ;
        RECT 52.110 121.875 52.430 122.835 ;
        RECT 52.600 122.875 52.770 123.335 ;
        RECT 53.045 123.255 53.255 123.785 ;
        RECT 53.515 123.045 53.845 123.570 ;
        RECT 54.015 123.175 54.185 123.785 ;
        RECT 54.355 123.130 54.685 123.565 ;
        RECT 54.855 123.270 55.025 123.785 ;
        RECT 55.365 123.240 60.710 123.785 ;
        RECT 54.355 123.045 54.735 123.130 ;
        RECT 53.645 122.875 53.845 123.045 ;
        RECT 54.510 123.005 54.735 123.045 ;
        RECT 52.600 122.545 53.475 122.875 ;
        RECT 53.645 122.545 54.395 122.875 ;
        RECT 51.410 121.405 51.660 121.735 ;
        RECT 52.600 121.705 52.770 122.545 ;
        RECT 53.645 122.340 53.835 122.545 ;
        RECT 54.565 122.425 54.735 123.005 ;
        RECT 54.520 122.375 54.735 122.425 ;
        RECT 56.950 122.410 57.290 123.240 ;
        RECT 60.885 123.015 62.555 123.785 ;
        RECT 62.725 123.060 63.015 123.785 ;
        RECT 63.185 123.240 68.530 123.785 ;
        RECT 68.705 123.240 74.050 123.785 ;
        RECT 74.225 123.240 79.570 123.785 ;
        RECT 79.745 123.240 85.090 123.785 ;
        RECT 52.940 121.965 53.835 122.340 ;
        RECT 54.345 122.295 54.735 122.375 ;
        RECT 51.885 121.535 52.770 121.705 ;
        RECT 52.950 121.235 53.265 121.735 ;
        RECT 53.495 121.405 53.835 121.965 ;
        RECT 54.005 121.235 54.175 122.245 ;
        RECT 54.345 121.450 54.675 122.295 ;
        RECT 54.845 121.235 55.015 122.150 ;
        RECT 58.770 121.670 59.120 122.920 ;
        RECT 60.885 122.495 61.635 123.015 ;
        RECT 61.805 122.325 62.555 122.845 ;
        RECT 64.770 122.410 65.110 123.240 ;
        RECT 55.365 121.235 60.710 121.670 ;
        RECT 60.885 121.235 62.555 122.325 ;
        RECT 62.725 121.235 63.015 122.400 ;
        RECT 66.590 121.670 66.940 122.920 ;
        RECT 70.290 122.410 70.630 123.240 ;
        RECT 72.110 121.670 72.460 122.920 ;
        RECT 75.810 122.410 76.150 123.240 ;
        RECT 77.630 121.670 77.980 122.920 ;
        RECT 81.330 122.410 81.670 123.240 ;
        RECT 85.265 123.015 87.855 123.785 ;
        RECT 88.485 123.060 88.775 123.785 ;
        RECT 88.945 123.240 94.290 123.785 ;
        RECT 94.465 123.240 99.810 123.785 ;
        RECT 99.985 123.240 105.330 123.785 ;
        RECT 105.505 123.240 110.850 123.785 ;
        RECT 83.150 121.670 83.500 122.920 ;
        RECT 85.265 122.495 86.475 123.015 ;
        RECT 86.645 122.325 87.855 122.845 ;
        RECT 90.530 122.410 90.870 123.240 ;
        RECT 63.185 121.235 68.530 121.670 ;
        RECT 68.705 121.235 74.050 121.670 ;
        RECT 74.225 121.235 79.570 121.670 ;
        RECT 79.745 121.235 85.090 121.670 ;
        RECT 85.265 121.235 87.855 122.325 ;
        RECT 88.485 121.235 88.775 122.400 ;
        RECT 92.350 121.670 92.700 122.920 ;
        RECT 96.050 122.410 96.390 123.240 ;
        RECT 97.870 121.670 98.220 122.920 ;
        RECT 101.570 122.410 101.910 123.240 ;
        RECT 103.390 121.670 103.740 122.920 ;
        RECT 107.090 122.410 107.430 123.240 ;
        RECT 111.025 123.015 113.615 123.785 ;
        RECT 114.245 123.060 114.535 123.785 ;
        RECT 114.705 123.240 120.050 123.785 ;
        RECT 120.225 123.240 125.570 123.785 ;
        RECT 125.745 123.240 131.090 123.785 ;
        RECT 131.265 123.240 136.610 123.785 ;
        RECT 108.910 121.670 109.260 122.920 ;
        RECT 111.025 122.495 112.235 123.015 ;
        RECT 112.405 122.325 113.615 122.845 ;
        RECT 116.290 122.410 116.630 123.240 ;
        RECT 88.945 121.235 94.290 121.670 ;
        RECT 94.465 121.235 99.810 121.670 ;
        RECT 99.985 121.235 105.330 121.670 ;
        RECT 105.505 121.235 110.850 121.670 ;
        RECT 111.025 121.235 113.615 122.325 ;
        RECT 114.245 121.235 114.535 122.400 ;
        RECT 118.110 121.670 118.460 122.920 ;
        RECT 121.810 122.410 122.150 123.240 ;
        RECT 123.630 121.670 123.980 122.920 ;
        RECT 127.330 122.410 127.670 123.240 ;
        RECT 129.150 121.670 129.500 122.920 ;
        RECT 132.850 122.410 133.190 123.240 ;
        RECT 136.785 123.015 139.375 123.785 ;
        RECT 140.005 123.060 140.295 123.785 ;
        RECT 140.465 123.240 145.810 123.785 ;
        RECT 134.670 121.670 135.020 122.920 ;
        RECT 136.785 122.495 137.995 123.015 ;
        RECT 138.165 122.325 139.375 122.845 ;
        RECT 142.050 122.410 142.390 123.240 ;
        RECT 145.985 123.015 148.575 123.785 ;
        RECT 149.205 123.035 150.415 123.785 ;
        RECT 114.705 121.235 120.050 121.670 ;
        RECT 120.225 121.235 125.570 121.670 ;
        RECT 125.745 121.235 131.090 121.670 ;
        RECT 131.265 121.235 136.610 121.670 ;
        RECT 136.785 121.235 139.375 122.325 ;
        RECT 140.005 121.235 140.295 122.400 ;
        RECT 143.870 121.670 144.220 122.920 ;
        RECT 145.985 122.495 147.195 123.015 ;
        RECT 147.365 122.325 148.575 122.845 ;
        RECT 140.465 121.235 145.810 121.670 ;
        RECT 145.985 121.235 148.575 122.325 ;
        RECT 149.205 122.325 149.725 122.865 ;
        RECT 149.895 122.495 150.415 123.035 ;
        RECT 149.205 121.235 150.415 122.325 ;
        RECT 11.120 121.065 150.500 121.235 ;
        RECT 11.205 119.975 12.415 121.065 ;
        RECT 12.585 120.630 17.930 121.065 ;
        RECT 18.105 120.630 23.450 121.065 ;
        RECT 11.205 119.265 11.725 119.805 ;
        RECT 11.895 119.435 12.415 119.975 ;
        RECT 11.205 118.515 12.415 119.265 ;
        RECT 14.170 119.060 14.510 119.890 ;
        RECT 15.990 119.380 16.340 120.630 ;
        RECT 19.690 119.060 20.030 119.890 ;
        RECT 21.510 119.380 21.860 120.630 ;
        RECT 24.085 119.900 24.375 121.065 ;
        RECT 24.545 120.630 29.890 121.065 ;
        RECT 30.065 120.630 35.410 121.065 ;
        RECT 35.585 120.630 40.930 121.065 ;
        RECT 41.105 120.630 46.450 121.065 ;
        RECT 12.585 118.515 17.930 119.060 ;
        RECT 18.105 118.515 23.450 119.060 ;
        RECT 24.085 118.515 24.375 119.240 ;
        RECT 26.130 119.060 26.470 119.890 ;
        RECT 27.950 119.380 28.300 120.630 ;
        RECT 31.650 119.060 31.990 119.890 ;
        RECT 33.470 119.380 33.820 120.630 ;
        RECT 37.170 119.060 37.510 119.890 ;
        RECT 38.990 119.380 39.340 120.630 ;
        RECT 42.690 119.060 43.030 119.890 ;
        RECT 44.510 119.380 44.860 120.630 ;
        RECT 46.625 119.975 49.215 121.065 ;
        RECT 46.625 119.285 47.835 119.805 ;
        RECT 48.005 119.455 49.215 119.975 ;
        RECT 49.845 119.900 50.135 121.065 ;
        RECT 50.305 120.630 55.650 121.065 ;
        RECT 55.825 120.630 61.170 121.065 ;
        RECT 61.345 120.630 66.690 121.065 ;
        RECT 66.865 120.630 72.210 121.065 ;
        RECT 24.545 118.515 29.890 119.060 ;
        RECT 30.065 118.515 35.410 119.060 ;
        RECT 35.585 118.515 40.930 119.060 ;
        RECT 41.105 118.515 46.450 119.060 ;
        RECT 46.625 118.515 49.215 119.285 ;
        RECT 49.845 118.515 50.135 119.240 ;
        RECT 51.890 119.060 52.230 119.890 ;
        RECT 53.710 119.380 54.060 120.630 ;
        RECT 57.410 119.060 57.750 119.890 ;
        RECT 59.230 119.380 59.580 120.630 ;
        RECT 62.930 119.060 63.270 119.890 ;
        RECT 64.750 119.380 65.100 120.630 ;
        RECT 68.450 119.060 68.790 119.890 ;
        RECT 70.270 119.380 70.620 120.630 ;
        RECT 72.385 119.975 74.975 121.065 ;
        RECT 72.385 119.285 73.595 119.805 ;
        RECT 73.765 119.455 74.975 119.975 ;
        RECT 75.605 119.900 75.895 121.065 ;
        RECT 76.065 120.630 81.410 121.065 ;
        RECT 81.585 120.630 86.930 121.065 ;
        RECT 87.105 120.630 92.450 121.065 ;
        RECT 92.625 120.630 97.970 121.065 ;
        RECT 50.305 118.515 55.650 119.060 ;
        RECT 55.825 118.515 61.170 119.060 ;
        RECT 61.345 118.515 66.690 119.060 ;
        RECT 66.865 118.515 72.210 119.060 ;
        RECT 72.385 118.515 74.975 119.285 ;
        RECT 75.605 118.515 75.895 119.240 ;
        RECT 77.650 119.060 77.990 119.890 ;
        RECT 79.470 119.380 79.820 120.630 ;
        RECT 83.170 119.060 83.510 119.890 ;
        RECT 84.990 119.380 85.340 120.630 ;
        RECT 88.690 119.060 89.030 119.890 ;
        RECT 90.510 119.380 90.860 120.630 ;
        RECT 94.210 119.060 94.550 119.890 ;
        RECT 96.030 119.380 96.380 120.630 ;
        RECT 98.145 119.975 100.735 121.065 ;
        RECT 98.145 119.285 99.355 119.805 ;
        RECT 99.525 119.455 100.735 119.975 ;
        RECT 101.365 119.900 101.655 121.065 ;
        RECT 101.825 120.630 107.170 121.065 ;
        RECT 107.345 120.630 112.690 121.065 ;
        RECT 112.865 120.630 118.210 121.065 ;
        RECT 118.385 120.630 123.730 121.065 ;
        RECT 76.065 118.515 81.410 119.060 ;
        RECT 81.585 118.515 86.930 119.060 ;
        RECT 87.105 118.515 92.450 119.060 ;
        RECT 92.625 118.515 97.970 119.060 ;
        RECT 98.145 118.515 100.735 119.285 ;
        RECT 101.365 118.515 101.655 119.240 ;
        RECT 103.410 119.060 103.750 119.890 ;
        RECT 105.230 119.380 105.580 120.630 ;
        RECT 108.930 119.060 109.270 119.890 ;
        RECT 110.750 119.380 111.100 120.630 ;
        RECT 114.450 119.060 114.790 119.890 ;
        RECT 116.270 119.380 116.620 120.630 ;
        RECT 119.970 119.060 120.310 119.890 ;
        RECT 121.790 119.380 122.140 120.630 ;
        RECT 123.905 119.975 126.495 121.065 ;
        RECT 123.905 119.285 125.115 119.805 ;
        RECT 125.285 119.455 126.495 119.975 ;
        RECT 127.125 119.900 127.415 121.065 ;
        RECT 127.585 120.630 132.930 121.065 ;
        RECT 133.105 120.630 138.450 121.065 ;
        RECT 138.625 120.630 143.970 121.065 ;
        RECT 101.825 118.515 107.170 119.060 ;
        RECT 107.345 118.515 112.690 119.060 ;
        RECT 112.865 118.515 118.210 119.060 ;
        RECT 118.385 118.515 123.730 119.060 ;
        RECT 123.905 118.515 126.495 119.285 ;
        RECT 127.125 118.515 127.415 119.240 ;
        RECT 129.170 119.060 129.510 119.890 ;
        RECT 130.990 119.380 131.340 120.630 ;
        RECT 134.690 119.060 135.030 119.890 ;
        RECT 136.510 119.380 136.860 120.630 ;
        RECT 140.210 119.060 140.550 119.890 ;
        RECT 142.030 119.380 142.380 120.630 ;
        RECT 144.145 119.975 147.655 121.065 ;
        RECT 147.825 119.975 149.035 121.065 ;
        RECT 144.145 119.285 145.795 119.805 ;
        RECT 145.965 119.455 147.655 119.975 ;
        RECT 127.585 118.515 132.930 119.060 ;
        RECT 133.105 118.515 138.450 119.060 ;
        RECT 138.625 118.515 143.970 119.060 ;
        RECT 144.145 118.515 147.655 119.285 ;
        RECT 147.825 119.265 148.345 119.805 ;
        RECT 148.515 119.435 149.035 119.975 ;
        RECT 149.205 119.975 150.415 121.065 ;
        RECT 149.205 119.435 149.725 119.975 ;
        RECT 149.895 119.265 150.415 119.805 ;
        RECT 147.825 118.515 149.035 119.265 ;
        RECT 149.205 118.515 150.415 119.265 ;
        RECT 11.120 118.345 150.500 118.515 ;
        RECT 11.205 117.595 12.415 118.345 ;
        RECT 12.585 117.800 17.930 118.345 ;
        RECT 18.105 117.800 23.450 118.345 ;
        RECT 23.625 117.800 28.970 118.345 ;
        RECT 29.145 117.800 34.490 118.345 ;
        RECT 11.205 117.055 11.725 117.595 ;
        RECT 11.895 116.885 12.415 117.425 ;
        RECT 14.170 116.970 14.510 117.800 ;
        RECT 11.205 115.795 12.415 116.885 ;
        RECT 15.990 116.230 16.340 117.480 ;
        RECT 19.690 116.970 20.030 117.800 ;
        RECT 21.510 116.230 21.860 117.480 ;
        RECT 25.210 116.970 25.550 117.800 ;
        RECT 27.030 116.230 27.380 117.480 ;
        RECT 30.730 116.970 31.070 117.800 ;
        RECT 34.665 117.575 36.335 118.345 ;
        RECT 36.965 117.620 37.255 118.345 ;
        RECT 37.425 117.800 42.770 118.345 ;
        RECT 42.945 117.800 48.290 118.345 ;
        RECT 48.465 117.800 53.810 118.345 ;
        RECT 53.985 117.800 59.330 118.345 ;
        RECT 32.550 116.230 32.900 117.480 ;
        RECT 34.665 117.055 35.415 117.575 ;
        RECT 35.585 116.885 36.335 117.405 ;
        RECT 39.010 116.970 39.350 117.800 ;
        RECT 12.585 115.795 17.930 116.230 ;
        RECT 18.105 115.795 23.450 116.230 ;
        RECT 23.625 115.795 28.970 116.230 ;
        RECT 29.145 115.795 34.490 116.230 ;
        RECT 34.665 115.795 36.335 116.885 ;
        RECT 36.965 115.795 37.255 116.960 ;
        RECT 40.830 116.230 41.180 117.480 ;
        RECT 44.530 116.970 44.870 117.800 ;
        RECT 46.350 116.230 46.700 117.480 ;
        RECT 50.050 116.970 50.390 117.800 ;
        RECT 51.870 116.230 52.220 117.480 ;
        RECT 55.570 116.970 55.910 117.800 ;
        RECT 59.505 117.575 62.095 118.345 ;
        RECT 62.725 117.620 63.015 118.345 ;
        RECT 63.185 117.800 68.530 118.345 ;
        RECT 68.705 117.800 74.050 118.345 ;
        RECT 74.225 117.800 79.570 118.345 ;
        RECT 79.745 117.800 85.090 118.345 ;
        RECT 57.390 116.230 57.740 117.480 ;
        RECT 59.505 117.055 60.715 117.575 ;
        RECT 60.885 116.885 62.095 117.405 ;
        RECT 64.770 116.970 65.110 117.800 ;
        RECT 37.425 115.795 42.770 116.230 ;
        RECT 42.945 115.795 48.290 116.230 ;
        RECT 48.465 115.795 53.810 116.230 ;
        RECT 53.985 115.795 59.330 116.230 ;
        RECT 59.505 115.795 62.095 116.885 ;
        RECT 62.725 115.795 63.015 116.960 ;
        RECT 66.590 116.230 66.940 117.480 ;
        RECT 70.290 116.970 70.630 117.800 ;
        RECT 72.110 116.230 72.460 117.480 ;
        RECT 75.810 116.970 76.150 117.800 ;
        RECT 77.630 116.230 77.980 117.480 ;
        RECT 81.330 116.970 81.670 117.800 ;
        RECT 85.265 117.575 87.855 118.345 ;
        RECT 88.485 117.620 88.775 118.345 ;
        RECT 88.945 117.800 94.290 118.345 ;
        RECT 94.465 117.800 99.810 118.345 ;
        RECT 99.985 117.800 105.330 118.345 ;
        RECT 105.505 117.800 110.850 118.345 ;
        RECT 83.150 116.230 83.500 117.480 ;
        RECT 85.265 117.055 86.475 117.575 ;
        RECT 86.645 116.885 87.855 117.405 ;
        RECT 90.530 116.970 90.870 117.800 ;
        RECT 63.185 115.795 68.530 116.230 ;
        RECT 68.705 115.795 74.050 116.230 ;
        RECT 74.225 115.795 79.570 116.230 ;
        RECT 79.745 115.795 85.090 116.230 ;
        RECT 85.265 115.795 87.855 116.885 ;
        RECT 88.485 115.795 88.775 116.960 ;
        RECT 92.350 116.230 92.700 117.480 ;
        RECT 96.050 116.970 96.390 117.800 ;
        RECT 97.870 116.230 98.220 117.480 ;
        RECT 101.570 116.970 101.910 117.800 ;
        RECT 103.390 116.230 103.740 117.480 ;
        RECT 107.090 116.970 107.430 117.800 ;
        RECT 111.025 117.575 113.615 118.345 ;
        RECT 114.245 117.620 114.535 118.345 ;
        RECT 114.705 117.800 120.050 118.345 ;
        RECT 120.225 117.800 125.570 118.345 ;
        RECT 125.745 117.800 131.090 118.345 ;
        RECT 131.265 117.800 136.610 118.345 ;
        RECT 108.910 116.230 109.260 117.480 ;
        RECT 111.025 117.055 112.235 117.575 ;
        RECT 112.405 116.885 113.615 117.405 ;
        RECT 116.290 116.970 116.630 117.800 ;
        RECT 88.945 115.795 94.290 116.230 ;
        RECT 94.465 115.795 99.810 116.230 ;
        RECT 99.985 115.795 105.330 116.230 ;
        RECT 105.505 115.795 110.850 116.230 ;
        RECT 111.025 115.795 113.615 116.885 ;
        RECT 114.245 115.795 114.535 116.960 ;
        RECT 118.110 116.230 118.460 117.480 ;
        RECT 121.810 116.970 122.150 117.800 ;
        RECT 123.630 116.230 123.980 117.480 ;
        RECT 127.330 116.970 127.670 117.800 ;
        RECT 129.150 116.230 129.500 117.480 ;
        RECT 132.850 116.970 133.190 117.800 ;
        RECT 136.785 117.575 139.375 118.345 ;
        RECT 140.005 117.620 140.295 118.345 ;
        RECT 140.465 117.800 145.810 118.345 ;
        RECT 134.670 116.230 135.020 117.480 ;
        RECT 136.785 117.055 137.995 117.575 ;
        RECT 138.165 116.885 139.375 117.405 ;
        RECT 142.050 116.970 142.390 117.800 ;
        RECT 145.985 117.575 148.575 118.345 ;
        RECT 149.205 117.595 150.415 118.345 ;
        RECT 114.705 115.795 120.050 116.230 ;
        RECT 120.225 115.795 125.570 116.230 ;
        RECT 125.745 115.795 131.090 116.230 ;
        RECT 131.265 115.795 136.610 116.230 ;
        RECT 136.785 115.795 139.375 116.885 ;
        RECT 140.005 115.795 140.295 116.960 ;
        RECT 143.870 116.230 144.220 117.480 ;
        RECT 145.985 117.055 147.195 117.575 ;
        RECT 147.365 116.885 148.575 117.405 ;
        RECT 140.465 115.795 145.810 116.230 ;
        RECT 145.985 115.795 148.575 116.885 ;
        RECT 149.205 116.885 149.725 117.425 ;
        RECT 149.895 117.055 150.415 117.595 ;
        RECT 149.205 115.795 150.415 116.885 ;
        RECT 11.120 115.625 150.500 115.795 ;
        RECT 11.205 114.535 12.415 115.625 ;
        RECT 12.585 115.190 17.930 115.625 ;
        RECT 18.105 115.190 23.450 115.625 ;
        RECT 11.205 113.825 11.725 114.365 ;
        RECT 11.895 113.995 12.415 114.535 ;
        RECT 11.205 113.075 12.415 113.825 ;
        RECT 14.170 113.620 14.510 114.450 ;
        RECT 15.990 113.940 16.340 115.190 ;
        RECT 19.690 113.620 20.030 114.450 ;
        RECT 21.510 113.940 21.860 115.190 ;
        RECT 24.085 114.460 24.375 115.625 ;
        RECT 24.545 115.190 29.890 115.625 ;
        RECT 30.065 115.190 35.410 115.625 ;
        RECT 35.585 115.190 40.930 115.625 ;
        RECT 41.105 115.190 46.450 115.625 ;
        RECT 12.585 113.075 17.930 113.620 ;
        RECT 18.105 113.075 23.450 113.620 ;
        RECT 24.085 113.075 24.375 113.800 ;
        RECT 26.130 113.620 26.470 114.450 ;
        RECT 27.950 113.940 28.300 115.190 ;
        RECT 31.650 113.620 31.990 114.450 ;
        RECT 33.470 113.940 33.820 115.190 ;
        RECT 37.170 113.620 37.510 114.450 ;
        RECT 38.990 113.940 39.340 115.190 ;
        RECT 42.690 113.620 43.030 114.450 ;
        RECT 44.510 113.940 44.860 115.190 ;
        RECT 46.625 114.535 49.215 115.625 ;
        RECT 46.625 113.845 47.835 114.365 ;
        RECT 48.005 114.015 49.215 114.535 ;
        RECT 49.845 114.460 50.135 115.625 ;
        RECT 50.305 115.190 55.650 115.625 ;
        RECT 55.825 115.190 61.170 115.625 ;
        RECT 61.345 115.190 66.690 115.625 ;
        RECT 66.865 115.190 72.210 115.625 ;
        RECT 24.545 113.075 29.890 113.620 ;
        RECT 30.065 113.075 35.410 113.620 ;
        RECT 35.585 113.075 40.930 113.620 ;
        RECT 41.105 113.075 46.450 113.620 ;
        RECT 46.625 113.075 49.215 113.845 ;
        RECT 49.845 113.075 50.135 113.800 ;
        RECT 51.890 113.620 52.230 114.450 ;
        RECT 53.710 113.940 54.060 115.190 ;
        RECT 57.410 113.620 57.750 114.450 ;
        RECT 59.230 113.940 59.580 115.190 ;
        RECT 62.930 113.620 63.270 114.450 ;
        RECT 64.750 113.940 65.100 115.190 ;
        RECT 68.450 113.620 68.790 114.450 ;
        RECT 70.270 113.940 70.620 115.190 ;
        RECT 72.385 114.535 74.975 115.625 ;
        RECT 72.385 113.845 73.595 114.365 ;
        RECT 73.765 114.015 74.975 114.535 ;
        RECT 75.605 114.460 75.895 115.625 ;
        RECT 76.065 115.190 81.410 115.625 ;
        RECT 81.585 115.190 86.930 115.625 ;
        RECT 87.105 115.190 92.450 115.625 ;
        RECT 92.625 115.190 97.970 115.625 ;
        RECT 50.305 113.075 55.650 113.620 ;
        RECT 55.825 113.075 61.170 113.620 ;
        RECT 61.345 113.075 66.690 113.620 ;
        RECT 66.865 113.075 72.210 113.620 ;
        RECT 72.385 113.075 74.975 113.845 ;
        RECT 75.605 113.075 75.895 113.800 ;
        RECT 77.650 113.620 77.990 114.450 ;
        RECT 79.470 113.940 79.820 115.190 ;
        RECT 83.170 113.620 83.510 114.450 ;
        RECT 84.990 113.940 85.340 115.190 ;
        RECT 88.690 113.620 89.030 114.450 ;
        RECT 90.510 113.940 90.860 115.190 ;
        RECT 94.210 113.620 94.550 114.450 ;
        RECT 96.030 113.940 96.380 115.190 ;
        RECT 98.145 114.535 100.735 115.625 ;
        RECT 98.145 113.845 99.355 114.365 ;
        RECT 99.525 114.015 100.735 114.535 ;
        RECT 101.365 114.460 101.655 115.625 ;
        RECT 101.825 115.190 107.170 115.625 ;
        RECT 107.345 115.190 112.690 115.625 ;
        RECT 112.865 115.190 118.210 115.625 ;
        RECT 118.385 115.190 123.730 115.625 ;
        RECT 76.065 113.075 81.410 113.620 ;
        RECT 81.585 113.075 86.930 113.620 ;
        RECT 87.105 113.075 92.450 113.620 ;
        RECT 92.625 113.075 97.970 113.620 ;
        RECT 98.145 113.075 100.735 113.845 ;
        RECT 101.365 113.075 101.655 113.800 ;
        RECT 103.410 113.620 103.750 114.450 ;
        RECT 105.230 113.940 105.580 115.190 ;
        RECT 108.930 113.620 109.270 114.450 ;
        RECT 110.750 113.940 111.100 115.190 ;
        RECT 114.450 113.620 114.790 114.450 ;
        RECT 116.270 113.940 116.620 115.190 ;
        RECT 119.970 113.620 120.310 114.450 ;
        RECT 121.790 113.940 122.140 115.190 ;
        RECT 123.905 114.535 126.495 115.625 ;
        RECT 123.905 113.845 125.115 114.365 ;
        RECT 125.285 114.015 126.495 114.535 ;
        RECT 127.125 114.460 127.415 115.625 ;
        RECT 127.585 115.190 132.930 115.625 ;
        RECT 133.105 115.190 138.450 115.625 ;
        RECT 138.625 115.190 143.970 115.625 ;
        RECT 101.825 113.075 107.170 113.620 ;
        RECT 107.345 113.075 112.690 113.620 ;
        RECT 112.865 113.075 118.210 113.620 ;
        RECT 118.385 113.075 123.730 113.620 ;
        RECT 123.905 113.075 126.495 113.845 ;
        RECT 127.125 113.075 127.415 113.800 ;
        RECT 129.170 113.620 129.510 114.450 ;
        RECT 130.990 113.940 131.340 115.190 ;
        RECT 134.690 113.620 135.030 114.450 ;
        RECT 136.510 113.940 136.860 115.190 ;
        RECT 140.210 113.620 140.550 114.450 ;
        RECT 142.030 113.940 142.380 115.190 ;
        RECT 144.145 114.535 147.655 115.625 ;
        RECT 147.825 114.535 149.035 115.625 ;
        RECT 144.145 113.845 145.795 114.365 ;
        RECT 145.965 114.015 147.655 114.535 ;
        RECT 127.585 113.075 132.930 113.620 ;
        RECT 133.105 113.075 138.450 113.620 ;
        RECT 138.625 113.075 143.970 113.620 ;
        RECT 144.145 113.075 147.655 113.845 ;
        RECT 147.825 113.825 148.345 114.365 ;
        RECT 148.515 113.995 149.035 114.535 ;
        RECT 149.205 114.535 150.415 115.625 ;
        RECT 149.205 113.995 149.725 114.535 ;
        RECT 149.895 113.825 150.415 114.365 ;
        RECT 147.825 113.075 149.035 113.825 ;
        RECT 149.205 113.075 150.415 113.825 ;
        RECT 11.120 112.905 150.500 113.075 ;
        RECT 11.205 112.155 12.415 112.905 ;
        RECT 12.585 112.360 17.930 112.905 ;
        RECT 18.105 112.360 23.450 112.905 ;
        RECT 23.625 112.360 28.970 112.905 ;
        RECT 29.145 112.360 34.490 112.905 ;
        RECT 11.205 111.615 11.725 112.155 ;
        RECT 11.895 111.445 12.415 111.985 ;
        RECT 14.170 111.530 14.510 112.360 ;
        RECT 11.205 110.355 12.415 111.445 ;
        RECT 15.990 110.790 16.340 112.040 ;
        RECT 19.690 111.530 20.030 112.360 ;
        RECT 21.510 110.790 21.860 112.040 ;
        RECT 25.210 111.530 25.550 112.360 ;
        RECT 27.030 110.790 27.380 112.040 ;
        RECT 30.730 111.530 31.070 112.360 ;
        RECT 34.665 112.135 36.335 112.905 ;
        RECT 36.965 112.180 37.255 112.905 ;
        RECT 37.425 112.360 42.770 112.905 ;
        RECT 42.945 112.360 48.290 112.905 ;
        RECT 48.465 112.360 53.810 112.905 ;
        RECT 53.985 112.360 59.330 112.905 ;
        RECT 32.550 110.790 32.900 112.040 ;
        RECT 34.665 111.615 35.415 112.135 ;
        RECT 35.585 111.445 36.335 111.965 ;
        RECT 39.010 111.530 39.350 112.360 ;
        RECT 12.585 110.355 17.930 110.790 ;
        RECT 18.105 110.355 23.450 110.790 ;
        RECT 23.625 110.355 28.970 110.790 ;
        RECT 29.145 110.355 34.490 110.790 ;
        RECT 34.665 110.355 36.335 111.445 ;
        RECT 36.965 110.355 37.255 111.520 ;
        RECT 40.830 110.790 41.180 112.040 ;
        RECT 44.530 111.530 44.870 112.360 ;
        RECT 46.350 110.790 46.700 112.040 ;
        RECT 50.050 111.530 50.390 112.360 ;
        RECT 51.870 110.790 52.220 112.040 ;
        RECT 55.570 111.530 55.910 112.360 ;
        RECT 59.505 112.135 62.095 112.905 ;
        RECT 62.725 112.180 63.015 112.905 ;
        RECT 63.185 112.360 68.530 112.905 ;
        RECT 68.705 112.360 74.050 112.905 ;
        RECT 74.225 112.360 79.570 112.905 ;
        RECT 79.745 112.360 85.090 112.905 ;
        RECT 57.390 110.790 57.740 112.040 ;
        RECT 59.505 111.615 60.715 112.135 ;
        RECT 60.885 111.445 62.095 111.965 ;
        RECT 64.770 111.530 65.110 112.360 ;
        RECT 37.425 110.355 42.770 110.790 ;
        RECT 42.945 110.355 48.290 110.790 ;
        RECT 48.465 110.355 53.810 110.790 ;
        RECT 53.985 110.355 59.330 110.790 ;
        RECT 59.505 110.355 62.095 111.445 ;
        RECT 62.725 110.355 63.015 111.520 ;
        RECT 66.590 110.790 66.940 112.040 ;
        RECT 70.290 111.530 70.630 112.360 ;
        RECT 72.110 110.790 72.460 112.040 ;
        RECT 75.810 111.530 76.150 112.360 ;
        RECT 77.630 110.790 77.980 112.040 ;
        RECT 81.330 111.530 81.670 112.360 ;
        RECT 85.265 112.135 87.855 112.905 ;
        RECT 88.485 112.180 88.775 112.905 ;
        RECT 88.945 112.360 94.290 112.905 ;
        RECT 94.465 112.360 99.810 112.905 ;
        RECT 99.985 112.360 105.330 112.905 ;
        RECT 105.505 112.360 110.850 112.905 ;
        RECT 83.150 110.790 83.500 112.040 ;
        RECT 85.265 111.615 86.475 112.135 ;
        RECT 86.645 111.445 87.855 111.965 ;
        RECT 90.530 111.530 90.870 112.360 ;
        RECT 63.185 110.355 68.530 110.790 ;
        RECT 68.705 110.355 74.050 110.790 ;
        RECT 74.225 110.355 79.570 110.790 ;
        RECT 79.745 110.355 85.090 110.790 ;
        RECT 85.265 110.355 87.855 111.445 ;
        RECT 88.485 110.355 88.775 111.520 ;
        RECT 92.350 110.790 92.700 112.040 ;
        RECT 96.050 111.530 96.390 112.360 ;
        RECT 97.870 110.790 98.220 112.040 ;
        RECT 101.570 111.530 101.910 112.360 ;
        RECT 103.390 110.790 103.740 112.040 ;
        RECT 107.090 111.530 107.430 112.360 ;
        RECT 111.025 112.135 113.615 112.905 ;
        RECT 114.245 112.180 114.535 112.905 ;
        RECT 114.705 112.360 120.050 112.905 ;
        RECT 120.225 112.360 125.570 112.905 ;
        RECT 125.745 112.360 131.090 112.905 ;
        RECT 131.265 112.360 136.610 112.905 ;
        RECT 108.910 110.790 109.260 112.040 ;
        RECT 111.025 111.615 112.235 112.135 ;
        RECT 112.405 111.445 113.615 111.965 ;
        RECT 116.290 111.530 116.630 112.360 ;
        RECT 88.945 110.355 94.290 110.790 ;
        RECT 94.465 110.355 99.810 110.790 ;
        RECT 99.985 110.355 105.330 110.790 ;
        RECT 105.505 110.355 110.850 110.790 ;
        RECT 111.025 110.355 113.615 111.445 ;
        RECT 114.245 110.355 114.535 111.520 ;
        RECT 118.110 110.790 118.460 112.040 ;
        RECT 121.810 111.530 122.150 112.360 ;
        RECT 123.630 110.790 123.980 112.040 ;
        RECT 127.330 111.530 127.670 112.360 ;
        RECT 129.150 110.790 129.500 112.040 ;
        RECT 132.850 111.530 133.190 112.360 ;
        RECT 136.785 112.135 139.375 112.905 ;
        RECT 140.005 112.180 140.295 112.905 ;
        RECT 140.465 112.360 145.810 112.905 ;
        RECT 134.670 110.790 135.020 112.040 ;
        RECT 136.785 111.615 137.995 112.135 ;
        RECT 138.165 111.445 139.375 111.965 ;
        RECT 142.050 111.530 142.390 112.360 ;
        RECT 145.985 112.135 148.575 112.905 ;
        RECT 149.205 112.155 150.415 112.905 ;
        RECT 114.705 110.355 120.050 110.790 ;
        RECT 120.225 110.355 125.570 110.790 ;
        RECT 125.745 110.355 131.090 110.790 ;
        RECT 131.265 110.355 136.610 110.790 ;
        RECT 136.785 110.355 139.375 111.445 ;
        RECT 140.005 110.355 140.295 111.520 ;
        RECT 143.870 110.790 144.220 112.040 ;
        RECT 145.985 111.615 147.195 112.135 ;
        RECT 147.365 111.445 148.575 111.965 ;
        RECT 140.465 110.355 145.810 110.790 ;
        RECT 145.985 110.355 148.575 111.445 ;
        RECT 149.205 111.445 149.725 111.985 ;
        RECT 149.895 111.615 150.415 112.155 ;
        RECT 149.205 110.355 150.415 111.445 ;
        RECT 11.120 110.185 150.500 110.355 ;
        RECT 11.205 109.095 12.415 110.185 ;
        RECT 12.585 109.750 17.930 110.185 ;
        RECT 18.105 109.750 23.450 110.185 ;
        RECT 11.205 108.385 11.725 108.925 ;
        RECT 11.895 108.555 12.415 109.095 ;
        RECT 11.205 107.635 12.415 108.385 ;
        RECT 14.170 108.180 14.510 109.010 ;
        RECT 15.990 108.500 16.340 109.750 ;
        RECT 19.690 108.180 20.030 109.010 ;
        RECT 21.510 108.500 21.860 109.750 ;
        RECT 24.085 109.020 24.375 110.185 ;
        RECT 24.545 109.750 29.890 110.185 ;
        RECT 30.065 109.750 35.410 110.185 ;
        RECT 35.585 109.750 40.930 110.185 ;
        RECT 41.105 109.750 46.450 110.185 ;
        RECT 12.585 107.635 17.930 108.180 ;
        RECT 18.105 107.635 23.450 108.180 ;
        RECT 24.085 107.635 24.375 108.360 ;
        RECT 26.130 108.180 26.470 109.010 ;
        RECT 27.950 108.500 28.300 109.750 ;
        RECT 31.650 108.180 31.990 109.010 ;
        RECT 33.470 108.500 33.820 109.750 ;
        RECT 37.170 108.180 37.510 109.010 ;
        RECT 38.990 108.500 39.340 109.750 ;
        RECT 42.690 108.180 43.030 109.010 ;
        RECT 44.510 108.500 44.860 109.750 ;
        RECT 46.625 109.095 49.215 110.185 ;
        RECT 46.625 108.405 47.835 108.925 ;
        RECT 48.005 108.575 49.215 109.095 ;
        RECT 49.845 109.020 50.135 110.185 ;
        RECT 50.305 109.750 55.650 110.185 ;
        RECT 55.825 109.750 61.170 110.185 ;
        RECT 61.345 109.750 66.690 110.185 ;
        RECT 66.865 109.750 72.210 110.185 ;
        RECT 24.545 107.635 29.890 108.180 ;
        RECT 30.065 107.635 35.410 108.180 ;
        RECT 35.585 107.635 40.930 108.180 ;
        RECT 41.105 107.635 46.450 108.180 ;
        RECT 46.625 107.635 49.215 108.405 ;
        RECT 49.845 107.635 50.135 108.360 ;
        RECT 51.890 108.180 52.230 109.010 ;
        RECT 53.710 108.500 54.060 109.750 ;
        RECT 57.410 108.180 57.750 109.010 ;
        RECT 59.230 108.500 59.580 109.750 ;
        RECT 62.930 108.180 63.270 109.010 ;
        RECT 64.750 108.500 65.100 109.750 ;
        RECT 68.450 108.180 68.790 109.010 ;
        RECT 70.270 108.500 70.620 109.750 ;
        RECT 72.385 109.095 74.975 110.185 ;
        RECT 72.385 108.405 73.595 108.925 ;
        RECT 73.765 108.575 74.975 109.095 ;
        RECT 75.605 109.020 75.895 110.185 ;
        RECT 76.065 109.750 81.410 110.185 ;
        RECT 81.585 109.750 86.930 110.185 ;
        RECT 87.105 109.750 92.450 110.185 ;
        RECT 92.625 109.750 97.970 110.185 ;
        RECT 50.305 107.635 55.650 108.180 ;
        RECT 55.825 107.635 61.170 108.180 ;
        RECT 61.345 107.635 66.690 108.180 ;
        RECT 66.865 107.635 72.210 108.180 ;
        RECT 72.385 107.635 74.975 108.405 ;
        RECT 75.605 107.635 75.895 108.360 ;
        RECT 77.650 108.180 77.990 109.010 ;
        RECT 79.470 108.500 79.820 109.750 ;
        RECT 83.170 108.180 83.510 109.010 ;
        RECT 84.990 108.500 85.340 109.750 ;
        RECT 88.690 108.180 89.030 109.010 ;
        RECT 90.510 108.500 90.860 109.750 ;
        RECT 94.210 108.180 94.550 109.010 ;
        RECT 96.030 108.500 96.380 109.750 ;
        RECT 98.145 109.095 100.735 110.185 ;
        RECT 98.145 108.405 99.355 108.925 ;
        RECT 99.525 108.575 100.735 109.095 ;
        RECT 101.365 109.020 101.655 110.185 ;
        RECT 101.825 109.750 107.170 110.185 ;
        RECT 107.345 109.750 112.690 110.185 ;
        RECT 112.865 109.750 118.210 110.185 ;
        RECT 118.385 109.750 123.730 110.185 ;
        RECT 76.065 107.635 81.410 108.180 ;
        RECT 81.585 107.635 86.930 108.180 ;
        RECT 87.105 107.635 92.450 108.180 ;
        RECT 92.625 107.635 97.970 108.180 ;
        RECT 98.145 107.635 100.735 108.405 ;
        RECT 101.365 107.635 101.655 108.360 ;
        RECT 103.410 108.180 103.750 109.010 ;
        RECT 105.230 108.500 105.580 109.750 ;
        RECT 108.930 108.180 109.270 109.010 ;
        RECT 110.750 108.500 111.100 109.750 ;
        RECT 114.450 108.180 114.790 109.010 ;
        RECT 116.270 108.500 116.620 109.750 ;
        RECT 119.970 108.180 120.310 109.010 ;
        RECT 121.790 108.500 122.140 109.750 ;
        RECT 123.905 109.095 126.495 110.185 ;
        RECT 123.905 108.405 125.115 108.925 ;
        RECT 125.285 108.575 126.495 109.095 ;
        RECT 127.125 109.020 127.415 110.185 ;
        RECT 127.585 109.750 132.930 110.185 ;
        RECT 133.105 109.750 138.450 110.185 ;
        RECT 138.625 109.750 143.970 110.185 ;
        RECT 101.825 107.635 107.170 108.180 ;
        RECT 107.345 107.635 112.690 108.180 ;
        RECT 112.865 107.635 118.210 108.180 ;
        RECT 118.385 107.635 123.730 108.180 ;
        RECT 123.905 107.635 126.495 108.405 ;
        RECT 127.125 107.635 127.415 108.360 ;
        RECT 129.170 108.180 129.510 109.010 ;
        RECT 130.990 108.500 131.340 109.750 ;
        RECT 134.690 108.180 135.030 109.010 ;
        RECT 136.510 108.500 136.860 109.750 ;
        RECT 140.210 108.180 140.550 109.010 ;
        RECT 142.030 108.500 142.380 109.750 ;
        RECT 144.145 109.095 147.655 110.185 ;
        RECT 147.825 109.095 149.035 110.185 ;
        RECT 144.145 108.405 145.795 108.925 ;
        RECT 145.965 108.575 147.655 109.095 ;
        RECT 127.585 107.635 132.930 108.180 ;
        RECT 133.105 107.635 138.450 108.180 ;
        RECT 138.625 107.635 143.970 108.180 ;
        RECT 144.145 107.635 147.655 108.405 ;
        RECT 147.825 108.385 148.345 108.925 ;
        RECT 148.515 108.555 149.035 109.095 ;
        RECT 149.205 109.095 150.415 110.185 ;
        RECT 149.205 108.555 149.725 109.095 ;
        RECT 149.895 108.385 150.415 108.925 ;
        RECT 147.825 107.635 149.035 108.385 ;
        RECT 149.205 107.635 150.415 108.385 ;
        RECT 11.120 107.465 150.500 107.635 ;
        RECT 11.205 106.715 12.415 107.465 ;
        RECT 12.585 106.920 17.930 107.465 ;
        RECT 18.105 106.920 23.450 107.465 ;
        RECT 23.625 106.920 28.970 107.465 ;
        RECT 29.145 106.920 34.490 107.465 ;
        RECT 11.205 106.175 11.725 106.715 ;
        RECT 11.895 106.005 12.415 106.545 ;
        RECT 14.170 106.090 14.510 106.920 ;
        RECT 11.205 104.915 12.415 106.005 ;
        RECT 15.990 105.350 16.340 106.600 ;
        RECT 19.690 106.090 20.030 106.920 ;
        RECT 21.510 105.350 21.860 106.600 ;
        RECT 25.210 106.090 25.550 106.920 ;
        RECT 27.030 105.350 27.380 106.600 ;
        RECT 30.730 106.090 31.070 106.920 ;
        RECT 34.665 106.695 36.335 107.465 ;
        RECT 36.965 106.740 37.255 107.465 ;
        RECT 37.425 106.920 42.770 107.465 ;
        RECT 42.945 106.920 48.290 107.465 ;
        RECT 48.465 106.920 53.810 107.465 ;
        RECT 53.985 106.920 59.330 107.465 ;
        RECT 32.550 105.350 32.900 106.600 ;
        RECT 34.665 106.175 35.415 106.695 ;
        RECT 35.585 106.005 36.335 106.525 ;
        RECT 39.010 106.090 39.350 106.920 ;
        RECT 12.585 104.915 17.930 105.350 ;
        RECT 18.105 104.915 23.450 105.350 ;
        RECT 23.625 104.915 28.970 105.350 ;
        RECT 29.145 104.915 34.490 105.350 ;
        RECT 34.665 104.915 36.335 106.005 ;
        RECT 36.965 104.915 37.255 106.080 ;
        RECT 40.830 105.350 41.180 106.600 ;
        RECT 44.530 106.090 44.870 106.920 ;
        RECT 46.350 105.350 46.700 106.600 ;
        RECT 50.050 106.090 50.390 106.920 ;
        RECT 51.870 105.350 52.220 106.600 ;
        RECT 55.570 106.090 55.910 106.920 ;
        RECT 59.505 106.695 62.095 107.465 ;
        RECT 62.725 106.740 63.015 107.465 ;
        RECT 63.185 106.920 68.530 107.465 ;
        RECT 68.705 106.920 74.050 107.465 ;
        RECT 74.225 106.920 79.570 107.465 ;
        RECT 79.745 106.920 85.090 107.465 ;
        RECT 57.390 105.350 57.740 106.600 ;
        RECT 59.505 106.175 60.715 106.695 ;
        RECT 60.885 106.005 62.095 106.525 ;
        RECT 64.770 106.090 65.110 106.920 ;
        RECT 37.425 104.915 42.770 105.350 ;
        RECT 42.945 104.915 48.290 105.350 ;
        RECT 48.465 104.915 53.810 105.350 ;
        RECT 53.985 104.915 59.330 105.350 ;
        RECT 59.505 104.915 62.095 106.005 ;
        RECT 62.725 104.915 63.015 106.080 ;
        RECT 66.590 105.350 66.940 106.600 ;
        RECT 70.290 106.090 70.630 106.920 ;
        RECT 72.110 105.350 72.460 106.600 ;
        RECT 75.810 106.090 76.150 106.920 ;
        RECT 77.630 105.350 77.980 106.600 ;
        RECT 81.330 106.090 81.670 106.920 ;
        RECT 85.265 106.695 87.855 107.465 ;
        RECT 88.485 106.740 88.775 107.465 ;
        RECT 88.945 106.920 94.290 107.465 ;
        RECT 94.465 106.920 99.810 107.465 ;
        RECT 99.985 106.920 105.330 107.465 ;
        RECT 105.505 106.920 110.850 107.465 ;
        RECT 83.150 105.350 83.500 106.600 ;
        RECT 85.265 106.175 86.475 106.695 ;
        RECT 86.645 106.005 87.855 106.525 ;
        RECT 90.530 106.090 90.870 106.920 ;
        RECT 63.185 104.915 68.530 105.350 ;
        RECT 68.705 104.915 74.050 105.350 ;
        RECT 74.225 104.915 79.570 105.350 ;
        RECT 79.745 104.915 85.090 105.350 ;
        RECT 85.265 104.915 87.855 106.005 ;
        RECT 88.485 104.915 88.775 106.080 ;
        RECT 92.350 105.350 92.700 106.600 ;
        RECT 96.050 106.090 96.390 106.920 ;
        RECT 97.870 105.350 98.220 106.600 ;
        RECT 101.570 106.090 101.910 106.920 ;
        RECT 103.390 105.350 103.740 106.600 ;
        RECT 107.090 106.090 107.430 106.920 ;
        RECT 111.025 106.695 113.615 107.465 ;
        RECT 114.245 106.740 114.535 107.465 ;
        RECT 114.705 106.920 120.050 107.465 ;
        RECT 120.225 106.920 125.570 107.465 ;
        RECT 125.745 106.920 131.090 107.465 ;
        RECT 131.265 106.920 136.610 107.465 ;
        RECT 108.910 105.350 109.260 106.600 ;
        RECT 111.025 106.175 112.235 106.695 ;
        RECT 112.405 106.005 113.615 106.525 ;
        RECT 116.290 106.090 116.630 106.920 ;
        RECT 88.945 104.915 94.290 105.350 ;
        RECT 94.465 104.915 99.810 105.350 ;
        RECT 99.985 104.915 105.330 105.350 ;
        RECT 105.505 104.915 110.850 105.350 ;
        RECT 111.025 104.915 113.615 106.005 ;
        RECT 114.245 104.915 114.535 106.080 ;
        RECT 118.110 105.350 118.460 106.600 ;
        RECT 121.810 106.090 122.150 106.920 ;
        RECT 123.630 105.350 123.980 106.600 ;
        RECT 127.330 106.090 127.670 106.920 ;
        RECT 129.150 105.350 129.500 106.600 ;
        RECT 132.850 106.090 133.190 106.920 ;
        RECT 136.785 106.695 139.375 107.465 ;
        RECT 140.005 106.740 140.295 107.465 ;
        RECT 140.465 106.920 145.810 107.465 ;
        RECT 134.670 105.350 135.020 106.600 ;
        RECT 136.785 106.175 137.995 106.695 ;
        RECT 138.165 106.005 139.375 106.525 ;
        RECT 142.050 106.090 142.390 106.920 ;
        RECT 145.985 106.695 148.575 107.465 ;
        RECT 149.205 106.715 150.415 107.465 ;
        RECT 114.705 104.915 120.050 105.350 ;
        RECT 120.225 104.915 125.570 105.350 ;
        RECT 125.745 104.915 131.090 105.350 ;
        RECT 131.265 104.915 136.610 105.350 ;
        RECT 136.785 104.915 139.375 106.005 ;
        RECT 140.005 104.915 140.295 106.080 ;
        RECT 143.870 105.350 144.220 106.600 ;
        RECT 145.985 106.175 147.195 106.695 ;
        RECT 147.365 106.005 148.575 106.525 ;
        RECT 140.465 104.915 145.810 105.350 ;
        RECT 145.985 104.915 148.575 106.005 ;
        RECT 149.205 106.005 149.725 106.545 ;
        RECT 149.895 106.175 150.415 106.715 ;
        RECT 149.205 104.915 150.415 106.005 ;
        RECT 11.120 104.745 150.500 104.915 ;
        RECT 11.205 103.655 12.415 104.745 ;
        RECT 12.585 104.310 17.930 104.745 ;
        RECT 18.105 104.310 23.450 104.745 ;
        RECT 11.205 102.945 11.725 103.485 ;
        RECT 11.895 103.115 12.415 103.655 ;
        RECT 11.205 102.195 12.415 102.945 ;
        RECT 14.170 102.740 14.510 103.570 ;
        RECT 15.990 103.060 16.340 104.310 ;
        RECT 19.690 102.740 20.030 103.570 ;
        RECT 21.510 103.060 21.860 104.310 ;
        RECT 24.085 103.580 24.375 104.745 ;
        RECT 24.545 104.310 29.890 104.745 ;
        RECT 30.065 104.310 35.410 104.745 ;
        RECT 35.585 104.310 40.930 104.745 ;
        RECT 41.105 104.310 46.450 104.745 ;
        RECT 12.585 102.195 17.930 102.740 ;
        RECT 18.105 102.195 23.450 102.740 ;
        RECT 24.085 102.195 24.375 102.920 ;
        RECT 26.130 102.740 26.470 103.570 ;
        RECT 27.950 103.060 28.300 104.310 ;
        RECT 31.650 102.740 31.990 103.570 ;
        RECT 33.470 103.060 33.820 104.310 ;
        RECT 37.170 102.740 37.510 103.570 ;
        RECT 38.990 103.060 39.340 104.310 ;
        RECT 42.690 102.740 43.030 103.570 ;
        RECT 44.510 103.060 44.860 104.310 ;
        RECT 46.625 103.655 49.215 104.745 ;
        RECT 46.625 102.965 47.835 103.485 ;
        RECT 48.005 103.135 49.215 103.655 ;
        RECT 49.845 103.580 50.135 104.745 ;
        RECT 50.305 104.310 55.650 104.745 ;
        RECT 55.825 104.310 61.170 104.745 ;
        RECT 61.345 104.310 66.690 104.745 ;
        RECT 66.865 104.310 72.210 104.745 ;
        RECT 24.545 102.195 29.890 102.740 ;
        RECT 30.065 102.195 35.410 102.740 ;
        RECT 35.585 102.195 40.930 102.740 ;
        RECT 41.105 102.195 46.450 102.740 ;
        RECT 46.625 102.195 49.215 102.965 ;
        RECT 49.845 102.195 50.135 102.920 ;
        RECT 51.890 102.740 52.230 103.570 ;
        RECT 53.710 103.060 54.060 104.310 ;
        RECT 57.410 102.740 57.750 103.570 ;
        RECT 59.230 103.060 59.580 104.310 ;
        RECT 62.930 102.740 63.270 103.570 ;
        RECT 64.750 103.060 65.100 104.310 ;
        RECT 68.450 102.740 68.790 103.570 ;
        RECT 70.270 103.060 70.620 104.310 ;
        RECT 72.385 103.655 74.975 104.745 ;
        RECT 72.385 102.965 73.595 103.485 ;
        RECT 73.765 103.135 74.975 103.655 ;
        RECT 75.605 103.580 75.895 104.745 ;
        RECT 76.065 104.310 81.410 104.745 ;
        RECT 81.585 104.310 86.930 104.745 ;
        RECT 87.105 104.310 92.450 104.745 ;
        RECT 92.625 104.310 97.970 104.745 ;
        RECT 50.305 102.195 55.650 102.740 ;
        RECT 55.825 102.195 61.170 102.740 ;
        RECT 61.345 102.195 66.690 102.740 ;
        RECT 66.865 102.195 72.210 102.740 ;
        RECT 72.385 102.195 74.975 102.965 ;
        RECT 75.605 102.195 75.895 102.920 ;
        RECT 77.650 102.740 77.990 103.570 ;
        RECT 79.470 103.060 79.820 104.310 ;
        RECT 83.170 102.740 83.510 103.570 ;
        RECT 84.990 103.060 85.340 104.310 ;
        RECT 88.690 102.740 89.030 103.570 ;
        RECT 90.510 103.060 90.860 104.310 ;
        RECT 94.210 102.740 94.550 103.570 ;
        RECT 96.030 103.060 96.380 104.310 ;
        RECT 98.145 103.655 100.735 104.745 ;
        RECT 98.145 102.965 99.355 103.485 ;
        RECT 99.525 103.135 100.735 103.655 ;
        RECT 101.365 103.580 101.655 104.745 ;
        RECT 101.825 104.310 107.170 104.745 ;
        RECT 107.345 104.310 112.690 104.745 ;
        RECT 112.865 104.310 118.210 104.745 ;
        RECT 118.385 104.310 123.730 104.745 ;
        RECT 76.065 102.195 81.410 102.740 ;
        RECT 81.585 102.195 86.930 102.740 ;
        RECT 87.105 102.195 92.450 102.740 ;
        RECT 92.625 102.195 97.970 102.740 ;
        RECT 98.145 102.195 100.735 102.965 ;
        RECT 101.365 102.195 101.655 102.920 ;
        RECT 103.410 102.740 103.750 103.570 ;
        RECT 105.230 103.060 105.580 104.310 ;
        RECT 108.930 102.740 109.270 103.570 ;
        RECT 110.750 103.060 111.100 104.310 ;
        RECT 114.450 102.740 114.790 103.570 ;
        RECT 116.270 103.060 116.620 104.310 ;
        RECT 119.970 102.740 120.310 103.570 ;
        RECT 121.790 103.060 122.140 104.310 ;
        RECT 123.905 103.655 126.495 104.745 ;
        RECT 123.905 102.965 125.115 103.485 ;
        RECT 125.285 103.135 126.495 103.655 ;
        RECT 127.125 103.580 127.415 104.745 ;
        RECT 127.585 104.310 132.930 104.745 ;
        RECT 133.105 104.310 138.450 104.745 ;
        RECT 138.625 104.310 143.970 104.745 ;
        RECT 101.825 102.195 107.170 102.740 ;
        RECT 107.345 102.195 112.690 102.740 ;
        RECT 112.865 102.195 118.210 102.740 ;
        RECT 118.385 102.195 123.730 102.740 ;
        RECT 123.905 102.195 126.495 102.965 ;
        RECT 127.125 102.195 127.415 102.920 ;
        RECT 129.170 102.740 129.510 103.570 ;
        RECT 130.990 103.060 131.340 104.310 ;
        RECT 134.690 102.740 135.030 103.570 ;
        RECT 136.510 103.060 136.860 104.310 ;
        RECT 140.210 102.740 140.550 103.570 ;
        RECT 142.030 103.060 142.380 104.310 ;
        RECT 144.145 103.655 147.655 104.745 ;
        RECT 147.825 103.655 149.035 104.745 ;
        RECT 144.145 102.965 145.795 103.485 ;
        RECT 145.965 103.135 147.655 103.655 ;
        RECT 127.585 102.195 132.930 102.740 ;
        RECT 133.105 102.195 138.450 102.740 ;
        RECT 138.625 102.195 143.970 102.740 ;
        RECT 144.145 102.195 147.655 102.965 ;
        RECT 147.825 102.945 148.345 103.485 ;
        RECT 148.515 103.115 149.035 103.655 ;
        RECT 149.205 103.655 150.415 104.745 ;
        RECT 149.205 103.115 149.725 103.655 ;
        RECT 149.895 102.945 150.415 103.485 ;
        RECT 147.825 102.195 149.035 102.945 ;
        RECT 149.205 102.195 150.415 102.945 ;
        RECT 11.120 102.025 150.500 102.195 ;
        RECT 11.205 101.275 12.415 102.025 ;
        RECT 12.585 101.480 17.930 102.025 ;
        RECT 18.105 101.480 23.450 102.025 ;
        RECT 23.625 101.480 28.970 102.025 ;
        RECT 29.145 101.480 34.490 102.025 ;
        RECT 11.205 100.735 11.725 101.275 ;
        RECT 11.895 100.565 12.415 101.105 ;
        RECT 14.170 100.650 14.510 101.480 ;
        RECT 11.205 99.475 12.415 100.565 ;
        RECT 15.990 99.910 16.340 101.160 ;
        RECT 19.690 100.650 20.030 101.480 ;
        RECT 21.510 99.910 21.860 101.160 ;
        RECT 25.210 100.650 25.550 101.480 ;
        RECT 27.030 99.910 27.380 101.160 ;
        RECT 30.730 100.650 31.070 101.480 ;
        RECT 34.665 101.255 36.335 102.025 ;
        RECT 36.965 101.300 37.255 102.025 ;
        RECT 37.425 101.480 42.770 102.025 ;
        RECT 42.945 101.480 48.290 102.025 ;
        RECT 48.465 101.480 53.810 102.025 ;
        RECT 53.985 101.480 59.330 102.025 ;
        RECT 32.550 99.910 32.900 101.160 ;
        RECT 34.665 100.735 35.415 101.255 ;
        RECT 35.585 100.565 36.335 101.085 ;
        RECT 39.010 100.650 39.350 101.480 ;
        RECT 12.585 99.475 17.930 99.910 ;
        RECT 18.105 99.475 23.450 99.910 ;
        RECT 23.625 99.475 28.970 99.910 ;
        RECT 29.145 99.475 34.490 99.910 ;
        RECT 34.665 99.475 36.335 100.565 ;
        RECT 36.965 99.475 37.255 100.640 ;
        RECT 40.830 99.910 41.180 101.160 ;
        RECT 44.530 100.650 44.870 101.480 ;
        RECT 46.350 99.910 46.700 101.160 ;
        RECT 50.050 100.650 50.390 101.480 ;
        RECT 51.870 99.910 52.220 101.160 ;
        RECT 55.570 100.650 55.910 101.480 ;
        RECT 59.505 101.255 62.095 102.025 ;
        RECT 62.725 101.300 63.015 102.025 ;
        RECT 63.185 101.480 68.530 102.025 ;
        RECT 68.705 101.480 74.050 102.025 ;
        RECT 74.225 101.480 79.570 102.025 ;
        RECT 79.745 101.480 85.090 102.025 ;
        RECT 57.390 99.910 57.740 101.160 ;
        RECT 59.505 100.735 60.715 101.255 ;
        RECT 60.885 100.565 62.095 101.085 ;
        RECT 64.770 100.650 65.110 101.480 ;
        RECT 37.425 99.475 42.770 99.910 ;
        RECT 42.945 99.475 48.290 99.910 ;
        RECT 48.465 99.475 53.810 99.910 ;
        RECT 53.985 99.475 59.330 99.910 ;
        RECT 59.505 99.475 62.095 100.565 ;
        RECT 62.725 99.475 63.015 100.640 ;
        RECT 66.590 99.910 66.940 101.160 ;
        RECT 70.290 100.650 70.630 101.480 ;
        RECT 72.110 99.910 72.460 101.160 ;
        RECT 75.810 100.650 76.150 101.480 ;
        RECT 77.630 99.910 77.980 101.160 ;
        RECT 81.330 100.650 81.670 101.480 ;
        RECT 85.265 101.255 87.855 102.025 ;
        RECT 88.485 101.300 88.775 102.025 ;
        RECT 88.945 101.480 94.290 102.025 ;
        RECT 94.465 101.480 99.810 102.025 ;
        RECT 99.985 101.480 105.330 102.025 ;
        RECT 105.505 101.480 110.850 102.025 ;
        RECT 83.150 99.910 83.500 101.160 ;
        RECT 85.265 100.735 86.475 101.255 ;
        RECT 86.645 100.565 87.855 101.085 ;
        RECT 90.530 100.650 90.870 101.480 ;
        RECT 63.185 99.475 68.530 99.910 ;
        RECT 68.705 99.475 74.050 99.910 ;
        RECT 74.225 99.475 79.570 99.910 ;
        RECT 79.745 99.475 85.090 99.910 ;
        RECT 85.265 99.475 87.855 100.565 ;
        RECT 88.485 99.475 88.775 100.640 ;
        RECT 92.350 99.910 92.700 101.160 ;
        RECT 96.050 100.650 96.390 101.480 ;
        RECT 97.870 99.910 98.220 101.160 ;
        RECT 101.570 100.650 101.910 101.480 ;
        RECT 103.390 99.910 103.740 101.160 ;
        RECT 107.090 100.650 107.430 101.480 ;
        RECT 111.025 101.255 113.615 102.025 ;
        RECT 114.245 101.300 114.535 102.025 ;
        RECT 114.705 101.480 120.050 102.025 ;
        RECT 120.225 101.480 125.570 102.025 ;
        RECT 125.745 101.480 131.090 102.025 ;
        RECT 131.265 101.480 136.610 102.025 ;
        RECT 108.910 99.910 109.260 101.160 ;
        RECT 111.025 100.735 112.235 101.255 ;
        RECT 112.405 100.565 113.615 101.085 ;
        RECT 116.290 100.650 116.630 101.480 ;
        RECT 88.945 99.475 94.290 99.910 ;
        RECT 94.465 99.475 99.810 99.910 ;
        RECT 99.985 99.475 105.330 99.910 ;
        RECT 105.505 99.475 110.850 99.910 ;
        RECT 111.025 99.475 113.615 100.565 ;
        RECT 114.245 99.475 114.535 100.640 ;
        RECT 118.110 99.910 118.460 101.160 ;
        RECT 121.810 100.650 122.150 101.480 ;
        RECT 123.630 99.910 123.980 101.160 ;
        RECT 127.330 100.650 127.670 101.480 ;
        RECT 129.150 99.910 129.500 101.160 ;
        RECT 132.850 100.650 133.190 101.480 ;
        RECT 136.785 101.255 139.375 102.025 ;
        RECT 140.005 101.300 140.295 102.025 ;
        RECT 140.465 101.480 145.810 102.025 ;
        RECT 134.670 99.910 135.020 101.160 ;
        RECT 136.785 100.735 137.995 101.255 ;
        RECT 138.165 100.565 139.375 101.085 ;
        RECT 142.050 100.650 142.390 101.480 ;
        RECT 145.985 101.255 148.575 102.025 ;
        RECT 149.205 101.275 150.415 102.025 ;
        RECT 114.705 99.475 120.050 99.910 ;
        RECT 120.225 99.475 125.570 99.910 ;
        RECT 125.745 99.475 131.090 99.910 ;
        RECT 131.265 99.475 136.610 99.910 ;
        RECT 136.785 99.475 139.375 100.565 ;
        RECT 140.005 99.475 140.295 100.640 ;
        RECT 143.870 99.910 144.220 101.160 ;
        RECT 145.985 100.735 147.195 101.255 ;
        RECT 147.365 100.565 148.575 101.085 ;
        RECT 140.465 99.475 145.810 99.910 ;
        RECT 145.985 99.475 148.575 100.565 ;
        RECT 149.205 100.565 149.725 101.105 ;
        RECT 149.895 100.735 150.415 101.275 ;
        RECT 149.205 99.475 150.415 100.565 ;
        RECT 11.120 99.305 150.500 99.475 ;
        RECT 11.205 98.215 12.415 99.305 ;
        RECT 12.585 98.870 17.930 99.305 ;
        RECT 18.105 98.870 23.450 99.305 ;
        RECT 11.205 97.505 11.725 98.045 ;
        RECT 11.895 97.675 12.415 98.215 ;
        RECT 11.205 96.755 12.415 97.505 ;
        RECT 14.170 97.300 14.510 98.130 ;
        RECT 15.990 97.620 16.340 98.870 ;
        RECT 19.690 97.300 20.030 98.130 ;
        RECT 21.510 97.620 21.860 98.870 ;
        RECT 24.085 98.140 24.375 99.305 ;
        RECT 24.545 98.870 29.890 99.305 ;
        RECT 30.065 98.870 35.410 99.305 ;
        RECT 35.585 98.870 40.930 99.305 ;
        RECT 41.105 98.870 46.450 99.305 ;
        RECT 12.585 96.755 17.930 97.300 ;
        RECT 18.105 96.755 23.450 97.300 ;
        RECT 24.085 96.755 24.375 97.480 ;
        RECT 26.130 97.300 26.470 98.130 ;
        RECT 27.950 97.620 28.300 98.870 ;
        RECT 31.650 97.300 31.990 98.130 ;
        RECT 33.470 97.620 33.820 98.870 ;
        RECT 37.170 97.300 37.510 98.130 ;
        RECT 38.990 97.620 39.340 98.870 ;
        RECT 42.690 97.300 43.030 98.130 ;
        RECT 44.510 97.620 44.860 98.870 ;
        RECT 46.625 98.215 49.215 99.305 ;
        RECT 46.625 97.525 47.835 98.045 ;
        RECT 48.005 97.695 49.215 98.215 ;
        RECT 49.845 98.140 50.135 99.305 ;
        RECT 50.305 98.870 55.650 99.305 ;
        RECT 55.825 98.870 61.170 99.305 ;
        RECT 61.345 98.870 66.690 99.305 ;
        RECT 66.865 98.870 72.210 99.305 ;
        RECT 24.545 96.755 29.890 97.300 ;
        RECT 30.065 96.755 35.410 97.300 ;
        RECT 35.585 96.755 40.930 97.300 ;
        RECT 41.105 96.755 46.450 97.300 ;
        RECT 46.625 96.755 49.215 97.525 ;
        RECT 49.845 96.755 50.135 97.480 ;
        RECT 51.890 97.300 52.230 98.130 ;
        RECT 53.710 97.620 54.060 98.870 ;
        RECT 57.410 97.300 57.750 98.130 ;
        RECT 59.230 97.620 59.580 98.870 ;
        RECT 62.930 97.300 63.270 98.130 ;
        RECT 64.750 97.620 65.100 98.870 ;
        RECT 68.450 97.300 68.790 98.130 ;
        RECT 70.270 97.620 70.620 98.870 ;
        RECT 72.385 98.215 74.975 99.305 ;
        RECT 72.385 97.525 73.595 98.045 ;
        RECT 73.765 97.695 74.975 98.215 ;
        RECT 75.605 98.140 75.895 99.305 ;
        RECT 76.065 98.870 81.410 99.305 ;
        RECT 81.585 98.870 86.930 99.305 ;
        RECT 87.105 98.870 92.450 99.305 ;
        RECT 92.625 98.870 97.970 99.305 ;
        RECT 50.305 96.755 55.650 97.300 ;
        RECT 55.825 96.755 61.170 97.300 ;
        RECT 61.345 96.755 66.690 97.300 ;
        RECT 66.865 96.755 72.210 97.300 ;
        RECT 72.385 96.755 74.975 97.525 ;
        RECT 75.605 96.755 75.895 97.480 ;
        RECT 77.650 97.300 77.990 98.130 ;
        RECT 79.470 97.620 79.820 98.870 ;
        RECT 83.170 97.300 83.510 98.130 ;
        RECT 84.990 97.620 85.340 98.870 ;
        RECT 88.690 97.300 89.030 98.130 ;
        RECT 90.510 97.620 90.860 98.870 ;
        RECT 94.210 97.300 94.550 98.130 ;
        RECT 96.030 97.620 96.380 98.870 ;
        RECT 98.145 98.215 100.735 99.305 ;
        RECT 98.145 97.525 99.355 98.045 ;
        RECT 99.525 97.695 100.735 98.215 ;
        RECT 101.365 98.140 101.655 99.305 ;
        RECT 101.825 98.870 107.170 99.305 ;
        RECT 107.345 98.870 112.690 99.305 ;
        RECT 112.865 98.870 118.210 99.305 ;
        RECT 118.385 98.870 123.730 99.305 ;
        RECT 76.065 96.755 81.410 97.300 ;
        RECT 81.585 96.755 86.930 97.300 ;
        RECT 87.105 96.755 92.450 97.300 ;
        RECT 92.625 96.755 97.970 97.300 ;
        RECT 98.145 96.755 100.735 97.525 ;
        RECT 101.365 96.755 101.655 97.480 ;
        RECT 103.410 97.300 103.750 98.130 ;
        RECT 105.230 97.620 105.580 98.870 ;
        RECT 108.930 97.300 109.270 98.130 ;
        RECT 110.750 97.620 111.100 98.870 ;
        RECT 114.450 97.300 114.790 98.130 ;
        RECT 116.270 97.620 116.620 98.870 ;
        RECT 119.970 97.300 120.310 98.130 ;
        RECT 121.790 97.620 122.140 98.870 ;
        RECT 123.905 98.215 126.495 99.305 ;
        RECT 123.905 97.525 125.115 98.045 ;
        RECT 125.285 97.695 126.495 98.215 ;
        RECT 127.125 98.140 127.415 99.305 ;
        RECT 127.585 98.870 132.930 99.305 ;
        RECT 133.105 98.870 138.450 99.305 ;
        RECT 138.625 98.870 143.970 99.305 ;
        RECT 101.825 96.755 107.170 97.300 ;
        RECT 107.345 96.755 112.690 97.300 ;
        RECT 112.865 96.755 118.210 97.300 ;
        RECT 118.385 96.755 123.730 97.300 ;
        RECT 123.905 96.755 126.495 97.525 ;
        RECT 127.125 96.755 127.415 97.480 ;
        RECT 129.170 97.300 129.510 98.130 ;
        RECT 130.990 97.620 131.340 98.870 ;
        RECT 134.690 97.300 135.030 98.130 ;
        RECT 136.510 97.620 136.860 98.870 ;
        RECT 140.210 97.300 140.550 98.130 ;
        RECT 142.030 97.620 142.380 98.870 ;
        RECT 144.145 98.215 147.655 99.305 ;
        RECT 147.825 98.215 149.035 99.305 ;
        RECT 144.145 97.525 145.795 98.045 ;
        RECT 145.965 97.695 147.655 98.215 ;
        RECT 127.585 96.755 132.930 97.300 ;
        RECT 133.105 96.755 138.450 97.300 ;
        RECT 138.625 96.755 143.970 97.300 ;
        RECT 144.145 96.755 147.655 97.525 ;
        RECT 147.825 97.505 148.345 98.045 ;
        RECT 148.515 97.675 149.035 98.215 ;
        RECT 149.205 98.215 150.415 99.305 ;
        RECT 149.205 97.675 149.725 98.215 ;
        RECT 149.895 97.505 150.415 98.045 ;
        RECT 147.825 96.755 149.035 97.505 ;
        RECT 149.205 96.755 150.415 97.505 ;
        RECT 11.120 96.585 150.500 96.755 ;
        RECT 11.205 95.835 12.415 96.585 ;
        RECT 12.585 96.040 17.930 96.585 ;
        RECT 18.105 96.040 23.450 96.585 ;
        RECT 23.625 96.040 28.970 96.585 ;
        RECT 29.145 96.040 34.490 96.585 ;
        RECT 11.205 95.295 11.725 95.835 ;
        RECT 11.895 95.125 12.415 95.665 ;
        RECT 14.170 95.210 14.510 96.040 ;
        RECT 11.205 94.035 12.415 95.125 ;
        RECT 15.990 94.470 16.340 95.720 ;
        RECT 19.690 95.210 20.030 96.040 ;
        RECT 21.510 94.470 21.860 95.720 ;
        RECT 25.210 95.210 25.550 96.040 ;
        RECT 27.030 94.470 27.380 95.720 ;
        RECT 30.730 95.210 31.070 96.040 ;
        RECT 34.665 95.815 36.335 96.585 ;
        RECT 36.965 95.860 37.255 96.585 ;
        RECT 37.425 96.040 42.770 96.585 ;
        RECT 42.945 96.040 48.290 96.585 ;
        RECT 48.465 96.040 53.810 96.585 ;
        RECT 53.985 96.040 59.330 96.585 ;
        RECT 32.550 94.470 32.900 95.720 ;
        RECT 34.665 95.295 35.415 95.815 ;
        RECT 35.585 95.125 36.335 95.645 ;
        RECT 39.010 95.210 39.350 96.040 ;
        RECT 12.585 94.035 17.930 94.470 ;
        RECT 18.105 94.035 23.450 94.470 ;
        RECT 23.625 94.035 28.970 94.470 ;
        RECT 29.145 94.035 34.490 94.470 ;
        RECT 34.665 94.035 36.335 95.125 ;
        RECT 36.965 94.035 37.255 95.200 ;
        RECT 40.830 94.470 41.180 95.720 ;
        RECT 44.530 95.210 44.870 96.040 ;
        RECT 46.350 94.470 46.700 95.720 ;
        RECT 50.050 95.210 50.390 96.040 ;
        RECT 51.870 94.470 52.220 95.720 ;
        RECT 55.570 95.210 55.910 96.040 ;
        RECT 59.505 95.815 62.095 96.585 ;
        RECT 62.725 95.860 63.015 96.585 ;
        RECT 63.185 96.040 68.530 96.585 ;
        RECT 68.705 96.040 74.050 96.585 ;
        RECT 74.225 96.040 79.570 96.585 ;
        RECT 79.745 96.040 85.090 96.585 ;
        RECT 57.390 94.470 57.740 95.720 ;
        RECT 59.505 95.295 60.715 95.815 ;
        RECT 60.885 95.125 62.095 95.645 ;
        RECT 64.770 95.210 65.110 96.040 ;
        RECT 37.425 94.035 42.770 94.470 ;
        RECT 42.945 94.035 48.290 94.470 ;
        RECT 48.465 94.035 53.810 94.470 ;
        RECT 53.985 94.035 59.330 94.470 ;
        RECT 59.505 94.035 62.095 95.125 ;
        RECT 62.725 94.035 63.015 95.200 ;
        RECT 66.590 94.470 66.940 95.720 ;
        RECT 70.290 95.210 70.630 96.040 ;
        RECT 72.110 94.470 72.460 95.720 ;
        RECT 75.810 95.210 76.150 96.040 ;
        RECT 77.630 94.470 77.980 95.720 ;
        RECT 81.330 95.210 81.670 96.040 ;
        RECT 85.265 95.815 87.855 96.585 ;
        RECT 88.485 95.860 88.775 96.585 ;
        RECT 88.945 96.040 94.290 96.585 ;
        RECT 94.465 96.040 99.810 96.585 ;
        RECT 99.985 96.040 105.330 96.585 ;
        RECT 105.505 96.040 110.850 96.585 ;
        RECT 83.150 94.470 83.500 95.720 ;
        RECT 85.265 95.295 86.475 95.815 ;
        RECT 86.645 95.125 87.855 95.645 ;
        RECT 90.530 95.210 90.870 96.040 ;
        RECT 63.185 94.035 68.530 94.470 ;
        RECT 68.705 94.035 74.050 94.470 ;
        RECT 74.225 94.035 79.570 94.470 ;
        RECT 79.745 94.035 85.090 94.470 ;
        RECT 85.265 94.035 87.855 95.125 ;
        RECT 88.485 94.035 88.775 95.200 ;
        RECT 92.350 94.470 92.700 95.720 ;
        RECT 96.050 95.210 96.390 96.040 ;
        RECT 97.870 94.470 98.220 95.720 ;
        RECT 101.570 95.210 101.910 96.040 ;
        RECT 103.390 94.470 103.740 95.720 ;
        RECT 107.090 95.210 107.430 96.040 ;
        RECT 111.025 95.815 113.615 96.585 ;
        RECT 114.245 95.860 114.535 96.585 ;
        RECT 114.705 96.040 120.050 96.585 ;
        RECT 120.225 96.040 125.570 96.585 ;
        RECT 125.745 96.040 131.090 96.585 ;
        RECT 131.265 96.040 136.610 96.585 ;
        RECT 108.910 94.470 109.260 95.720 ;
        RECT 111.025 95.295 112.235 95.815 ;
        RECT 112.405 95.125 113.615 95.645 ;
        RECT 116.290 95.210 116.630 96.040 ;
        RECT 88.945 94.035 94.290 94.470 ;
        RECT 94.465 94.035 99.810 94.470 ;
        RECT 99.985 94.035 105.330 94.470 ;
        RECT 105.505 94.035 110.850 94.470 ;
        RECT 111.025 94.035 113.615 95.125 ;
        RECT 114.245 94.035 114.535 95.200 ;
        RECT 118.110 94.470 118.460 95.720 ;
        RECT 121.810 95.210 122.150 96.040 ;
        RECT 123.630 94.470 123.980 95.720 ;
        RECT 127.330 95.210 127.670 96.040 ;
        RECT 129.150 94.470 129.500 95.720 ;
        RECT 132.850 95.210 133.190 96.040 ;
        RECT 136.785 95.815 139.375 96.585 ;
        RECT 140.005 95.860 140.295 96.585 ;
        RECT 140.465 96.040 145.810 96.585 ;
        RECT 134.670 94.470 135.020 95.720 ;
        RECT 136.785 95.295 137.995 95.815 ;
        RECT 138.165 95.125 139.375 95.645 ;
        RECT 142.050 95.210 142.390 96.040 ;
        RECT 145.985 95.815 148.575 96.585 ;
        RECT 149.205 95.835 150.415 96.585 ;
        RECT 114.705 94.035 120.050 94.470 ;
        RECT 120.225 94.035 125.570 94.470 ;
        RECT 125.745 94.035 131.090 94.470 ;
        RECT 131.265 94.035 136.610 94.470 ;
        RECT 136.785 94.035 139.375 95.125 ;
        RECT 140.005 94.035 140.295 95.200 ;
        RECT 143.870 94.470 144.220 95.720 ;
        RECT 145.985 95.295 147.195 95.815 ;
        RECT 147.365 95.125 148.575 95.645 ;
        RECT 140.465 94.035 145.810 94.470 ;
        RECT 145.985 94.035 148.575 95.125 ;
        RECT 149.205 95.125 149.725 95.665 ;
        RECT 149.895 95.295 150.415 95.835 ;
        RECT 149.205 94.035 150.415 95.125 ;
        RECT 11.120 93.865 150.500 94.035 ;
        RECT 11.205 92.775 12.415 93.865 ;
        RECT 12.585 93.430 17.930 93.865 ;
        RECT 18.105 93.430 23.450 93.865 ;
        RECT 11.205 92.065 11.725 92.605 ;
        RECT 11.895 92.235 12.415 92.775 ;
        RECT 11.205 91.315 12.415 92.065 ;
        RECT 14.170 91.860 14.510 92.690 ;
        RECT 15.990 92.180 16.340 93.430 ;
        RECT 19.690 91.860 20.030 92.690 ;
        RECT 21.510 92.180 21.860 93.430 ;
        RECT 24.085 92.700 24.375 93.865 ;
        RECT 24.545 93.430 29.890 93.865 ;
        RECT 30.065 93.430 35.410 93.865 ;
        RECT 35.585 93.430 40.930 93.865 ;
        RECT 41.105 93.430 46.450 93.865 ;
        RECT 12.585 91.315 17.930 91.860 ;
        RECT 18.105 91.315 23.450 91.860 ;
        RECT 24.085 91.315 24.375 92.040 ;
        RECT 26.130 91.860 26.470 92.690 ;
        RECT 27.950 92.180 28.300 93.430 ;
        RECT 31.650 91.860 31.990 92.690 ;
        RECT 33.470 92.180 33.820 93.430 ;
        RECT 37.170 91.860 37.510 92.690 ;
        RECT 38.990 92.180 39.340 93.430 ;
        RECT 42.690 91.860 43.030 92.690 ;
        RECT 44.510 92.180 44.860 93.430 ;
        RECT 46.625 92.775 49.215 93.865 ;
        RECT 46.625 92.085 47.835 92.605 ;
        RECT 48.005 92.255 49.215 92.775 ;
        RECT 49.845 92.700 50.135 93.865 ;
        RECT 50.305 93.430 55.650 93.865 ;
        RECT 55.825 93.430 61.170 93.865 ;
        RECT 61.345 93.430 66.690 93.865 ;
        RECT 66.865 93.430 72.210 93.865 ;
        RECT 24.545 91.315 29.890 91.860 ;
        RECT 30.065 91.315 35.410 91.860 ;
        RECT 35.585 91.315 40.930 91.860 ;
        RECT 41.105 91.315 46.450 91.860 ;
        RECT 46.625 91.315 49.215 92.085 ;
        RECT 49.845 91.315 50.135 92.040 ;
        RECT 51.890 91.860 52.230 92.690 ;
        RECT 53.710 92.180 54.060 93.430 ;
        RECT 57.410 91.860 57.750 92.690 ;
        RECT 59.230 92.180 59.580 93.430 ;
        RECT 62.930 91.860 63.270 92.690 ;
        RECT 64.750 92.180 65.100 93.430 ;
        RECT 68.450 91.860 68.790 92.690 ;
        RECT 70.270 92.180 70.620 93.430 ;
        RECT 72.385 92.775 74.975 93.865 ;
        RECT 72.385 92.085 73.595 92.605 ;
        RECT 73.765 92.255 74.975 92.775 ;
        RECT 75.605 92.700 75.895 93.865 ;
        RECT 76.065 93.430 81.410 93.865 ;
        RECT 81.585 93.430 86.930 93.865 ;
        RECT 87.105 93.430 92.450 93.865 ;
        RECT 92.625 93.430 97.970 93.865 ;
        RECT 50.305 91.315 55.650 91.860 ;
        RECT 55.825 91.315 61.170 91.860 ;
        RECT 61.345 91.315 66.690 91.860 ;
        RECT 66.865 91.315 72.210 91.860 ;
        RECT 72.385 91.315 74.975 92.085 ;
        RECT 75.605 91.315 75.895 92.040 ;
        RECT 77.650 91.860 77.990 92.690 ;
        RECT 79.470 92.180 79.820 93.430 ;
        RECT 83.170 91.860 83.510 92.690 ;
        RECT 84.990 92.180 85.340 93.430 ;
        RECT 88.690 91.860 89.030 92.690 ;
        RECT 90.510 92.180 90.860 93.430 ;
        RECT 94.210 91.860 94.550 92.690 ;
        RECT 96.030 92.180 96.380 93.430 ;
        RECT 98.145 92.775 100.735 93.865 ;
        RECT 98.145 92.085 99.355 92.605 ;
        RECT 99.525 92.255 100.735 92.775 ;
        RECT 101.365 92.700 101.655 93.865 ;
        RECT 101.825 93.430 107.170 93.865 ;
        RECT 107.345 93.430 112.690 93.865 ;
        RECT 112.865 93.430 118.210 93.865 ;
        RECT 118.385 93.430 123.730 93.865 ;
        RECT 76.065 91.315 81.410 91.860 ;
        RECT 81.585 91.315 86.930 91.860 ;
        RECT 87.105 91.315 92.450 91.860 ;
        RECT 92.625 91.315 97.970 91.860 ;
        RECT 98.145 91.315 100.735 92.085 ;
        RECT 101.365 91.315 101.655 92.040 ;
        RECT 103.410 91.860 103.750 92.690 ;
        RECT 105.230 92.180 105.580 93.430 ;
        RECT 108.930 91.860 109.270 92.690 ;
        RECT 110.750 92.180 111.100 93.430 ;
        RECT 114.450 91.860 114.790 92.690 ;
        RECT 116.270 92.180 116.620 93.430 ;
        RECT 119.970 91.860 120.310 92.690 ;
        RECT 121.790 92.180 122.140 93.430 ;
        RECT 123.905 92.775 126.495 93.865 ;
        RECT 123.905 92.085 125.115 92.605 ;
        RECT 125.285 92.255 126.495 92.775 ;
        RECT 127.125 92.700 127.415 93.865 ;
        RECT 127.585 93.430 132.930 93.865 ;
        RECT 133.105 93.430 138.450 93.865 ;
        RECT 138.625 93.430 143.970 93.865 ;
        RECT 101.825 91.315 107.170 91.860 ;
        RECT 107.345 91.315 112.690 91.860 ;
        RECT 112.865 91.315 118.210 91.860 ;
        RECT 118.385 91.315 123.730 91.860 ;
        RECT 123.905 91.315 126.495 92.085 ;
        RECT 127.125 91.315 127.415 92.040 ;
        RECT 129.170 91.860 129.510 92.690 ;
        RECT 130.990 92.180 131.340 93.430 ;
        RECT 134.690 91.860 135.030 92.690 ;
        RECT 136.510 92.180 136.860 93.430 ;
        RECT 140.210 91.860 140.550 92.690 ;
        RECT 142.030 92.180 142.380 93.430 ;
        RECT 144.145 92.775 147.655 93.865 ;
        RECT 147.825 92.775 149.035 93.865 ;
        RECT 144.145 92.085 145.795 92.605 ;
        RECT 145.965 92.255 147.655 92.775 ;
        RECT 127.585 91.315 132.930 91.860 ;
        RECT 133.105 91.315 138.450 91.860 ;
        RECT 138.625 91.315 143.970 91.860 ;
        RECT 144.145 91.315 147.655 92.085 ;
        RECT 147.825 92.065 148.345 92.605 ;
        RECT 148.515 92.235 149.035 92.775 ;
        RECT 149.205 92.775 150.415 93.865 ;
        RECT 149.205 92.235 149.725 92.775 ;
        RECT 149.895 92.065 150.415 92.605 ;
        RECT 147.825 91.315 149.035 92.065 ;
        RECT 149.205 91.315 150.415 92.065 ;
        RECT 11.120 91.145 150.500 91.315 ;
        RECT 11.205 90.395 12.415 91.145 ;
        RECT 12.585 90.600 17.930 91.145 ;
        RECT 18.105 90.600 23.450 91.145 ;
        RECT 23.625 90.600 28.970 91.145 ;
        RECT 29.145 90.600 34.490 91.145 ;
        RECT 11.205 89.855 11.725 90.395 ;
        RECT 11.895 89.685 12.415 90.225 ;
        RECT 14.170 89.770 14.510 90.600 ;
        RECT 11.205 88.595 12.415 89.685 ;
        RECT 15.990 89.030 16.340 90.280 ;
        RECT 19.690 89.770 20.030 90.600 ;
        RECT 21.510 89.030 21.860 90.280 ;
        RECT 25.210 89.770 25.550 90.600 ;
        RECT 27.030 89.030 27.380 90.280 ;
        RECT 30.730 89.770 31.070 90.600 ;
        RECT 34.665 90.375 36.335 91.145 ;
        RECT 36.965 90.420 37.255 91.145 ;
        RECT 37.425 90.600 42.770 91.145 ;
        RECT 42.945 90.600 48.290 91.145 ;
        RECT 48.465 90.600 53.810 91.145 ;
        RECT 53.985 90.600 59.330 91.145 ;
        RECT 32.550 89.030 32.900 90.280 ;
        RECT 34.665 89.855 35.415 90.375 ;
        RECT 35.585 89.685 36.335 90.205 ;
        RECT 39.010 89.770 39.350 90.600 ;
        RECT 12.585 88.595 17.930 89.030 ;
        RECT 18.105 88.595 23.450 89.030 ;
        RECT 23.625 88.595 28.970 89.030 ;
        RECT 29.145 88.595 34.490 89.030 ;
        RECT 34.665 88.595 36.335 89.685 ;
        RECT 36.965 88.595 37.255 89.760 ;
        RECT 40.830 89.030 41.180 90.280 ;
        RECT 44.530 89.770 44.870 90.600 ;
        RECT 46.350 89.030 46.700 90.280 ;
        RECT 50.050 89.770 50.390 90.600 ;
        RECT 51.870 89.030 52.220 90.280 ;
        RECT 55.570 89.770 55.910 90.600 ;
        RECT 59.505 90.375 62.095 91.145 ;
        RECT 62.725 90.420 63.015 91.145 ;
        RECT 63.185 90.600 68.530 91.145 ;
        RECT 68.705 90.600 74.050 91.145 ;
        RECT 74.225 90.600 79.570 91.145 ;
        RECT 79.745 90.600 85.090 91.145 ;
        RECT 57.390 89.030 57.740 90.280 ;
        RECT 59.505 89.855 60.715 90.375 ;
        RECT 60.885 89.685 62.095 90.205 ;
        RECT 64.770 89.770 65.110 90.600 ;
        RECT 37.425 88.595 42.770 89.030 ;
        RECT 42.945 88.595 48.290 89.030 ;
        RECT 48.465 88.595 53.810 89.030 ;
        RECT 53.985 88.595 59.330 89.030 ;
        RECT 59.505 88.595 62.095 89.685 ;
        RECT 62.725 88.595 63.015 89.760 ;
        RECT 66.590 89.030 66.940 90.280 ;
        RECT 70.290 89.770 70.630 90.600 ;
        RECT 72.110 89.030 72.460 90.280 ;
        RECT 75.810 89.770 76.150 90.600 ;
        RECT 77.630 89.030 77.980 90.280 ;
        RECT 81.330 89.770 81.670 90.600 ;
        RECT 85.265 90.375 87.855 91.145 ;
        RECT 88.485 90.420 88.775 91.145 ;
        RECT 88.945 90.600 94.290 91.145 ;
        RECT 94.465 90.600 99.810 91.145 ;
        RECT 99.985 90.600 105.330 91.145 ;
        RECT 105.505 90.600 110.850 91.145 ;
        RECT 83.150 89.030 83.500 90.280 ;
        RECT 85.265 89.855 86.475 90.375 ;
        RECT 86.645 89.685 87.855 90.205 ;
        RECT 90.530 89.770 90.870 90.600 ;
        RECT 63.185 88.595 68.530 89.030 ;
        RECT 68.705 88.595 74.050 89.030 ;
        RECT 74.225 88.595 79.570 89.030 ;
        RECT 79.745 88.595 85.090 89.030 ;
        RECT 85.265 88.595 87.855 89.685 ;
        RECT 88.485 88.595 88.775 89.760 ;
        RECT 92.350 89.030 92.700 90.280 ;
        RECT 96.050 89.770 96.390 90.600 ;
        RECT 97.870 89.030 98.220 90.280 ;
        RECT 101.570 89.770 101.910 90.600 ;
        RECT 103.390 89.030 103.740 90.280 ;
        RECT 107.090 89.770 107.430 90.600 ;
        RECT 111.025 90.375 113.615 91.145 ;
        RECT 114.245 90.420 114.535 91.145 ;
        RECT 114.705 90.600 120.050 91.145 ;
        RECT 120.225 90.600 125.570 91.145 ;
        RECT 125.745 90.600 131.090 91.145 ;
        RECT 131.265 90.600 136.610 91.145 ;
        RECT 108.910 89.030 109.260 90.280 ;
        RECT 111.025 89.855 112.235 90.375 ;
        RECT 112.405 89.685 113.615 90.205 ;
        RECT 116.290 89.770 116.630 90.600 ;
        RECT 88.945 88.595 94.290 89.030 ;
        RECT 94.465 88.595 99.810 89.030 ;
        RECT 99.985 88.595 105.330 89.030 ;
        RECT 105.505 88.595 110.850 89.030 ;
        RECT 111.025 88.595 113.615 89.685 ;
        RECT 114.245 88.595 114.535 89.760 ;
        RECT 118.110 89.030 118.460 90.280 ;
        RECT 121.810 89.770 122.150 90.600 ;
        RECT 123.630 89.030 123.980 90.280 ;
        RECT 127.330 89.770 127.670 90.600 ;
        RECT 129.150 89.030 129.500 90.280 ;
        RECT 132.850 89.770 133.190 90.600 ;
        RECT 136.785 90.375 139.375 91.145 ;
        RECT 140.005 90.420 140.295 91.145 ;
        RECT 140.465 90.600 145.810 91.145 ;
        RECT 134.670 89.030 135.020 90.280 ;
        RECT 136.785 89.855 137.995 90.375 ;
        RECT 138.165 89.685 139.375 90.205 ;
        RECT 142.050 89.770 142.390 90.600 ;
        RECT 145.985 90.375 148.575 91.145 ;
        RECT 149.205 90.395 150.415 91.145 ;
        RECT 114.705 88.595 120.050 89.030 ;
        RECT 120.225 88.595 125.570 89.030 ;
        RECT 125.745 88.595 131.090 89.030 ;
        RECT 131.265 88.595 136.610 89.030 ;
        RECT 136.785 88.595 139.375 89.685 ;
        RECT 140.005 88.595 140.295 89.760 ;
        RECT 143.870 89.030 144.220 90.280 ;
        RECT 145.985 89.855 147.195 90.375 ;
        RECT 147.365 89.685 148.575 90.205 ;
        RECT 140.465 88.595 145.810 89.030 ;
        RECT 145.985 88.595 148.575 89.685 ;
        RECT 149.205 89.685 149.725 90.225 ;
        RECT 149.895 89.855 150.415 90.395 ;
        RECT 149.205 88.595 150.415 89.685 ;
        RECT 11.120 88.425 150.500 88.595 ;
        RECT 11.205 87.335 12.415 88.425 ;
        RECT 12.585 87.990 17.930 88.425 ;
        RECT 18.105 87.990 23.450 88.425 ;
        RECT 11.205 86.625 11.725 87.165 ;
        RECT 11.895 86.795 12.415 87.335 ;
        RECT 11.205 85.875 12.415 86.625 ;
        RECT 14.170 86.420 14.510 87.250 ;
        RECT 15.990 86.740 16.340 87.990 ;
        RECT 19.690 86.420 20.030 87.250 ;
        RECT 21.510 86.740 21.860 87.990 ;
        RECT 24.085 87.260 24.375 88.425 ;
        RECT 24.545 87.990 29.890 88.425 ;
        RECT 30.065 87.990 35.410 88.425 ;
        RECT 35.585 87.990 40.930 88.425 ;
        RECT 41.105 87.990 46.450 88.425 ;
        RECT 12.585 85.875 17.930 86.420 ;
        RECT 18.105 85.875 23.450 86.420 ;
        RECT 24.085 85.875 24.375 86.600 ;
        RECT 26.130 86.420 26.470 87.250 ;
        RECT 27.950 86.740 28.300 87.990 ;
        RECT 31.650 86.420 31.990 87.250 ;
        RECT 33.470 86.740 33.820 87.990 ;
        RECT 37.170 86.420 37.510 87.250 ;
        RECT 38.990 86.740 39.340 87.990 ;
        RECT 42.690 86.420 43.030 87.250 ;
        RECT 44.510 86.740 44.860 87.990 ;
        RECT 46.625 87.335 49.215 88.425 ;
        RECT 46.625 86.645 47.835 87.165 ;
        RECT 48.005 86.815 49.215 87.335 ;
        RECT 49.845 87.260 50.135 88.425 ;
        RECT 50.305 87.990 55.650 88.425 ;
        RECT 55.825 87.990 61.170 88.425 ;
        RECT 61.345 87.990 66.690 88.425 ;
        RECT 66.865 87.990 72.210 88.425 ;
        RECT 24.545 85.875 29.890 86.420 ;
        RECT 30.065 85.875 35.410 86.420 ;
        RECT 35.585 85.875 40.930 86.420 ;
        RECT 41.105 85.875 46.450 86.420 ;
        RECT 46.625 85.875 49.215 86.645 ;
        RECT 49.845 85.875 50.135 86.600 ;
        RECT 51.890 86.420 52.230 87.250 ;
        RECT 53.710 86.740 54.060 87.990 ;
        RECT 57.410 86.420 57.750 87.250 ;
        RECT 59.230 86.740 59.580 87.990 ;
        RECT 62.930 86.420 63.270 87.250 ;
        RECT 64.750 86.740 65.100 87.990 ;
        RECT 68.450 86.420 68.790 87.250 ;
        RECT 70.270 86.740 70.620 87.990 ;
        RECT 72.385 87.335 74.975 88.425 ;
        RECT 72.385 86.645 73.595 87.165 ;
        RECT 73.765 86.815 74.975 87.335 ;
        RECT 75.605 87.260 75.895 88.425 ;
        RECT 76.065 87.990 81.410 88.425 ;
        RECT 81.585 87.990 86.930 88.425 ;
        RECT 87.105 87.990 92.450 88.425 ;
        RECT 92.625 87.990 97.970 88.425 ;
        RECT 50.305 85.875 55.650 86.420 ;
        RECT 55.825 85.875 61.170 86.420 ;
        RECT 61.345 85.875 66.690 86.420 ;
        RECT 66.865 85.875 72.210 86.420 ;
        RECT 72.385 85.875 74.975 86.645 ;
        RECT 75.605 85.875 75.895 86.600 ;
        RECT 77.650 86.420 77.990 87.250 ;
        RECT 79.470 86.740 79.820 87.990 ;
        RECT 83.170 86.420 83.510 87.250 ;
        RECT 84.990 86.740 85.340 87.990 ;
        RECT 88.690 86.420 89.030 87.250 ;
        RECT 90.510 86.740 90.860 87.990 ;
        RECT 94.210 86.420 94.550 87.250 ;
        RECT 96.030 86.740 96.380 87.990 ;
        RECT 98.145 87.335 100.735 88.425 ;
        RECT 98.145 86.645 99.355 87.165 ;
        RECT 99.525 86.815 100.735 87.335 ;
        RECT 101.365 87.260 101.655 88.425 ;
        RECT 101.825 87.990 107.170 88.425 ;
        RECT 107.345 87.990 112.690 88.425 ;
        RECT 112.865 87.990 118.210 88.425 ;
        RECT 118.385 87.990 123.730 88.425 ;
        RECT 76.065 85.875 81.410 86.420 ;
        RECT 81.585 85.875 86.930 86.420 ;
        RECT 87.105 85.875 92.450 86.420 ;
        RECT 92.625 85.875 97.970 86.420 ;
        RECT 98.145 85.875 100.735 86.645 ;
        RECT 101.365 85.875 101.655 86.600 ;
        RECT 103.410 86.420 103.750 87.250 ;
        RECT 105.230 86.740 105.580 87.990 ;
        RECT 108.930 86.420 109.270 87.250 ;
        RECT 110.750 86.740 111.100 87.990 ;
        RECT 114.450 86.420 114.790 87.250 ;
        RECT 116.270 86.740 116.620 87.990 ;
        RECT 119.970 86.420 120.310 87.250 ;
        RECT 121.790 86.740 122.140 87.990 ;
        RECT 123.905 87.335 126.495 88.425 ;
        RECT 123.905 86.645 125.115 87.165 ;
        RECT 125.285 86.815 126.495 87.335 ;
        RECT 127.125 87.260 127.415 88.425 ;
        RECT 127.585 87.990 132.930 88.425 ;
        RECT 133.105 87.990 138.450 88.425 ;
        RECT 138.625 87.990 143.970 88.425 ;
        RECT 101.825 85.875 107.170 86.420 ;
        RECT 107.345 85.875 112.690 86.420 ;
        RECT 112.865 85.875 118.210 86.420 ;
        RECT 118.385 85.875 123.730 86.420 ;
        RECT 123.905 85.875 126.495 86.645 ;
        RECT 127.125 85.875 127.415 86.600 ;
        RECT 129.170 86.420 129.510 87.250 ;
        RECT 130.990 86.740 131.340 87.990 ;
        RECT 134.690 86.420 135.030 87.250 ;
        RECT 136.510 86.740 136.860 87.990 ;
        RECT 140.210 86.420 140.550 87.250 ;
        RECT 142.030 86.740 142.380 87.990 ;
        RECT 144.145 87.335 147.655 88.425 ;
        RECT 147.825 87.335 149.035 88.425 ;
        RECT 144.145 86.645 145.795 87.165 ;
        RECT 145.965 86.815 147.655 87.335 ;
        RECT 127.585 85.875 132.930 86.420 ;
        RECT 133.105 85.875 138.450 86.420 ;
        RECT 138.625 85.875 143.970 86.420 ;
        RECT 144.145 85.875 147.655 86.645 ;
        RECT 147.825 86.625 148.345 87.165 ;
        RECT 148.515 86.795 149.035 87.335 ;
        RECT 149.205 87.335 150.415 88.425 ;
        RECT 149.205 86.795 149.725 87.335 ;
        RECT 149.895 86.625 150.415 87.165 ;
        RECT 147.825 85.875 149.035 86.625 ;
        RECT 149.205 85.875 150.415 86.625 ;
        RECT 11.120 85.705 150.500 85.875 ;
        RECT 11.205 84.955 12.415 85.705 ;
        RECT 12.585 85.160 17.930 85.705 ;
        RECT 18.105 85.160 23.450 85.705 ;
        RECT 23.625 85.160 28.970 85.705 ;
        RECT 29.145 85.160 34.490 85.705 ;
        RECT 11.205 84.415 11.725 84.955 ;
        RECT 11.895 84.245 12.415 84.785 ;
        RECT 14.170 84.330 14.510 85.160 ;
        RECT 11.205 83.155 12.415 84.245 ;
        RECT 15.990 83.590 16.340 84.840 ;
        RECT 19.690 84.330 20.030 85.160 ;
        RECT 21.510 83.590 21.860 84.840 ;
        RECT 25.210 84.330 25.550 85.160 ;
        RECT 27.030 83.590 27.380 84.840 ;
        RECT 30.730 84.330 31.070 85.160 ;
        RECT 34.665 84.935 36.335 85.705 ;
        RECT 36.965 84.980 37.255 85.705 ;
        RECT 37.425 85.160 42.770 85.705 ;
        RECT 42.945 85.160 48.290 85.705 ;
        RECT 48.465 85.160 53.810 85.705 ;
        RECT 53.985 85.160 59.330 85.705 ;
        RECT 32.550 83.590 32.900 84.840 ;
        RECT 34.665 84.415 35.415 84.935 ;
        RECT 35.585 84.245 36.335 84.765 ;
        RECT 39.010 84.330 39.350 85.160 ;
        RECT 12.585 83.155 17.930 83.590 ;
        RECT 18.105 83.155 23.450 83.590 ;
        RECT 23.625 83.155 28.970 83.590 ;
        RECT 29.145 83.155 34.490 83.590 ;
        RECT 34.665 83.155 36.335 84.245 ;
        RECT 36.965 83.155 37.255 84.320 ;
        RECT 40.830 83.590 41.180 84.840 ;
        RECT 44.530 84.330 44.870 85.160 ;
        RECT 46.350 83.590 46.700 84.840 ;
        RECT 50.050 84.330 50.390 85.160 ;
        RECT 51.870 83.590 52.220 84.840 ;
        RECT 55.570 84.330 55.910 85.160 ;
        RECT 59.505 84.935 62.095 85.705 ;
        RECT 62.725 84.980 63.015 85.705 ;
        RECT 63.185 85.160 68.530 85.705 ;
        RECT 68.705 85.160 74.050 85.705 ;
        RECT 74.225 85.160 79.570 85.705 ;
        RECT 79.745 85.160 85.090 85.705 ;
        RECT 57.390 83.590 57.740 84.840 ;
        RECT 59.505 84.415 60.715 84.935 ;
        RECT 60.885 84.245 62.095 84.765 ;
        RECT 64.770 84.330 65.110 85.160 ;
        RECT 37.425 83.155 42.770 83.590 ;
        RECT 42.945 83.155 48.290 83.590 ;
        RECT 48.465 83.155 53.810 83.590 ;
        RECT 53.985 83.155 59.330 83.590 ;
        RECT 59.505 83.155 62.095 84.245 ;
        RECT 62.725 83.155 63.015 84.320 ;
        RECT 66.590 83.590 66.940 84.840 ;
        RECT 70.290 84.330 70.630 85.160 ;
        RECT 72.110 83.590 72.460 84.840 ;
        RECT 75.810 84.330 76.150 85.160 ;
        RECT 77.630 83.590 77.980 84.840 ;
        RECT 81.330 84.330 81.670 85.160 ;
        RECT 85.265 84.935 87.855 85.705 ;
        RECT 88.485 84.980 88.775 85.705 ;
        RECT 88.945 85.160 94.290 85.705 ;
        RECT 94.465 85.160 99.810 85.705 ;
        RECT 99.985 85.160 105.330 85.705 ;
        RECT 105.505 85.160 110.850 85.705 ;
        RECT 83.150 83.590 83.500 84.840 ;
        RECT 85.265 84.415 86.475 84.935 ;
        RECT 86.645 84.245 87.855 84.765 ;
        RECT 90.530 84.330 90.870 85.160 ;
        RECT 63.185 83.155 68.530 83.590 ;
        RECT 68.705 83.155 74.050 83.590 ;
        RECT 74.225 83.155 79.570 83.590 ;
        RECT 79.745 83.155 85.090 83.590 ;
        RECT 85.265 83.155 87.855 84.245 ;
        RECT 88.485 83.155 88.775 84.320 ;
        RECT 92.350 83.590 92.700 84.840 ;
        RECT 96.050 84.330 96.390 85.160 ;
        RECT 97.870 83.590 98.220 84.840 ;
        RECT 101.570 84.330 101.910 85.160 ;
        RECT 103.390 83.590 103.740 84.840 ;
        RECT 107.090 84.330 107.430 85.160 ;
        RECT 111.025 84.935 113.615 85.705 ;
        RECT 114.245 84.980 114.535 85.705 ;
        RECT 114.705 85.160 120.050 85.705 ;
        RECT 120.225 85.160 125.570 85.705 ;
        RECT 125.745 85.160 131.090 85.705 ;
        RECT 131.265 85.160 136.610 85.705 ;
        RECT 108.910 83.590 109.260 84.840 ;
        RECT 111.025 84.415 112.235 84.935 ;
        RECT 112.405 84.245 113.615 84.765 ;
        RECT 116.290 84.330 116.630 85.160 ;
        RECT 88.945 83.155 94.290 83.590 ;
        RECT 94.465 83.155 99.810 83.590 ;
        RECT 99.985 83.155 105.330 83.590 ;
        RECT 105.505 83.155 110.850 83.590 ;
        RECT 111.025 83.155 113.615 84.245 ;
        RECT 114.245 83.155 114.535 84.320 ;
        RECT 118.110 83.590 118.460 84.840 ;
        RECT 121.810 84.330 122.150 85.160 ;
        RECT 123.630 83.590 123.980 84.840 ;
        RECT 127.330 84.330 127.670 85.160 ;
        RECT 129.150 83.590 129.500 84.840 ;
        RECT 132.850 84.330 133.190 85.160 ;
        RECT 136.785 84.935 139.375 85.705 ;
        RECT 140.005 84.980 140.295 85.705 ;
        RECT 140.465 85.160 145.810 85.705 ;
        RECT 134.670 83.590 135.020 84.840 ;
        RECT 136.785 84.415 137.995 84.935 ;
        RECT 138.165 84.245 139.375 84.765 ;
        RECT 142.050 84.330 142.390 85.160 ;
        RECT 145.985 84.935 148.575 85.705 ;
        RECT 149.205 84.955 150.415 85.705 ;
        RECT 114.705 83.155 120.050 83.590 ;
        RECT 120.225 83.155 125.570 83.590 ;
        RECT 125.745 83.155 131.090 83.590 ;
        RECT 131.265 83.155 136.610 83.590 ;
        RECT 136.785 83.155 139.375 84.245 ;
        RECT 140.005 83.155 140.295 84.320 ;
        RECT 143.870 83.590 144.220 84.840 ;
        RECT 145.985 84.415 147.195 84.935 ;
        RECT 147.365 84.245 148.575 84.765 ;
        RECT 140.465 83.155 145.810 83.590 ;
        RECT 145.985 83.155 148.575 84.245 ;
        RECT 149.205 84.245 149.725 84.785 ;
        RECT 149.895 84.415 150.415 84.955 ;
        RECT 149.205 83.155 150.415 84.245 ;
        RECT 11.120 82.985 150.500 83.155 ;
        RECT 11.205 81.895 12.415 82.985 ;
        RECT 12.585 82.550 17.930 82.985 ;
        RECT 18.105 82.550 23.450 82.985 ;
        RECT 11.205 81.185 11.725 81.725 ;
        RECT 11.895 81.355 12.415 81.895 ;
        RECT 11.205 80.435 12.415 81.185 ;
        RECT 14.170 80.980 14.510 81.810 ;
        RECT 15.990 81.300 16.340 82.550 ;
        RECT 19.690 80.980 20.030 81.810 ;
        RECT 21.510 81.300 21.860 82.550 ;
        RECT 24.085 81.820 24.375 82.985 ;
        RECT 24.545 82.550 29.890 82.985 ;
        RECT 30.065 82.550 35.410 82.985 ;
        RECT 35.585 82.550 40.930 82.985 ;
        RECT 41.105 82.550 46.450 82.985 ;
        RECT 12.585 80.435 17.930 80.980 ;
        RECT 18.105 80.435 23.450 80.980 ;
        RECT 24.085 80.435 24.375 81.160 ;
        RECT 26.130 80.980 26.470 81.810 ;
        RECT 27.950 81.300 28.300 82.550 ;
        RECT 31.650 80.980 31.990 81.810 ;
        RECT 33.470 81.300 33.820 82.550 ;
        RECT 37.170 80.980 37.510 81.810 ;
        RECT 38.990 81.300 39.340 82.550 ;
        RECT 42.690 80.980 43.030 81.810 ;
        RECT 44.510 81.300 44.860 82.550 ;
        RECT 46.625 81.895 49.215 82.985 ;
        RECT 46.625 81.205 47.835 81.725 ;
        RECT 48.005 81.375 49.215 81.895 ;
        RECT 49.845 81.820 50.135 82.985 ;
        RECT 50.305 82.550 55.650 82.985 ;
        RECT 55.825 82.550 61.170 82.985 ;
        RECT 61.345 82.550 66.690 82.985 ;
        RECT 66.865 82.550 72.210 82.985 ;
        RECT 24.545 80.435 29.890 80.980 ;
        RECT 30.065 80.435 35.410 80.980 ;
        RECT 35.585 80.435 40.930 80.980 ;
        RECT 41.105 80.435 46.450 80.980 ;
        RECT 46.625 80.435 49.215 81.205 ;
        RECT 49.845 80.435 50.135 81.160 ;
        RECT 51.890 80.980 52.230 81.810 ;
        RECT 53.710 81.300 54.060 82.550 ;
        RECT 57.410 80.980 57.750 81.810 ;
        RECT 59.230 81.300 59.580 82.550 ;
        RECT 62.930 80.980 63.270 81.810 ;
        RECT 64.750 81.300 65.100 82.550 ;
        RECT 68.450 80.980 68.790 81.810 ;
        RECT 70.270 81.300 70.620 82.550 ;
        RECT 72.385 81.895 74.975 82.985 ;
        RECT 72.385 81.205 73.595 81.725 ;
        RECT 73.765 81.375 74.975 81.895 ;
        RECT 75.605 81.820 75.895 82.985 ;
        RECT 76.065 82.550 81.410 82.985 ;
        RECT 81.585 82.550 86.930 82.985 ;
        RECT 87.105 82.550 92.450 82.985 ;
        RECT 92.625 82.550 97.970 82.985 ;
        RECT 50.305 80.435 55.650 80.980 ;
        RECT 55.825 80.435 61.170 80.980 ;
        RECT 61.345 80.435 66.690 80.980 ;
        RECT 66.865 80.435 72.210 80.980 ;
        RECT 72.385 80.435 74.975 81.205 ;
        RECT 75.605 80.435 75.895 81.160 ;
        RECT 77.650 80.980 77.990 81.810 ;
        RECT 79.470 81.300 79.820 82.550 ;
        RECT 83.170 80.980 83.510 81.810 ;
        RECT 84.990 81.300 85.340 82.550 ;
        RECT 88.690 80.980 89.030 81.810 ;
        RECT 90.510 81.300 90.860 82.550 ;
        RECT 94.210 80.980 94.550 81.810 ;
        RECT 96.030 81.300 96.380 82.550 ;
        RECT 98.145 81.895 100.735 82.985 ;
        RECT 98.145 81.205 99.355 81.725 ;
        RECT 99.525 81.375 100.735 81.895 ;
        RECT 101.365 81.820 101.655 82.985 ;
        RECT 101.825 82.550 107.170 82.985 ;
        RECT 107.345 82.550 112.690 82.985 ;
        RECT 112.865 82.550 118.210 82.985 ;
        RECT 118.385 82.550 123.730 82.985 ;
        RECT 76.065 80.435 81.410 80.980 ;
        RECT 81.585 80.435 86.930 80.980 ;
        RECT 87.105 80.435 92.450 80.980 ;
        RECT 92.625 80.435 97.970 80.980 ;
        RECT 98.145 80.435 100.735 81.205 ;
        RECT 101.365 80.435 101.655 81.160 ;
        RECT 103.410 80.980 103.750 81.810 ;
        RECT 105.230 81.300 105.580 82.550 ;
        RECT 108.930 80.980 109.270 81.810 ;
        RECT 110.750 81.300 111.100 82.550 ;
        RECT 114.450 80.980 114.790 81.810 ;
        RECT 116.270 81.300 116.620 82.550 ;
        RECT 119.970 80.980 120.310 81.810 ;
        RECT 121.790 81.300 122.140 82.550 ;
        RECT 123.905 81.895 126.495 82.985 ;
        RECT 123.905 81.205 125.115 81.725 ;
        RECT 125.285 81.375 126.495 81.895 ;
        RECT 127.125 81.820 127.415 82.985 ;
        RECT 127.585 82.550 132.930 82.985 ;
        RECT 133.105 82.550 138.450 82.985 ;
        RECT 138.625 82.550 143.970 82.985 ;
        RECT 101.825 80.435 107.170 80.980 ;
        RECT 107.345 80.435 112.690 80.980 ;
        RECT 112.865 80.435 118.210 80.980 ;
        RECT 118.385 80.435 123.730 80.980 ;
        RECT 123.905 80.435 126.495 81.205 ;
        RECT 127.125 80.435 127.415 81.160 ;
        RECT 129.170 80.980 129.510 81.810 ;
        RECT 130.990 81.300 131.340 82.550 ;
        RECT 134.690 80.980 135.030 81.810 ;
        RECT 136.510 81.300 136.860 82.550 ;
        RECT 140.210 80.980 140.550 81.810 ;
        RECT 142.030 81.300 142.380 82.550 ;
        RECT 144.145 81.895 147.655 82.985 ;
        RECT 147.825 81.895 149.035 82.985 ;
        RECT 144.145 81.205 145.795 81.725 ;
        RECT 145.965 81.375 147.655 81.895 ;
        RECT 127.585 80.435 132.930 80.980 ;
        RECT 133.105 80.435 138.450 80.980 ;
        RECT 138.625 80.435 143.970 80.980 ;
        RECT 144.145 80.435 147.655 81.205 ;
        RECT 147.825 81.185 148.345 81.725 ;
        RECT 148.515 81.355 149.035 81.895 ;
        RECT 149.205 81.895 150.415 82.985 ;
        RECT 149.205 81.355 149.725 81.895 ;
        RECT 149.895 81.185 150.415 81.725 ;
        RECT 147.825 80.435 149.035 81.185 ;
        RECT 149.205 80.435 150.415 81.185 ;
        RECT 11.120 80.265 150.500 80.435 ;
        RECT 11.205 79.515 12.415 80.265 ;
        RECT 12.585 79.720 17.930 80.265 ;
        RECT 18.105 79.720 23.450 80.265 ;
        RECT 23.625 79.720 28.970 80.265 ;
        RECT 29.145 79.720 34.490 80.265 ;
        RECT 11.205 78.975 11.725 79.515 ;
        RECT 11.895 78.805 12.415 79.345 ;
        RECT 14.170 78.890 14.510 79.720 ;
        RECT 11.205 77.715 12.415 78.805 ;
        RECT 15.990 78.150 16.340 79.400 ;
        RECT 19.690 78.890 20.030 79.720 ;
        RECT 21.510 78.150 21.860 79.400 ;
        RECT 25.210 78.890 25.550 79.720 ;
        RECT 27.030 78.150 27.380 79.400 ;
        RECT 30.730 78.890 31.070 79.720 ;
        RECT 34.665 79.495 36.335 80.265 ;
        RECT 36.965 79.540 37.255 80.265 ;
        RECT 37.425 79.720 42.770 80.265 ;
        RECT 42.945 79.720 48.290 80.265 ;
        RECT 48.465 79.720 53.810 80.265 ;
        RECT 53.985 79.720 59.330 80.265 ;
        RECT 32.550 78.150 32.900 79.400 ;
        RECT 34.665 78.975 35.415 79.495 ;
        RECT 35.585 78.805 36.335 79.325 ;
        RECT 39.010 78.890 39.350 79.720 ;
        RECT 12.585 77.715 17.930 78.150 ;
        RECT 18.105 77.715 23.450 78.150 ;
        RECT 23.625 77.715 28.970 78.150 ;
        RECT 29.145 77.715 34.490 78.150 ;
        RECT 34.665 77.715 36.335 78.805 ;
        RECT 36.965 77.715 37.255 78.880 ;
        RECT 40.830 78.150 41.180 79.400 ;
        RECT 44.530 78.890 44.870 79.720 ;
        RECT 46.350 78.150 46.700 79.400 ;
        RECT 50.050 78.890 50.390 79.720 ;
        RECT 51.870 78.150 52.220 79.400 ;
        RECT 55.570 78.890 55.910 79.720 ;
        RECT 59.505 79.495 62.095 80.265 ;
        RECT 62.725 79.540 63.015 80.265 ;
        RECT 63.185 79.720 68.530 80.265 ;
        RECT 68.705 79.720 74.050 80.265 ;
        RECT 74.225 79.720 79.570 80.265 ;
        RECT 79.745 79.720 85.090 80.265 ;
        RECT 57.390 78.150 57.740 79.400 ;
        RECT 59.505 78.975 60.715 79.495 ;
        RECT 60.885 78.805 62.095 79.325 ;
        RECT 64.770 78.890 65.110 79.720 ;
        RECT 37.425 77.715 42.770 78.150 ;
        RECT 42.945 77.715 48.290 78.150 ;
        RECT 48.465 77.715 53.810 78.150 ;
        RECT 53.985 77.715 59.330 78.150 ;
        RECT 59.505 77.715 62.095 78.805 ;
        RECT 62.725 77.715 63.015 78.880 ;
        RECT 66.590 78.150 66.940 79.400 ;
        RECT 70.290 78.890 70.630 79.720 ;
        RECT 72.110 78.150 72.460 79.400 ;
        RECT 75.810 78.890 76.150 79.720 ;
        RECT 77.630 78.150 77.980 79.400 ;
        RECT 81.330 78.890 81.670 79.720 ;
        RECT 85.265 79.495 87.855 80.265 ;
        RECT 88.485 79.540 88.775 80.265 ;
        RECT 88.945 79.720 94.290 80.265 ;
        RECT 94.465 79.720 99.810 80.265 ;
        RECT 99.985 79.720 105.330 80.265 ;
        RECT 105.505 79.720 110.850 80.265 ;
        RECT 83.150 78.150 83.500 79.400 ;
        RECT 85.265 78.975 86.475 79.495 ;
        RECT 86.645 78.805 87.855 79.325 ;
        RECT 90.530 78.890 90.870 79.720 ;
        RECT 63.185 77.715 68.530 78.150 ;
        RECT 68.705 77.715 74.050 78.150 ;
        RECT 74.225 77.715 79.570 78.150 ;
        RECT 79.745 77.715 85.090 78.150 ;
        RECT 85.265 77.715 87.855 78.805 ;
        RECT 88.485 77.715 88.775 78.880 ;
        RECT 92.350 78.150 92.700 79.400 ;
        RECT 96.050 78.890 96.390 79.720 ;
        RECT 97.870 78.150 98.220 79.400 ;
        RECT 101.570 78.890 101.910 79.720 ;
        RECT 103.390 78.150 103.740 79.400 ;
        RECT 107.090 78.890 107.430 79.720 ;
        RECT 111.025 79.495 113.615 80.265 ;
        RECT 114.245 79.540 114.535 80.265 ;
        RECT 114.705 79.720 120.050 80.265 ;
        RECT 120.225 79.720 125.570 80.265 ;
        RECT 125.745 79.720 131.090 80.265 ;
        RECT 131.265 79.720 136.610 80.265 ;
        RECT 108.910 78.150 109.260 79.400 ;
        RECT 111.025 78.975 112.235 79.495 ;
        RECT 112.405 78.805 113.615 79.325 ;
        RECT 116.290 78.890 116.630 79.720 ;
        RECT 88.945 77.715 94.290 78.150 ;
        RECT 94.465 77.715 99.810 78.150 ;
        RECT 99.985 77.715 105.330 78.150 ;
        RECT 105.505 77.715 110.850 78.150 ;
        RECT 111.025 77.715 113.615 78.805 ;
        RECT 114.245 77.715 114.535 78.880 ;
        RECT 118.110 78.150 118.460 79.400 ;
        RECT 121.810 78.890 122.150 79.720 ;
        RECT 123.630 78.150 123.980 79.400 ;
        RECT 127.330 78.890 127.670 79.720 ;
        RECT 129.150 78.150 129.500 79.400 ;
        RECT 132.850 78.890 133.190 79.720 ;
        RECT 136.785 79.495 139.375 80.265 ;
        RECT 140.005 79.540 140.295 80.265 ;
        RECT 140.465 79.720 145.810 80.265 ;
        RECT 134.670 78.150 135.020 79.400 ;
        RECT 136.785 78.975 137.995 79.495 ;
        RECT 138.165 78.805 139.375 79.325 ;
        RECT 142.050 78.890 142.390 79.720 ;
        RECT 145.985 79.495 148.575 80.265 ;
        RECT 149.205 79.515 150.415 80.265 ;
        RECT 114.705 77.715 120.050 78.150 ;
        RECT 120.225 77.715 125.570 78.150 ;
        RECT 125.745 77.715 131.090 78.150 ;
        RECT 131.265 77.715 136.610 78.150 ;
        RECT 136.785 77.715 139.375 78.805 ;
        RECT 140.005 77.715 140.295 78.880 ;
        RECT 143.870 78.150 144.220 79.400 ;
        RECT 145.985 78.975 147.195 79.495 ;
        RECT 147.365 78.805 148.575 79.325 ;
        RECT 140.465 77.715 145.810 78.150 ;
        RECT 145.985 77.715 148.575 78.805 ;
        RECT 149.205 78.805 149.725 79.345 ;
        RECT 149.895 78.975 150.415 79.515 ;
        RECT 149.205 77.715 150.415 78.805 ;
        RECT 11.120 77.545 150.500 77.715 ;
        RECT 11.205 76.455 12.415 77.545 ;
        RECT 12.585 77.110 17.930 77.545 ;
        RECT 18.105 77.110 23.450 77.545 ;
        RECT 11.205 75.745 11.725 76.285 ;
        RECT 11.895 75.915 12.415 76.455 ;
        RECT 11.205 74.995 12.415 75.745 ;
        RECT 14.170 75.540 14.510 76.370 ;
        RECT 15.990 75.860 16.340 77.110 ;
        RECT 19.690 75.540 20.030 76.370 ;
        RECT 21.510 75.860 21.860 77.110 ;
        RECT 24.085 76.380 24.375 77.545 ;
        RECT 24.545 77.110 29.890 77.545 ;
        RECT 30.065 77.110 35.410 77.545 ;
        RECT 12.585 74.995 17.930 75.540 ;
        RECT 18.105 74.995 23.450 75.540 ;
        RECT 24.085 74.995 24.375 75.720 ;
        RECT 26.130 75.540 26.470 76.370 ;
        RECT 27.950 75.860 28.300 77.110 ;
        RECT 31.650 75.540 31.990 76.370 ;
        RECT 33.470 75.860 33.820 77.110 ;
        RECT 35.585 76.455 36.795 77.545 ;
        RECT 35.585 75.745 36.105 76.285 ;
        RECT 36.275 75.915 36.795 76.455 ;
        RECT 36.965 76.380 37.255 77.545 ;
        RECT 37.425 77.110 42.770 77.545 ;
        RECT 42.945 77.110 48.290 77.545 ;
        RECT 24.545 74.995 29.890 75.540 ;
        RECT 30.065 74.995 35.410 75.540 ;
        RECT 35.585 74.995 36.795 75.745 ;
        RECT 36.965 74.995 37.255 75.720 ;
        RECT 39.010 75.540 39.350 76.370 ;
        RECT 40.830 75.860 41.180 77.110 ;
        RECT 44.530 75.540 44.870 76.370 ;
        RECT 46.350 75.860 46.700 77.110 ;
        RECT 48.465 76.455 49.675 77.545 ;
        RECT 48.465 75.745 48.985 76.285 ;
        RECT 49.155 75.915 49.675 76.455 ;
        RECT 49.845 76.380 50.135 77.545 ;
        RECT 50.305 77.110 55.650 77.545 ;
        RECT 55.825 77.110 61.170 77.545 ;
        RECT 37.425 74.995 42.770 75.540 ;
        RECT 42.945 74.995 48.290 75.540 ;
        RECT 48.465 74.995 49.675 75.745 ;
        RECT 49.845 74.995 50.135 75.720 ;
        RECT 51.890 75.540 52.230 76.370 ;
        RECT 53.710 75.860 54.060 77.110 ;
        RECT 57.410 75.540 57.750 76.370 ;
        RECT 59.230 75.860 59.580 77.110 ;
        RECT 61.345 76.455 62.555 77.545 ;
        RECT 61.345 75.745 61.865 76.285 ;
        RECT 62.035 75.915 62.555 76.455 ;
        RECT 62.725 76.380 63.015 77.545 ;
        RECT 63.185 77.110 68.530 77.545 ;
        RECT 68.705 77.110 74.050 77.545 ;
        RECT 50.305 74.995 55.650 75.540 ;
        RECT 55.825 74.995 61.170 75.540 ;
        RECT 61.345 74.995 62.555 75.745 ;
        RECT 62.725 74.995 63.015 75.720 ;
        RECT 64.770 75.540 65.110 76.370 ;
        RECT 66.590 75.860 66.940 77.110 ;
        RECT 70.290 75.540 70.630 76.370 ;
        RECT 72.110 75.860 72.460 77.110 ;
        RECT 74.225 76.455 75.435 77.545 ;
        RECT 74.225 75.745 74.745 76.285 ;
        RECT 74.915 75.915 75.435 76.455 ;
        RECT 75.605 76.380 75.895 77.545 ;
        RECT 76.065 77.110 81.410 77.545 ;
        RECT 81.585 77.110 86.930 77.545 ;
        RECT 63.185 74.995 68.530 75.540 ;
        RECT 68.705 74.995 74.050 75.540 ;
        RECT 74.225 74.995 75.435 75.745 ;
        RECT 75.605 74.995 75.895 75.720 ;
        RECT 77.650 75.540 77.990 76.370 ;
        RECT 79.470 75.860 79.820 77.110 ;
        RECT 83.170 75.540 83.510 76.370 ;
        RECT 84.990 75.860 85.340 77.110 ;
        RECT 87.105 76.455 88.315 77.545 ;
        RECT 87.105 75.745 87.625 76.285 ;
        RECT 87.795 75.915 88.315 76.455 ;
        RECT 88.485 76.380 88.775 77.545 ;
        RECT 88.945 77.110 94.290 77.545 ;
        RECT 94.465 77.110 99.810 77.545 ;
        RECT 76.065 74.995 81.410 75.540 ;
        RECT 81.585 74.995 86.930 75.540 ;
        RECT 87.105 74.995 88.315 75.745 ;
        RECT 88.485 74.995 88.775 75.720 ;
        RECT 90.530 75.540 90.870 76.370 ;
        RECT 92.350 75.860 92.700 77.110 ;
        RECT 96.050 75.540 96.390 76.370 ;
        RECT 97.870 75.860 98.220 77.110 ;
        RECT 99.985 76.455 101.195 77.545 ;
        RECT 99.985 75.745 100.505 76.285 ;
        RECT 100.675 75.915 101.195 76.455 ;
        RECT 101.365 76.380 101.655 77.545 ;
        RECT 101.825 77.110 107.170 77.545 ;
        RECT 107.345 77.110 112.690 77.545 ;
        RECT 88.945 74.995 94.290 75.540 ;
        RECT 94.465 74.995 99.810 75.540 ;
        RECT 99.985 74.995 101.195 75.745 ;
        RECT 101.365 74.995 101.655 75.720 ;
        RECT 103.410 75.540 103.750 76.370 ;
        RECT 105.230 75.860 105.580 77.110 ;
        RECT 108.930 75.540 109.270 76.370 ;
        RECT 110.750 75.860 111.100 77.110 ;
        RECT 112.865 76.455 114.075 77.545 ;
        RECT 112.865 75.745 113.385 76.285 ;
        RECT 113.555 75.915 114.075 76.455 ;
        RECT 114.245 76.380 114.535 77.545 ;
        RECT 114.705 77.110 120.050 77.545 ;
        RECT 120.225 77.110 125.570 77.545 ;
        RECT 101.825 74.995 107.170 75.540 ;
        RECT 107.345 74.995 112.690 75.540 ;
        RECT 112.865 74.995 114.075 75.745 ;
        RECT 114.245 74.995 114.535 75.720 ;
        RECT 116.290 75.540 116.630 76.370 ;
        RECT 118.110 75.860 118.460 77.110 ;
        RECT 121.810 75.540 122.150 76.370 ;
        RECT 123.630 75.860 123.980 77.110 ;
        RECT 125.745 76.455 126.955 77.545 ;
        RECT 125.745 75.745 126.265 76.285 ;
        RECT 126.435 75.915 126.955 76.455 ;
        RECT 127.125 76.380 127.415 77.545 ;
        RECT 127.585 77.110 132.930 77.545 ;
        RECT 133.105 77.110 138.450 77.545 ;
        RECT 114.705 74.995 120.050 75.540 ;
        RECT 120.225 74.995 125.570 75.540 ;
        RECT 125.745 74.995 126.955 75.745 ;
        RECT 127.125 74.995 127.415 75.720 ;
        RECT 129.170 75.540 129.510 76.370 ;
        RECT 130.990 75.860 131.340 77.110 ;
        RECT 134.690 75.540 135.030 76.370 ;
        RECT 136.510 75.860 136.860 77.110 ;
        RECT 138.625 76.455 139.835 77.545 ;
        RECT 138.625 75.745 139.145 76.285 ;
        RECT 139.315 75.915 139.835 76.455 ;
        RECT 140.005 76.380 140.295 77.545 ;
        RECT 140.465 77.110 145.810 77.545 ;
        RECT 127.585 74.995 132.930 75.540 ;
        RECT 133.105 74.995 138.450 75.540 ;
        RECT 138.625 74.995 139.835 75.745 ;
        RECT 140.005 74.995 140.295 75.720 ;
        RECT 142.050 75.540 142.390 76.370 ;
        RECT 143.870 75.860 144.220 77.110 ;
        RECT 145.985 76.455 148.575 77.545 ;
        RECT 145.985 75.765 147.195 76.285 ;
        RECT 147.365 75.935 148.575 76.455 ;
        RECT 149.205 76.455 150.415 77.545 ;
        RECT 149.205 75.915 149.725 76.455 ;
        RECT 140.465 74.995 145.810 75.540 ;
        RECT 145.985 74.995 148.575 75.765 ;
        RECT 149.895 75.745 150.415 76.285 ;
        RECT 149.205 74.995 150.415 75.745 ;
        RECT 11.120 74.825 150.500 74.995 ;
        RECT 54.840 49.890 84.840 52.430 ;
        RECT 94.360 50.340 106.510 51.780 ;
        RECT 54.840 35.180 61.230 49.890 ;
        RECT 61.955 49.320 62.995 49.490 ;
        RECT 61.570 47.260 61.740 49.260 ;
        RECT 63.210 47.260 63.380 49.260 ;
        RECT 61.955 47.030 62.995 47.200 ;
        RECT 61.570 44.970 61.740 46.970 ;
        RECT 63.210 44.970 63.380 46.970 ;
        RECT 61.955 44.740 62.995 44.910 ;
        RECT 61.570 42.680 61.740 44.680 ;
        RECT 63.210 42.680 63.380 44.680 ;
        RECT 61.955 42.450 62.995 42.620 ;
        RECT 61.570 40.390 61.740 42.390 ;
        RECT 63.210 40.390 63.380 42.390 ;
        RECT 61.955 40.160 62.995 40.330 ;
        RECT 61.570 38.100 61.740 40.100 ;
        RECT 63.210 38.100 63.380 40.100 ;
        RECT 61.955 37.870 62.995 38.040 ;
        RECT 61.570 35.810 61.740 37.810 ;
        RECT 63.210 35.810 63.380 37.810 ;
        RECT 61.955 35.580 62.995 35.750 ;
        RECT 63.720 35.180 63.890 49.890 ;
        RECT 66.380 49.880 84.840 49.890 ;
        RECT 64.615 49.320 65.655 49.490 ;
        RECT 64.230 47.260 64.400 49.260 ;
        RECT 65.870 47.260 66.040 49.260 ;
        RECT 64.615 47.030 65.655 47.200 ;
        RECT 64.230 44.970 64.400 46.970 ;
        RECT 65.870 44.970 66.040 46.970 ;
        RECT 64.615 44.740 65.655 44.910 ;
        RECT 64.230 42.680 64.400 44.680 ;
        RECT 65.870 42.680 66.040 44.680 ;
        RECT 66.380 43.690 78.000 49.880 ;
        RECT 78.725 49.310 79.765 49.480 ;
        RECT 78.340 48.750 78.510 49.250 ;
        RECT 79.980 48.750 80.150 49.250 ;
        RECT 78.725 48.520 79.765 48.690 ;
        RECT 78.340 47.960 78.510 48.460 ;
        RECT 79.980 47.960 80.150 48.460 ;
        RECT 78.725 47.730 79.765 47.900 ;
        RECT 78.340 47.170 78.510 47.670 ;
        RECT 79.980 47.170 80.150 47.670 ;
        RECT 78.725 46.940 79.765 47.110 ;
        RECT 78.340 46.380 78.510 46.880 ;
        RECT 79.980 46.380 80.150 46.880 ;
        RECT 78.725 46.150 79.765 46.320 ;
        RECT 78.340 45.590 78.510 46.090 ;
        RECT 79.980 45.590 80.150 46.090 ;
        RECT 78.725 45.360 79.765 45.530 ;
        RECT 78.340 44.800 78.510 45.300 ;
        RECT 79.980 44.800 80.150 45.300 ;
        RECT 78.725 44.570 79.765 44.740 ;
        RECT 78.340 44.010 78.510 44.510 ;
        RECT 79.980 44.010 80.150 44.510 ;
        RECT 78.725 43.780 79.765 43.950 ;
        RECT 64.615 42.450 65.655 42.620 ;
        RECT 64.230 40.390 64.400 42.390 ;
        RECT 65.870 40.390 66.040 42.390 ;
        RECT 64.615 40.160 65.655 40.330 ;
        RECT 64.230 38.100 64.400 40.100 ;
        RECT 65.870 38.100 66.040 40.100 ;
        RECT 64.615 37.870 65.655 38.040 ;
        RECT 64.230 35.810 64.400 37.810 ;
        RECT 65.870 35.810 66.040 37.810 ;
        RECT 64.615 35.580 65.655 35.750 ;
        RECT 66.380 35.180 71.810 43.690 ;
        RECT 54.840 34.810 71.810 35.180 ;
        RECT 72.690 42.720 75.430 42.890 ;
        RECT 54.840 34.800 71.660 34.810 ;
        RECT 72.690 34.280 72.860 42.720 ;
        RECT 73.540 42.150 74.580 42.320 ;
        RECT 73.200 40.090 73.370 42.090 ;
        RECT 74.750 40.090 74.920 42.090 ;
        RECT 73.540 39.860 74.580 40.030 ;
        RECT 73.200 37.800 73.370 39.800 ;
        RECT 74.750 37.800 74.920 39.800 ;
        RECT 73.540 37.570 74.580 37.740 ;
        RECT 73.200 35.510 73.370 37.510 ;
        RECT 74.750 35.510 74.920 37.510 ;
        RECT 73.540 35.280 74.580 35.450 ;
        RECT 54.840 34.110 72.860 34.280 ;
        RECT 54.840 30.210 61.940 34.110 ;
        RECT 62.570 33.600 63.070 33.770 ;
        RECT 62.340 30.890 62.510 33.430 ;
        RECT 63.130 30.890 63.300 33.430 ;
        RECT 62.570 30.550 63.070 30.720 ;
        RECT 63.700 30.210 63.870 34.110 ;
        RECT 64.500 33.600 65.000 33.770 ;
        RECT 64.270 30.890 64.440 33.430 ;
        RECT 65.060 30.890 65.230 33.430 ;
        RECT 64.500 30.550 65.000 30.720 ;
        RECT 65.630 30.210 72.860 34.110 ;
        RECT 73.200 33.220 73.370 35.220 ;
        RECT 74.750 33.220 74.920 35.220 ;
        RECT 73.540 32.990 74.580 33.160 ;
        RECT 73.200 30.930 73.370 32.930 ;
        RECT 74.750 30.930 74.920 32.930 ;
        RECT 75.260 31.730 75.430 42.720 ;
        RECT 76.330 33.220 78.000 43.690 ;
        RECT 78.340 43.220 78.510 43.720 ;
        RECT 79.980 43.220 80.150 43.720 ;
        RECT 78.725 42.990 79.765 43.160 ;
        RECT 78.340 42.430 78.510 42.930 ;
        RECT 79.980 42.430 80.150 42.930 ;
        RECT 78.725 42.200 79.765 42.370 ;
        RECT 78.340 41.640 78.510 42.140 ;
        RECT 79.980 41.640 80.150 42.140 ;
        RECT 78.725 41.410 79.765 41.580 ;
        RECT 78.340 40.850 78.510 41.350 ;
        RECT 79.980 40.850 80.150 41.350 ;
        RECT 78.725 40.620 79.765 40.790 ;
        RECT 78.340 40.060 78.510 40.560 ;
        RECT 79.980 40.060 80.150 40.560 ;
        RECT 78.725 39.830 79.765 40.000 ;
        RECT 78.340 39.270 78.510 39.770 ;
        RECT 79.980 39.270 80.150 39.770 ;
        RECT 78.725 39.040 79.765 39.210 ;
        RECT 78.340 38.480 78.510 38.980 ;
        RECT 79.980 38.480 80.150 38.980 ;
        RECT 78.725 38.250 79.765 38.420 ;
        RECT 78.340 37.690 78.510 38.190 ;
        RECT 79.980 37.690 80.150 38.190 ;
        RECT 78.725 37.460 79.765 37.630 ;
        RECT 78.340 36.900 78.510 37.400 ;
        RECT 79.980 36.900 80.150 37.400 ;
        RECT 78.725 36.670 79.765 36.840 ;
        RECT 78.340 36.110 78.510 36.610 ;
        RECT 79.980 36.110 80.150 36.610 ;
        RECT 78.725 35.880 79.765 36.050 ;
        RECT 78.340 35.320 78.510 35.820 ;
        RECT 79.980 35.320 80.150 35.820 ;
        RECT 78.725 35.090 79.765 35.260 ;
        RECT 78.340 34.530 78.510 35.030 ;
        RECT 79.980 34.530 80.150 35.030 ;
        RECT 78.725 34.300 79.765 34.470 ;
        RECT 78.340 33.740 78.510 34.240 ;
        RECT 79.980 33.740 80.150 34.240 ;
        RECT 78.725 33.510 79.765 33.680 ;
        RECT 80.490 33.220 84.840 49.880 ;
        RECT 94.380 49.800 99.650 49.870 ;
        RECT 101.120 49.800 106.490 49.810 ;
        RECT 94.380 49.630 106.490 49.800 ;
        RECT 94.380 41.710 99.750 49.630 ;
        RECT 100.230 46.990 100.580 49.150 ;
        RECT 100.230 42.190 100.580 44.350 ;
        RECT 101.060 41.710 106.490 49.630 ;
        RECT 94.380 39.790 106.490 41.710 ;
        RECT 94.380 37.390 95.140 39.790 ;
        RECT 95.770 39.280 97.770 39.450 ;
        RECT 98.060 39.280 100.060 39.450 ;
        RECT 100.350 39.280 102.350 39.450 ;
        RECT 102.640 39.280 104.640 39.450 ;
        RECT 95.540 38.070 95.710 39.110 ;
        RECT 97.830 38.070 98.000 39.110 ;
        RECT 100.120 38.070 100.290 39.110 ;
        RECT 102.410 38.070 102.580 39.110 ;
        RECT 104.700 38.070 104.870 39.110 ;
        RECT 95.770 37.730 97.770 37.900 ;
        RECT 98.060 37.730 100.060 37.900 ;
        RECT 100.350 37.730 102.350 37.900 ;
        RECT 102.640 37.730 104.640 37.900 ;
        RECT 105.270 37.390 106.490 39.790 ;
        RECT 94.380 36.810 106.490 37.390 ;
        RECT 94.360 35.380 106.490 36.810 ;
        RECT 94.340 34.100 106.490 35.380 ;
        RECT 117.070 49.490 147.070 52.030 ;
        RECT 117.070 34.780 123.460 49.490 ;
        RECT 124.185 48.920 125.225 49.090 ;
        RECT 123.800 46.860 123.970 48.860 ;
        RECT 125.440 46.860 125.610 48.860 ;
        RECT 124.185 46.630 125.225 46.800 ;
        RECT 123.800 44.570 123.970 46.570 ;
        RECT 125.440 44.570 125.610 46.570 ;
        RECT 124.185 44.340 125.225 44.510 ;
        RECT 123.800 42.280 123.970 44.280 ;
        RECT 125.440 42.280 125.610 44.280 ;
        RECT 124.185 42.050 125.225 42.220 ;
        RECT 123.800 39.990 123.970 41.990 ;
        RECT 125.440 39.990 125.610 41.990 ;
        RECT 124.185 39.760 125.225 39.930 ;
        RECT 123.800 37.700 123.970 39.700 ;
        RECT 125.440 37.700 125.610 39.700 ;
        RECT 124.185 37.470 125.225 37.640 ;
        RECT 123.800 35.410 123.970 37.410 ;
        RECT 125.440 35.410 125.610 37.410 ;
        RECT 124.185 35.180 125.225 35.350 ;
        RECT 125.950 34.780 126.120 49.490 ;
        RECT 128.610 49.480 147.070 49.490 ;
        RECT 126.845 48.920 127.885 49.090 ;
        RECT 126.460 46.860 126.630 48.860 ;
        RECT 128.100 46.860 128.270 48.860 ;
        RECT 126.845 46.630 127.885 46.800 ;
        RECT 126.460 44.570 126.630 46.570 ;
        RECT 128.100 44.570 128.270 46.570 ;
        RECT 126.845 44.340 127.885 44.510 ;
        RECT 126.460 42.280 126.630 44.280 ;
        RECT 128.100 42.280 128.270 44.280 ;
        RECT 128.610 43.290 140.230 49.480 ;
        RECT 140.955 48.910 141.995 49.080 ;
        RECT 140.570 48.350 140.740 48.850 ;
        RECT 142.210 48.350 142.380 48.850 ;
        RECT 140.955 48.120 141.995 48.290 ;
        RECT 140.570 47.560 140.740 48.060 ;
        RECT 142.210 47.560 142.380 48.060 ;
        RECT 140.955 47.330 141.995 47.500 ;
        RECT 140.570 46.770 140.740 47.270 ;
        RECT 142.210 46.770 142.380 47.270 ;
        RECT 140.955 46.540 141.995 46.710 ;
        RECT 140.570 45.980 140.740 46.480 ;
        RECT 142.210 45.980 142.380 46.480 ;
        RECT 140.955 45.750 141.995 45.920 ;
        RECT 140.570 45.190 140.740 45.690 ;
        RECT 142.210 45.190 142.380 45.690 ;
        RECT 140.955 44.960 141.995 45.130 ;
        RECT 140.570 44.400 140.740 44.900 ;
        RECT 142.210 44.400 142.380 44.900 ;
        RECT 140.955 44.170 141.995 44.340 ;
        RECT 140.570 43.610 140.740 44.110 ;
        RECT 142.210 43.610 142.380 44.110 ;
        RECT 140.955 43.380 141.995 43.550 ;
        RECT 126.845 42.050 127.885 42.220 ;
        RECT 126.460 39.990 126.630 41.990 ;
        RECT 128.100 39.990 128.270 41.990 ;
        RECT 126.845 39.760 127.885 39.930 ;
        RECT 126.460 37.700 126.630 39.700 ;
        RECT 128.100 37.700 128.270 39.700 ;
        RECT 126.845 37.470 127.885 37.640 ;
        RECT 126.460 35.410 126.630 37.410 ;
        RECT 128.100 35.410 128.270 37.410 ;
        RECT 126.845 35.180 127.885 35.350 ;
        RECT 128.610 34.780 134.040 43.290 ;
        RECT 117.070 34.410 134.040 34.780 ;
        RECT 134.920 42.320 137.660 42.490 ;
        RECT 117.070 34.400 133.890 34.410 ;
        RECT 134.920 33.880 135.090 42.320 ;
        RECT 135.770 41.750 136.810 41.920 ;
        RECT 135.430 39.690 135.600 41.690 ;
        RECT 136.980 39.690 137.150 41.690 ;
        RECT 135.770 39.460 136.810 39.630 ;
        RECT 135.430 37.400 135.600 39.400 ;
        RECT 136.980 37.400 137.150 39.400 ;
        RECT 135.770 37.170 136.810 37.340 ;
        RECT 135.430 35.110 135.600 37.110 ;
        RECT 136.980 35.110 137.150 37.110 ;
        RECT 135.770 34.880 136.810 35.050 ;
        RECT 76.330 32.690 84.840 33.220 ;
        RECT 117.070 33.710 135.090 33.880 ;
        RECT 73.540 30.700 74.580 30.870 ;
        RECT 54.840 27.170 72.860 30.210 ;
        RECT 73.200 28.640 73.370 30.640 ;
        RECT 74.750 28.640 74.920 30.640 ;
        RECT 73.540 28.410 74.580 28.580 ;
        RECT 54.840 24.770 55.200 27.170 ;
        RECT 55.830 26.660 57.830 26.830 ;
        RECT 58.120 26.660 60.120 26.830 ;
        RECT 60.410 26.660 62.410 26.830 ;
        RECT 62.700 26.660 64.700 26.830 ;
        RECT 55.600 25.450 55.770 26.490 ;
        RECT 57.890 25.450 58.060 26.490 ;
        RECT 60.180 25.450 60.350 26.490 ;
        RECT 62.470 25.450 62.640 26.490 ;
        RECT 64.760 25.450 64.930 26.490 ;
        RECT 65.330 25.720 72.860 27.170 ;
        RECT 73.200 26.350 73.370 28.350 ;
        RECT 74.750 26.350 74.920 28.350 ;
        RECT 73.540 26.120 74.580 26.290 ;
        RECT 75.260 25.720 84.840 31.730 ;
        RECT 55.830 25.110 57.830 25.280 ;
        RECT 58.120 25.110 60.120 25.280 ;
        RECT 60.410 25.110 62.410 25.280 ;
        RECT 62.700 25.110 64.700 25.280 ;
        RECT 65.330 24.770 84.840 25.720 ;
        RECT 54.840 22.450 84.840 24.770 ;
        RECT 117.070 29.810 124.170 33.710 ;
        RECT 124.800 33.200 125.300 33.370 ;
        RECT 124.570 30.490 124.740 33.030 ;
        RECT 125.360 30.490 125.530 33.030 ;
        RECT 124.800 30.150 125.300 30.320 ;
        RECT 125.930 29.810 126.100 33.710 ;
        RECT 126.730 33.200 127.230 33.370 ;
        RECT 126.500 30.490 126.670 33.030 ;
        RECT 127.290 30.490 127.460 33.030 ;
        RECT 126.730 30.150 127.230 30.320 ;
        RECT 127.860 29.810 135.090 33.710 ;
        RECT 135.430 32.820 135.600 34.820 ;
        RECT 136.980 32.820 137.150 34.820 ;
        RECT 135.770 32.590 136.810 32.760 ;
        RECT 135.430 30.530 135.600 32.530 ;
        RECT 136.980 30.530 137.150 32.530 ;
        RECT 137.490 31.330 137.660 42.320 ;
        RECT 138.560 32.820 140.230 43.290 ;
        RECT 140.570 42.820 140.740 43.320 ;
        RECT 142.210 42.820 142.380 43.320 ;
        RECT 140.955 42.590 141.995 42.760 ;
        RECT 140.570 42.030 140.740 42.530 ;
        RECT 142.210 42.030 142.380 42.530 ;
        RECT 140.955 41.800 141.995 41.970 ;
        RECT 140.570 41.240 140.740 41.740 ;
        RECT 142.210 41.240 142.380 41.740 ;
        RECT 140.955 41.010 141.995 41.180 ;
        RECT 140.570 40.450 140.740 40.950 ;
        RECT 142.210 40.450 142.380 40.950 ;
        RECT 140.955 40.220 141.995 40.390 ;
        RECT 140.570 39.660 140.740 40.160 ;
        RECT 142.210 39.660 142.380 40.160 ;
        RECT 140.955 39.430 141.995 39.600 ;
        RECT 140.570 38.870 140.740 39.370 ;
        RECT 142.210 38.870 142.380 39.370 ;
        RECT 140.955 38.640 141.995 38.810 ;
        RECT 140.570 38.080 140.740 38.580 ;
        RECT 142.210 38.080 142.380 38.580 ;
        RECT 140.955 37.850 141.995 38.020 ;
        RECT 140.570 37.290 140.740 37.790 ;
        RECT 142.210 37.290 142.380 37.790 ;
        RECT 140.955 37.060 141.995 37.230 ;
        RECT 140.570 36.500 140.740 37.000 ;
        RECT 142.210 36.500 142.380 37.000 ;
        RECT 140.955 36.270 141.995 36.440 ;
        RECT 140.570 35.710 140.740 36.210 ;
        RECT 142.210 35.710 142.380 36.210 ;
        RECT 140.955 35.480 141.995 35.650 ;
        RECT 140.570 34.920 140.740 35.420 ;
        RECT 142.210 34.920 142.380 35.420 ;
        RECT 140.955 34.690 141.995 34.860 ;
        RECT 140.570 34.130 140.740 34.630 ;
        RECT 142.210 34.130 142.380 34.630 ;
        RECT 140.955 33.900 141.995 34.070 ;
        RECT 140.570 33.340 140.740 33.840 ;
        RECT 142.210 33.340 142.380 33.840 ;
        RECT 140.955 33.110 141.995 33.280 ;
        RECT 142.720 32.820 147.070 49.480 ;
        RECT 138.560 32.290 147.070 32.820 ;
        RECT 135.770 30.300 136.810 30.470 ;
        RECT 117.070 26.770 135.090 29.810 ;
        RECT 135.430 28.240 135.600 30.240 ;
        RECT 136.980 28.240 137.150 30.240 ;
        RECT 135.770 28.010 136.810 28.180 ;
        RECT 117.070 24.370 117.430 26.770 ;
        RECT 118.060 26.260 120.060 26.430 ;
        RECT 120.350 26.260 122.350 26.430 ;
        RECT 122.640 26.260 124.640 26.430 ;
        RECT 124.930 26.260 126.930 26.430 ;
        RECT 117.830 25.050 118.000 26.090 ;
        RECT 120.120 25.050 120.290 26.090 ;
        RECT 122.410 25.050 122.580 26.090 ;
        RECT 124.700 25.050 124.870 26.090 ;
        RECT 126.990 25.050 127.160 26.090 ;
        RECT 127.560 25.320 135.090 26.770 ;
        RECT 135.430 25.950 135.600 27.950 ;
        RECT 136.980 25.950 137.150 27.950 ;
        RECT 135.770 25.720 136.810 25.890 ;
        RECT 137.490 25.320 147.070 31.330 ;
        RECT 118.060 24.710 120.060 24.880 ;
        RECT 120.350 24.710 122.350 24.880 ;
        RECT 122.640 24.710 124.640 24.880 ;
        RECT 124.930 24.710 126.930 24.880 ;
        RECT 127.560 24.370 147.070 25.320 ;
        RECT 54.840 22.430 84.290 22.450 ;
        RECT 117.070 22.050 147.070 24.370 ;
        RECT 117.070 22.030 146.520 22.050 ;
      LAYER mcon ;
        RECT 11.265 213.545 11.435 213.715 ;
        RECT 11.725 213.545 11.895 213.715 ;
        RECT 12.185 213.545 12.355 213.715 ;
        RECT 12.645 213.545 12.815 213.715 ;
        RECT 13.105 213.545 13.275 213.715 ;
        RECT 13.565 213.545 13.735 213.715 ;
        RECT 14.025 213.545 14.195 213.715 ;
        RECT 14.485 213.545 14.655 213.715 ;
        RECT 14.945 213.545 15.115 213.715 ;
        RECT 15.405 213.545 15.575 213.715 ;
        RECT 15.865 213.545 16.035 213.715 ;
        RECT 16.325 213.545 16.495 213.715 ;
        RECT 16.785 213.545 16.955 213.715 ;
        RECT 17.245 213.545 17.415 213.715 ;
        RECT 17.705 213.545 17.875 213.715 ;
        RECT 18.165 213.545 18.335 213.715 ;
        RECT 18.625 213.545 18.795 213.715 ;
        RECT 19.085 213.545 19.255 213.715 ;
        RECT 19.545 213.545 19.715 213.715 ;
        RECT 20.005 213.545 20.175 213.715 ;
        RECT 20.465 213.545 20.635 213.715 ;
        RECT 20.925 213.545 21.095 213.715 ;
        RECT 21.385 213.545 21.555 213.715 ;
        RECT 21.845 213.545 22.015 213.715 ;
        RECT 22.305 213.545 22.475 213.715 ;
        RECT 22.765 213.545 22.935 213.715 ;
        RECT 23.225 213.545 23.395 213.715 ;
        RECT 23.685 213.545 23.855 213.715 ;
        RECT 24.145 213.545 24.315 213.715 ;
        RECT 24.605 213.545 24.775 213.715 ;
        RECT 25.065 213.545 25.235 213.715 ;
        RECT 25.525 213.545 25.695 213.715 ;
        RECT 25.985 213.545 26.155 213.715 ;
        RECT 26.445 213.545 26.615 213.715 ;
        RECT 26.905 213.545 27.075 213.715 ;
        RECT 27.365 213.545 27.535 213.715 ;
        RECT 27.825 213.545 27.995 213.715 ;
        RECT 28.285 213.545 28.455 213.715 ;
        RECT 28.745 213.545 28.915 213.715 ;
        RECT 29.205 213.545 29.375 213.715 ;
        RECT 29.665 213.545 29.835 213.715 ;
        RECT 30.125 213.545 30.295 213.715 ;
        RECT 30.585 213.545 30.755 213.715 ;
        RECT 31.045 213.545 31.215 213.715 ;
        RECT 31.505 213.545 31.675 213.715 ;
        RECT 31.965 213.545 32.135 213.715 ;
        RECT 32.425 213.545 32.595 213.715 ;
        RECT 32.885 213.545 33.055 213.715 ;
        RECT 33.345 213.545 33.515 213.715 ;
        RECT 33.805 213.545 33.975 213.715 ;
        RECT 34.265 213.545 34.435 213.715 ;
        RECT 34.725 213.545 34.895 213.715 ;
        RECT 35.185 213.545 35.355 213.715 ;
        RECT 35.645 213.545 35.815 213.715 ;
        RECT 36.105 213.545 36.275 213.715 ;
        RECT 36.565 213.545 36.735 213.715 ;
        RECT 37.025 213.545 37.195 213.715 ;
        RECT 37.485 213.545 37.655 213.715 ;
        RECT 37.945 213.545 38.115 213.715 ;
        RECT 38.405 213.545 38.575 213.715 ;
        RECT 38.865 213.545 39.035 213.715 ;
        RECT 39.325 213.545 39.495 213.715 ;
        RECT 39.785 213.545 39.955 213.715 ;
        RECT 40.245 213.545 40.415 213.715 ;
        RECT 40.705 213.545 40.875 213.715 ;
        RECT 41.165 213.545 41.335 213.715 ;
        RECT 41.625 213.545 41.795 213.715 ;
        RECT 42.085 213.545 42.255 213.715 ;
        RECT 42.545 213.545 42.715 213.715 ;
        RECT 43.005 213.545 43.175 213.715 ;
        RECT 43.465 213.545 43.635 213.715 ;
        RECT 43.925 213.545 44.095 213.715 ;
        RECT 44.385 213.545 44.555 213.715 ;
        RECT 44.845 213.545 45.015 213.715 ;
        RECT 45.305 213.545 45.475 213.715 ;
        RECT 45.765 213.545 45.935 213.715 ;
        RECT 46.225 213.545 46.395 213.715 ;
        RECT 46.685 213.545 46.855 213.715 ;
        RECT 47.145 213.545 47.315 213.715 ;
        RECT 47.605 213.545 47.775 213.715 ;
        RECT 48.065 213.545 48.235 213.715 ;
        RECT 48.525 213.545 48.695 213.715 ;
        RECT 48.985 213.545 49.155 213.715 ;
        RECT 49.445 213.545 49.615 213.715 ;
        RECT 49.905 213.545 50.075 213.715 ;
        RECT 50.365 213.545 50.535 213.715 ;
        RECT 50.825 213.545 50.995 213.715 ;
        RECT 51.285 213.545 51.455 213.715 ;
        RECT 51.745 213.545 51.915 213.715 ;
        RECT 52.205 213.545 52.375 213.715 ;
        RECT 52.665 213.545 52.835 213.715 ;
        RECT 53.125 213.545 53.295 213.715 ;
        RECT 53.585 213.545 53.755 213.715 ;
        RECT 54.045 213.545 54.215 213.715 ;
        RECT 54.505 213.545 54.675 213.715 ;
        RECT 54.965 213.545 55.135 213.715 ;
        RECT 55.425 213.545 55.595 213.715 ;
        RECT 55.885 213.545 56.055 213.715 ;
        RECT 56.345 213.545 56.515 213.715 ;
        RECT 56.805 213.545 56.975 213.715 ;
        RECT 57.265 213.545 57.435 213.715 ;
        RECT 57.725 213.545 57.895 213.715 ;
        RECT 58.185 213.545 58.355 213.715 ;
        RECT 58.645 213.545 58.815 213.715 ;
        RECT 59.105 213.545 59.275 213.715 ;
        RECT 59.565 213.545 59.735 213.715 ;
        RECT 60.025 213.545 60.195 213.715 ;
        RECT 60.485 213.545 60.655 213.715 ;
        RECT 60.945 213.545 61.115 213.715 ;
        RECT 61.405 213.545 61.575 213.715 ;
        RECT 61.865 213.545 62.035 213.715 ;
        RECT 62.325 213.545 62.495 213.715 ;
        RECT 62.785 213.545 62.955 213.715 ;
        RECT 63.245 213.545 63.415 213.715 ;
        RECT 63.705 213.545 63.875 213.715 ;
        RECT 64.165 213.545 64.335 213.715 ;
        RECT 64.625 213.545 64.795 213.715 ;
        RECT 65.085 213.545 65.255 213.715 ;
        RECT 65.545 213.545 65.715 213.715 ;
        RECT 66.005 213.545 66.175 213.715 ;
        RECT 66.465 213.545 66.635 213.715 ;
        RECT 66.925 213.545 67.095 213.715 ;
        RECT 67.385 213.545 67.555 213.715 ;
        RECT 67.845 213.545 68.015 213.715 ;
        RECT 68.305 213.545 68.475 213.715 ;
        RECT 68.765 213.545 68.935 213.715 ;
        RECT 69.225 213.545 69.395 213.715 ;
        RECT 69.685 213.545 69.855 213.715 ;
        RECT 70.145 213.545 70.315 213.715 ;
        RECT 70.605 213.545 70.775 213.715 ;
        RECT 71.065 213.545 71.235 213.715 ;
        RECT 71.525 213.545 71.695 213.715 ;
        RECT 71.985 213.545 72.155 213.715 ;
        RECT 72.445 213.545 72.615 213.715 ;
        RECT 72.905 213.545 73.075 213.715 ;
        RECT 73.365 213.545 73.535 213.715 ;
        RECT 73.825 213.545 73.995 213.715 ;
        RECT 74.285 213.545 74.455 213.715 ;
        RECT 74.745 213.545 74.915 213.715 ;
        RECT 75.205 213.545 75.375 213.715 ;
        RECT 75.665 213.545 75.835 213.715 ;
        RECT 76.125 213.545 76.295 213.715 ;
        RECT 76.585 213.545 76.755 213.715 ;
        RECT 77.045 213.545 77.215 213.715 ;
        RECT 77.505 213.545 77.675 213.715 ;
        RECT 77.965 213.545 78.135 213.715 ;
        RECT 78.425 213.545 78.595 213.715 ;
        RECT 78.885 213.545 79.055 213.715 ;
        RECT 79.345 213.545 79.515 213.715 ;
        RECT 79.805 213.545 79.975 213.715 ;
        RECT 80.265 213.545 80.435 213.715 ;
        RECT 80.725 213.545 80.895 213.715 ;
        RECT 81.185 213.545 81.355 213.715 ;
        RECT 81.645 213.545 81.815 213.715 ;
        RECT 82.105 213.545 82.275 213.715 ;
        RECT 82.565 213.545 82.735 213.715 ;
        RECT 83.025 213.545 83.195 213.715 ;
        RECT 83.485 213.545 83.655 213.715 ;
        RECT 83.945 213.545 84.115 213.715 ;
        RECT 84.405 213.545 84.575 213.715 ;
        RECT 84.865 213.545 85.035 213.715 ;
        RECT 85.325 213.545 85.495 213.715 ;
        RECT 85.785 213.545 85.955 213.715 ;
        RECT 86.245 213.545 86.415 213.715 ;
        RECT 86.705 213.545 86.875 213.715 ;
        RECT 87.165 213.545 87.335 213.715 ;
        RECT 87.625 213.545 87.795 213.715 ;
        RECT 88.085 213.545 88.255 213.715 ;
        RECT 88.545 213.545 88.715 213.715 ;
        RECT 89.005 213.545 89.175 213.715 ;
        RECT 89.465 213.545 89.635 213.715 ;
        RECT 89.925 213.545 90.095 213.715 ;
        RECT 90.385 213.545 90.555 213.715 ;
        RECT 90.845 213.545 91.015 213.715 ;
        RECT 91.305 213.545 91.475 213.715 ;
        RECT 91.765 213.545 91.935 213.715 ;
        RECT 92.225 213.545 92.395 213.715 ;
        RECT 92.685 213.545 92.855 213.715 ;
        RECT 93.145 213.545 93.315 213.715 ;
        RECT 93.605 213.545 93.775 213.715 ;
        RECT 94.065 213.545 94.235 213.715 ;
        RECT 94.525 213.545 94.695 213.715 ;
        RECT 94.985 213.545 95.155 213.715 ;
        RECT 95.445 213.545 95.615 213.715 ;
        RECT 95.905 213.545 96.075 213.715 ;
        RECT 96.365 213.545 96.535 213.715 ;
        RECT 96.825 213.545 96.995 213.715 ;
        RECT 97.285 213.545 97.455 213.715 ;
        RECT 97.745 213.545 97.915 213.715 ;
        RECT 98.205 213.545 98.375 213.715 ;
        RECT 98.665 213.545 98.835 213.715 ;
        RECT 99.125 213.545 99.295 213.715 ;
        RECT 99.585 213.545 99.755 213.715 ;
        RECT 100.045 213.545 100.215 213.715 ;
        RECT 100.505 213.545 100.675 213.715 ;
        RECT 100.965 213.545 101.135 213.715 ;
        RECT 101.425 213.545 101.595 213.715 ;
        RECT 101.885 213.545 102.055 213.715 ;
        RECT 102.345 213.545 102.515 213.715 ;
        RECT 102.805 213.545 102.975 213.715 ;
        RECT 103.265 213.545 103.435 213.715 ;
        RECT 103.725 213.545 103.895 213.715 ;
        RECT 104.185 213.545 104.355 213.715 ;
        RECT 104.645 213.545 104.815 213.715 ;
        RECT 105.105 213.545 105.275 213.715 ;
        RECT 105.565 213.545 105.735 213.715 ;
        RECT 106.025 213.545 106.195 213.715 ;
        RECT 106.485 213.545 106.655 213.715 ;
        RECT 106.945 213.545 107.115 213.715 ;
        RECT 107.405 213.545 107.575 213.715 ;
        RECT 107.865 213.545 108.035 213.715 ;
        RECT 108.325 213.545 108.495 213.715 ;
        RECT 108.785 213.545 108.955 213.715 ;
        RECT 109.245 213.545 109.415 213.715 ;
        RECT 109.705 213.545 109.875 213.715 ;
        RECT 110.165 213.545 110.335 213.715 ;
        RECT 110.625 213.545 110.795 213.715 ;
        RECT 111.085 213.545 111.255 213.715 ;
        RECT 111.545 213.545 111.715 213.715 ;
        RECT 112.005 213.545 112.175 213.715 ;
        RECT 112.465 213.545 112.635 213.715 ;
        RECT 112.925 213.545 113.095 213.715 ;
        RECT 113.385 213.545 113.555 213.715 ;
        RECT 113.845 213.545 114.015 213.715 ;
        RECT 114.305 213.545 114.475 213.715 ;
        RECT 114.765 213.545 114.935 213.715 ;
        RECT 115.225 213.545 115.395 213.715 ;
        RECT 115.685 213.545 115.855 213.715 ;
        RECT 116.145 213.545 116.315 213.715 ;
        RECT 116.605 213.545 116.775 213.715 ;
        RECT 117.065 213.545 117.235 213.715 ;
        RECT 117.525 213.545 117.695 213.715 ;
        RECT 117.985 213.545 118.155 213.715 ;
        RECT 118.445 213.545 118.615 213.715 ;
        RECT 118.905 213.545 119.075 213.715 ;
        RECT 119.365 213.545 119.535 213.715 ;
        RECT 119.825 213.545 119.995 213.715 ;
        RECT 120.285 213.545 120.455 213.715 ;
        RECT 120.745 213.545 120.915 213.715 ;
        RECT 121.205 213.545 121.375 213.715 ;
        RECT 121.665 213.545 121.835 213.715 ;
        RECT 122.125 213.545 122.295 213.715 ;
        RECT 122.585 213.545 122.755 213.715 ;
        RECT 123.045 213.545 123.215 213.715 ;
        RECT 123.505 213.545 123.675 213.715 ;
        RECT 123.965 213.545 124.135 213.715 ;
        RECT 124.425 213.545 124.595 213.715 ;
        RECT 124.885 213.545 125.055 213.715 ;
        RECT 125.345 213.545 125.515 213.715 ;
        RECT 125.805 213.545 125.975 213.715 ;
        RECT 126.265 213.545 126.435 213.715 ;
        RECT 126.725 213.545 126.895 213.715 ;
        RECT 127.185 213.545 127.355 213.715 ;
        RECT 127.645 213.545 127.815 213.715 ;
        RECT 128.105 213.545 128.275 213.715 ;
        RECT 128.565 213.545 128.735 213.715 ;
        RECT 129.025 213.545 129.195 213.715 ;
        RECT 129.485 213.545 129.655 213.715 ;
        RECT 129.945 213.545 130.115 213.715 ;
        RECT 130.405 213.545 130.575 213.715 ;
        RECT 130.865 213.545 131.035 213.715 ;
        RECT 131.325 213.545 131.495 213.715 ;
        RECT 131.785 213.545 131.955 213.715 ;
        RECT 132.245 213.545 132.415 213.715 ;
        RECT 132.705 213.545 132.875 213.715 ;
        RECT 133.165 213.545 133.335 213.715 ;
        RECT 133.625 213.545 133.795 213.715 ;
        RECT 134.085 213.545 134.255 213.715 ;
        RECT 134.545 213.545 134.715 213.715 ;
        RECT 135.005 213.545 135.175 213.715 ;
        RECT 135.465 213.545 135.635 213.715 ;
        RECT 135.925 213.545 136.095 213.715 ;
        RECT 136.385 213.545 136.555 213.715 ;
        RECT 136.845 213.545 137.015 213.715 ;
        RECT 137.305 213.545 137.475 213.715 ;
        RECT 137.765 213.545 137.935 213.715 ;
        RECT 138.225 213.545 138.395 213.715 ;
        RECT 138.685 213.545 138.855 213.715 ;
        RECT 139.145 213.545 139.315 213.715 ;
        RECT 139.605 213.545 139.775 213.715 ;
        RECT 140.065 213.545 140.235 213.715 ;
        RECT 140.525 213.545 140.695 213.715 ;
        RECT 140.985 213.545 141.155 213.715 ;
        RECT 141.445 213.545 141.615 213.715 ;
        RECT 141.905 213.545 142.075 213.715 ;
        RECT 142.365 213.545 142.535 213.715 ;
        RECT 142.825 213.545 142.995 213.715 ;
        RECT 143.285 213.545 143.455 213.715 ;
        RECT 143.745 213.545 143.915 213.715 ;
        RECT 144.205 213.545 144.375 213.715 ;
        RECT 144.665 213.545 144.835 213.715 ;
        RECT 145.125 213.545 145.295 213.715 ;
        RECT 145.585 213.545 145.755 213.715 ;
        RECT 146.045 213.545 146.215 213.715 ;
        RECT 146.505 213.545 146.675 213.715 ;
        RECT 146.965 213.545 147.135 213.715 ;
        RECT 147.425 213.545 147.595 213.715 ;
        RECT 147.885 213.545 148.055 213.715 ;
        RECT 148.345 213.545 148.515 213.715 ;
        RECT 148.805 213.545 148.975 213.715 ;
        RECT 149.265 213.545 149.435 213.715 ;
        RECT 149.725 213.545 149.895 213.715 ;
        RECT 150.185 213.545 150.355 213.715 ;
        RECT 65.085 213.035 65.255 213.205 ;
        RECT 64.165 212.015 64.335 212.185 ;
        RECT 86.705 212.015 86.875 212.185 ;
        RECT 87.625 211.335 87.795 211.505 ;
        RECT 96.365 212.015 96.535 212.185 ;
        RECT 97.285 211.335 97.455 211.505 ;
        RECT 104.645 212.015 104.815 212.185 ;
        RECT 107.865 211.335 108.035 211.505 ;
        RECT 109.245 212.015 109.415 212.185 ;
        RECT 108.785 211.335 108.955 211.505 ;
        RECT 110.625 212.015 110.795 212.185 ;
        RECT 109.705 211.335 109.875 211.505 ;
        RECT 117.525 212.015 117.695 212.185 ;
        RECT 116.605 211.335 116.775 211.505 ;
        RECT 128.565 212.015 128.735 212.185 ;
        RECT 127.645 211.335 127.815 211.505 ;
        RECT 137.305 212.015 137.475 212.185 ;
        RECT 137.765 211.335 137.935 211.505 ;
        RECT 11.265 210.825 11.435 210.995 ;
        RECT 11.725 210.825 11.895 210.995 ;
        RECT 12.185 210.825 12.355 210.995 ;
        RECT 12.645 210.825 12.815 210.995 ;
        RECT 13.105 210.825 13.275 210.995 ;
        RECT 13.565 210.825 13.735 210.995 ;
        RECT 14.025 210.825 14.195 210.995 ;
        RECT 14.485 210.825 14.655 210.995 ;
        RECT 14.945 210.825 15.115 210.995 ;
        RECT 15.405 210.825 15.575 210.995 ;
        RECT 15.865 210.825 16.035 210.995 ;
        RECT 16.325 210.825 16.495 210.995 ;
        RECT 16.785 210.825 16.955 210.995 ;
        RECT 17.245 210.825 17.415 210.995 ;
        RECT 17.705 210.825 17.875 210.995 ;
        RECT 18.165 210.825 18.335 210.995 ;
        RECT 18.625 210.825 18.795 210.995 ;
        RECT 19.085 210.825 19.255 210.995 ;
        RECT 19.545 210.825 19.715 210.995 ;
        RECT 20.005 210.825 20.175 210.995 ;
        RECT 20.465 210.825 20.635 210.995 ;
        RECT 20.925 210.825 21.095 210.995 ;
        RECT 21.385 210.825 21.555 210.995 ;
        RECT 21.845 210.825 22.015 210.995 ;
        RECT 22.305 210.825 22.475 210.995 ;
        RECT 22.765 210.825 22.935 210.995 ;
        RECT 23.225 210.825 23.395 210.995 ;
        RECT 23.685 210.825 23.855 210.995 ;
        RECT 24.145 210.825 24.315 210.995 ;
        RECT 24.605 210.825 24.775 210.995 ;
        RECT 25.065 210.825 25.235 210.995 ;
        RECT 25.525 210.825 25.695 210.995 ;
        RECT 25.985 210.825 26.155 210.995 ;
        RECT 26.445 210.825 26.615 210.995 ;
        RECT 26.905 210.825 27.075 210.995 ;
        RECT 27.365 210.825 27.535 210.995 ;
        RECT 27.825 210.825 27.995 210.995 ;
        RECT 28.285 210.825 28.455 210.995 ;
        RECT 28.745 210.825 28.915 210.995 ;
        RECT 29.205 210.825 29.375 210.995 ;
        RECT 29.665 210.825 29.835 210.995 ;
        RECT 30.125 210.825 30.295 210.995 ;
        RECT 30.585 210.825 30.755 210.995 ;
        RECT 31.045 210.825 31.215 210.995 ;
        RECT 31.505 210.825 31.675 210.995 ;
        RECT 31.965 210.825 32.135 210.995 ;
        RECT 32.425 210.825 32.595 210.995 ;
        RECT 32.885 210.825 33.055 210.995 ;
        RECT 33.345 210.825 33.515 210.995 ;
        RECT 33.805 210.825 33.975 210.995 ;
        RECT 34.265 210.825 34.435 210.995 ;
        RECT 34.725 210.825 34.895 210.995 ;
        RECT 35.185 210.825 35.355 210.995 ;
        RECT 35.645 210.825 35.815 210.995 ;
        RECT 36.105 210.825 36.275 210.995 ;
        RECT 36.565 210.825 36.735 210.995 ;
        RECT 37.025 210.825 37.195 210.995 ;
        RECT 37.485 210.825 37.655 210.995 ;
        RECT 37.945 210.825 38.115 210.995 ;
        RECT 38.405 210.825 38.575 210.995 ;
        RECT 38.865 210.825 39.035 210.995 ;
        RECT 39.325 210.825 39.495 210.995 ;
        RECT 39.785 210.825 39.955 210.995 ;
        RECT 40.245 210.825 40.415 210.995 ;
        RECT 40.705 210.825 40.875 210.995 ;
        RECT 41.165 210.825 41.335 210.995 ;
        RECT 41.625 210.825 41.795 210.995 ;
        RECT 42.085 210.825 42.255 210.995 ;
        RECT 42.545 210.825 42.715 210.995 ;
        RECT 43.005 210.825 43.175 210.995 ;
        RECT 43.465 210.825 43.635 210.995 ;
        RECT 43.925 210.825 44.095 210.995 ;
        RECT 44.385 210.825 44.555 210.995 ;
        RECT 44.845 210.825 45.015 210.995 ;
        RECT 45.305 210.825 45.475 210.995 ;
        RECT 45.765 210.825 45.935 210.995 ;
        RECT 46.225 210.825 46.395 210.995 ;
        RECT 46.685 210.825 46.855 210.995 ;
        RECT 47.145 210.825 47.315 210.995 ;
        RECT 47.605 210.825 47.775 210.995 ;
        RECT 48.065 210.825 48.235 210.995 ;
        RECT 48.525 210.825 48.695 210.995 ;
        RECT 48.985 210.825 49.155 210.995 ;
        RECT 49.445 210.825 49.615 210.995 ;
        RECT 49.905 210.825 50.075 210.995 ;
        RECT 50.365 210.825 50.535 210.995 ;
        RECT 50.825 210.825 50.995 210.995 ;
        RECT 51.285 210.825 51.455 210.995 ;
        RECT 51.745 210.825 51.915 210.995 ;
        RECT 52.205 210.825 52.375 210.995 ;
        RECT 52.665 210.825 52.835 210.995 ;
        RECT 53.125 210.825 53.295 210.995 ;
        RECT 53.585 210.825 53.755 210.995 ;
        RECT 54.045 210.825 54.215 210.995 ;
        RECT 54.505 210.825 54.675 210.995 ;
        RECT 54.965 210.825 55.135 210.995 ;
        RECT 55.425 210.825 55.595 210.995 ;
        RECT 55.885 210.825 56.055 210.995 ;
        RECT 56.345 210.825 56.515 210.995 ;
        RECT 56.805 210.825 56.975 210.995 ;
        RECT 57.265 210.825 57.435 210.995 ;
        RECT 57.725 210.825 57.895 210.995 ;
        RECT 58.185 210.825 58.355 210.995 ;
        RECT 58.645 210.825 58.815 210.995 ;
        RECT 59.105 210.825 59.275 210.995 ;
        RECT 59.565 210.825 59.735 210.995 ;
        RECT 60.025 210.825 60.195 210.995 ;
        RECT 60.485 210.825 60.655 210.995 ;
        RECT 60.945 210.825 61.115 210.995 ;
        RECT 61.405 210.825 61.575 210.995 ;
        RECT 61.865 210.825 62.035 210.995 ;
        RECT 62.325 210.825 62.495 210.995 ;
        RECT 62.785 210.825 62.955 210.995 ;
        RECT 63.245 210.825 63.415 210.995 ;
        RECT 63.705 210.825 63.875 210.995 ;
        RECT 64.165 210.825 64.335 210.995 ;
        RECT 64.625 210.825 64.795 210.995 ;
        RECT 65.085 210.825 65.255 210.995 ;
        RECT 65.545 210.825 65.715 210.995 ;
        RECT 66.005 210.825 66.175 210.995 ;
        RECT 66.465 210.825 66.635 210.995 ;
        RECT 66.925 210.825 67.095 210.995 ;
        RECT 67.385 210.825 67.555 210.995 ;
        RECT 67.845 210.825 68.015 210.995 ;
        RECT 68.305 210.825 68.475 210.995 ;
        RECT 68.765 210.825 68.935 210.995 ;
        RECT 69.225 210.825 69.395 210.995 ;
        RECT 69.685 210.825 69.855 210.995 ;
        RECT 70.145 210.825 70.315 210.995 ;
        RECT 70.605 210.825 70.775 210.995 ;
        RECT 71.065 210.825 71.235 210.995 ;
        RECT 71.525 210.825 71.695 210.995 ;
        RECT 71.985 210.825 72.155 210.995 ;
        RECT 72.445 210.825 72.615 210.995 ;
        RECT 72.905 210.825 73.075 210.995 ;
        RECT 73.365 210.825 73.535 210.995 ;
        RECT 73.825 210.825 73.995 210.995 ;
        RECT 74.285 210.825 74.455 210.995 ;
        RECT 74.745 210.825 74.915 210.995 ;
        RECT 75.205 210.825 75.375 210.995 ;
        RECT 75.665 210.825 75.835 210.995 ;
        RECT 76.125 210.825 76.295 210.995 ;
        RECT 76.585 210.825 76.755 210.995 ;
        RECT 77.045 210.825 77.215 210.995 ;
        RECT 77.505 210.825 77.675 210.995 ;
        RECT 77.965 210.825 78.135 210.995 ;
        RECT 78.425 210.825 78.595 210.995 ;
        RECT 78.885 210.825 79.055 210.995 ;
        RECT 79.345 210.825 79.515 210.995 ;
        RECT 79.805 210.825 79.975 210.995 ;
        RECT 80.265 210.825 80.435 210.995 ;
        RECT 80.725 210.825 80.895 210.995 ;
        RECT 81.185 210.825 81.355 210.995 ;
        RECT 81.645 210.825 81.815 210.995 ;
        RECT 82.105 210.825 82.275 210.995 ;
        RECT 82.565 210.825 82.735 210.995 ;
        RECT 83.025 210.825 83.195 210.995 ;
        RECT 83.485 210.825 83.655 210.995 ;
        RECT 83.945 210.825 84.115 210.995 ;
        RECT 84.405 210.825 84.575 210.995 ;
        RECT 84.865 210.825 85.035 210.995 ;
        RECT 85.325 210.825 85.495 210.995 ;
        RECT 85.785 210.825 85.955 210.995 ;
        RECT 86.245 210.825 86.415 210.995 ;
        RECT 86.705 210.825 86.875 210.995 ;
        RECT 87.165 210.825 87.335 210.995 ;
        RECT 87.625 210.825 87.795 210.995 ;
        RECT 88.085 210.825 88.255 210.995 ;
        RECT 88.545 210.825 88.715 210.995 ;
        RECT 89.005 210.825 89.175 210.995 ;
        RECT 89.465 210.825 89.635 210.995 ;
        RECT 89.925 210.825 90.095 210.995 ;
        RECT 90.385 210.825 90.555 210.995 ;
        RECT 90.845 210.825 91.015 210.995 ;
        RECT 91.305 210.825 91.475 210.995 ;
        RECT 91.765 210.825 91.935 210.995 ;
        RECT 92.225 210.825 92.395 210.995 ;
        RECT 92.685 210.825 92.855 210.995 ;
        RECT 93.145 210.825 93.315 210.995 ;
        RECT 93.605 210.825 93.775 210.995 ;
        RECT 94.065 210.825 94.235 210.995 ;
        RECT 94.525 210.825 94.695 210.995 ;
        RECT 94.985 210.825 95.155 210.995 ;
        RECT 95.445 210.825 95.615 210.995 ;
        RECT 95.905 210.825 96.075 210.995 ;
        RECT 96.365 210.825 96.535 210.995 ;
        RECT 96.825 210.825 96.995 210.995 ;
        RECT 97.285 210.825 97.455 210.995 ;
        RECT 97.745 210.825 97.915 210.995 ;
        RECT 98.205 210.825 98.375 210.995 ;
        RECT 98.665 210.825 98.835 210.995 ;
        RECT 99.125 210.825 99.295 210.995 ;
        RECT 99.585 210.825 99.755 210.995 ;
        RECT 100.045 210.825 100.215 210.995 ;
        RECT 100.505 210.825 100.675 210.995 ;
        RECT 100.965 210.825 101.135 210.995 ;
        RECT 101.425 210.825 101.595 210.995 ;
        RECT 101.885 210.825 102.055 210.995 ;
        RECT 102.345 210.825 102.515 210.995 ;
        RECT 102.805 210.825 102.975 210.995 ;
        RECT 103.265 210.825 103.435 210.995 ;
        RECT 103.725 210.825 103.895 210.995 ;
        RECT 104.185 210.825 104.355 210.995 ;
        RECT 104.645 210.825 104.815 210.995 ;
        RECT 105.105 210.825 105.275 210.995 ;
        RECT 105.565 210.825 105.735 210.995 ;
        RECT 106.025 210.825 106.195 210.995 ;
        RECT 106.485 210.825 106.655 210.995 ;
        RECT 106.945 210.825 107.115 210.995 ;
        RECT 107.405 210.825 107.575 210.995 ;
        RECT 107.865 210.825 108.035 210.995 ;
        RECT 108.325 210.825 108.495 210.995 ;
        RECT 108.785 210.825 108.955 210.995 ;
        RECT 109.245 210.825 109.415 210.995 ;
        RECT 109.705 210.825 109.875 210.995 ;
        RECT 110.165 210.825 110.335 210.995 ;
        RECT 110.625 210.825 110.795 210.995 ;
        RECT 111.085 210.825 111.255 210.995 ;
        RECT 111.545 210.825 111.715 210.995 ;
        RECT 112.005 210.825 112.175 210.995 ;
        RECT 112.465 210.825 112.635 210.995 ;
        RECT 112.925 210.825 113.095 210.995 ;
        RECT 113.385 210.825 113.555 210.995 ;
        RECT 113.845 210.825 114.015 210.995 ;
        RECT 114.305 210.825 114.475 210.995 ;
        RECT 114.765 210.825 114.935 210.995 ;
        RECT 115.225 210.825 115.395 210.995 ;
        RECT 115.685 210.825 115.855 210.995 ;
        RECT 116.145 210.825 116.315 210.995 ;
        RECT 116.605 210.825 116.775 210.995 ;
        RECT 117.065 210.825 117.235 210.995 ;
        RECT 117.525 210.825 117.695 210.995 ;
        RECT 117.985 210.825 118.155 210.995 ;
        RECT 118.445 210.825 118.615 210.995 ;
        RECT 118.905 210.825 119.075 210.995 ;
        RECT 119.365 210.825 119.535 210.995 ;
        RECT 119.825 210.825 119.995 210.995 ;
        RECT 120.285 210.825 120.455 210.995 ;
        RECT 120.745 210.825 120.915 210.995 ;
        RECT 121.205 210.825 121.375 210.995 ;
        RECT 121.665 210.825 121.835 210.995 ;
        RECT 122.125 210.825 122.295 210.995 ;
        RECT 122.585 210.825 122.755 210.995 ;
        RECT 123.045 210.825 123.215 210.995 ;
        RECT 123.505 210.825 123.675 210.995 ;
        RECT 123.965 210.825 124.135 210.995 ;
        RECT 124.425 210.825 124.595 210.995 ;
        RECT 124.885 210.825 125.055 210.995 ;
        RECT 125.345 210.825 125.515 210.995 ;
        RECT 125.805 210.825 125.975 210.995 ;
        RECT 126.265 210.825 126.435 210.995 ;
        RECT 126.725 210.825 126.895 210.995 ;
        RECT 127.185 210.825 127.355 210.995 ;
        RECT 127.645 210.825 127.815 210.995 ;
        RECT 128.105 210.825 128.275 210.995 ;
        RECT 128.565 210.825 128.735 210.995 ;
        RECT 129.025 210.825 129.195 210.995 ;
        RECT 129.485 210.825 129.655 210.995 ;
        RECT 129.945 210.825 130.115 210.995 ;
        RECT 130.405 210.825 130.575 210.995 ;
        RECT 130.865 210.825 131.035 210.995 ;
        RECT 131.325 210.825 131.495 210.995 ;
        RECT 131.785 210.825 131.955 210.995 ;
        RECT 132.245 210.825 132.415 210.995 ;
        RECT 132.705 210.825 132.875 210.995 ;
        RECT 133.165 210.825 133.335 210.995 ;
        RECT 133.625 210.825 133.795 210.995 ;
        RECT 134.085 210.825 134.255 210.995 ;
        RECT 134.545 210.825 134.715 210.995 ;
        RECT 135.005 210.825 135.175 210.995 ;
        RECT 135.465 210.825 135.635 210.995 ;
        RECT 135.925 210.825 136.095 210.995 ;
        RECT 136.385 210.825 136.555 210.995 ;
        RECT 136.845 210.825 137.015 210.995 ;
        RECT 137.305 210.825 137.475 210.995 ;
        RECT 137.765 210.825 137.935 210.995 ;
        RECT 138.225 210.825 138.395 210.995 ;
        RECT 138.685 210.825 138.855 210.995 ;
        RECT 139.145 210.825 139.315 210.995 ;
        RECT 139.605 210.825 139.775 210.995 ;
        RECT 140.065 210.825 140.235 210.995 ;
        RECT 140.525 210.825 140.695 210.995 ;
        RECT 140.985 210.825 141.155 210.995 ;
        RECT 141.445 210.825 141.615 210.995 ;
        RECT 141.905 210.825 142.075 210.995 ;
        RECT 142.365 210.825 142.535 210.995 ;
        RECT 142.825 210.825 142.995 210.995 ;
        RECT 143.285 210.825 143.455 210.995 ;
        RECT 143.745 210.825 143.915 210.995 ;
        RECT 144.205 210.825 144.375 210.995 ;
        RECT 144.665 210.825 144.835 210.995 ;
        RECT 145.125 210.825 145.295 210.995 ;
        RECT 145.585 210.825 145.755 210.995 ;
        RECT 146.045 210.825 146.215 210.995 ;
        RECT 146.505 210.825 146.675 210.995 ;
        RECT 146.965 210.825 147.135 210.995 ;
        RECT 147.425 210.825 147.595 210.995 ;
        RECT 147.885 210.825 148.055 210.995 ;
        RECT 148.345 210.825 148.515 210.995 ;
        RECT 148.805 210.825 148.975 210.995 ;
        RECT 149.265 210.825 149.435 210.995 ;
        RECT 149.725 210.825 149.895 210.995 ;
        RECT 150.185 210.825 150.355 210.995 ;
        RECT 15.405 209.975 15.575 210.145 ;
        RECT 17.245 209.635 17.415 209.805 ;
        RECT 20.005 209.295 20.175 209.465 ;
        RECT 20.490 208.955 20.660 209.125 ;
        RECT 20.885 209.295 21.055 209.465 ;
        RECT 21.340 209.635 21.510 209.805 ;
        RECT 22.075 209.295 22.245 209.465 ;
        RECT 22.590 208.955 22.760 209.125 ;
        RECT 24.160 208.955 24.330 209.125 ;
        RECT 24.595 209.295 24.765 209.465 ;
        RECT 27.365 209.975 27.535 210.145 ;
        RECT 26.905 208.615 27.075 208.785 ;
        RECT 29.205 209.635 29.375 209.805 ;
        RECT 31.505 209.975 31.675 210.145 ;
        RECT 32.425 209.635 32.595 209.805 ;
        RECT 32.885 209.635 33.055 209.805 ;
        RECT 34.265 209.975 34.435 210.145 ;
        RECT 33.805 209.635 33.975 209.805 ;
        RECT 30.585 208.615 30.755 208.785 ;
        RECT 33.345 208.615 33.515 208.785 ;
        RECT 36.105 209.635 36.275 209.805 ;
        RECT 38.405 209.635 38.575 209.805 ;
        RECT 37.485 208.615 37.655 208.785 ;
        RECT 42.085 210.315 42.255 210.485 ;
        RECT 40.245 209.635 40.415 209.805 ;
        RECT 39.785 209.295 39.955 209.465 ;
        RECT 44.385 209.635 44.555 209.805 ;
        RECT 43.465 208.955 43.635 209.125 ;
        RECT 46.225 209.635 46.395 209.805 ;
        RECT 46.685 209.295 46.855 209.465 ;
        RECT 48.065 208.955 48.235 209.125 ;
        RECT 49.445 209.635 49.615 209.805 ;
        RECT 48.985 209.295 49.155 209.465 ;
        RECT 51.285 209.295 51.455 209.465 ;
        RECT 53.125 209.635 53.295 209.805 ;
        RECT 52.665 209.295 52.835 209.465 ;
        RECT 55.425 209.635 55.595 209.805 ;
        RECT 55.910 208.955 56.080 209.125 ;
        RECT 56.305 209.295 56.475 209.465 ;
        RECT 54.505 208.615 54.675 208.785 ;
        RECT 56.760 209.635 56.930 209.805 ;
        RECT 57.495 209.295 57.665 209.465 ;
        RECT 58.010 208.955 58.180 209.125 ;
        RECT 59.580 208.955 59.750 209.125 ;
        RECT 60.015 209.295 60.185 209.465 ;
        RECT 64.165 209.635 64.335 209.805 ;
        RECT 62.325 208.615 62.495 208.785 ;
        RECT 64.650 208.955 64.820 209.125 ;
        RECT 65.045 209.295 65.215 209.465 ;
        RECT 65.445 209.635 65.615 209.805 ;
        RECT 66.235 209.295 66.405 209.465 ;
        RECT 66.750 208.955 66.920 209.125 ;
        RECT 68.320 208.955 68.490 209.125 ;
        RECT 68.755 209.295 68.925 209.465 ;
        RECT 71.985 209.635 72.155 209.805 ;
        RECT 71.065 208.955 71.235 209.125 ;
        RECT 74.285 209.635 74.455 209.805 ;
        RECT 73.365 208.615 73.535 208.785 ;
        RECT 74.770 208.955 74.940 209.125 ;
        RECT 75.165 209.295 75.335 209.465 ;
        RECT 75.565 209.635 75.735 209.805 ;
        RECT 76.355 209.295 76.525 209.465 ;
        RECT 76.870 208.955 77.040 209.125 ;
        RECT 78.440 208.955 78.610 209.125 ;
        RECT 78.875 209.295 79.045 209.465 ;
        RECT 81.185 210.315 81.355 210.485 ;
        RECT 81.645 208.955 81.815 209.125 ;
        RECT 84.405 210.315 84.575 210.485 ;
        RECT 83.485 209.975 83.655 210.145 ;
        RECT 83.485 208.615 83.655 208.785 ;
        RECT 85.325 209.975 85.495 210.145 ;
        RECT 87.165 209.975 87.335 210.145 ;
        RECT 89.005 209.295 89.175 209.465 ;
        RECT 89.490 208.955 89.660 209.125 ;
        RECT 89.885 209.295 90.055 209.465 ;
        RECT 90.285 209.635 90.455 209.805 ;
        RECT 91.075 209.295 91.245 209.465 ;
        RECT 91.590 208.955 91.760 209.125 ;
        RECT 93.160 208.955 93.330 209.125 ;
        RECT 93.595 209.295 93.765 209.465 ;
        RECT 96.825 209.635 96.995 209.805 ;
        RECT 95.905 208.615 96.075 208.785 ;
        RECT 97.310 208.955 97.480 209.125 ;
        RECT 97.705 209.295 97.875 209.465 ;
        RECT 98.160 209.635 98.330 209.805 ;
        RECT 98.895 209.295 99.065 209.465 ;
        RECT 99.410 208.955 99.580 209.125 ;
        RECT 100.980 208.955 101.150 209.125 ;
        RECT 101.415 209.295 101.585 209.465 ;
        RECT 103.725 210.315 103.895 210.485 ;
        RECT 104.185 209.295 104.355 209.465 ;
        RECT 104.670 208.955 104.840 209.125 ;
        RECT 105.065 209.295 105.235 209.465 ;
        RECT 105.520 209.975 105.690 210.145 ;
        RECT 106.255 209.295 106.425 209.465 ;
        RECT 106.770 208.955 106.940 209.125 ;
        RECT 108.340 208.955 108.510 209.125 ;
        RECT 108.775 209.295 108.945 209.465 ;
        RECT 111.545 209.635 111.715 209.805 ;
        RECT 111.085 208.955 111.255 209.125 ;
        RECT 113.845 209.635 114.015 209.805 ;
        RECT 112.005 208.615 112.175 208.785 ;
        RECT 113.385 208.615 113.555 208.785 ;
        RECT 116.145 208.955 116.315 209.125 ;
        RECT 118.455 209.295 118.625 209.465 ;
        RECT 118.890 208.955 119.060 209.125 ;
        RECT 120.975 209.295 121.145 209.465 ;
        RECT 120.460 208.955 120.630 209.125 ;
        RECT 121.765 209.635 121.935 209.805 ;
        RECT 122.165 209.295 122.335 209.465 ;
        RECT 123.045 209.295 123.215 209.465 ;
        RECT 123.505 209.295 123.675 209.465 ;
        RECT 122.560 208.955 122.730 209.125 ;
        RECT 123.990 208.955 124.160 209.125 ;
        RECT 124.385 209.295 124.555 209.465 ;
        RECT 124.840 209.635 125.010 209.805 ;
        RECT 125.575 209.295 125.745 209.465 ;
        RECT 126.090 208.955 126.260 209.125 ;
        RECT 127.660 208.955 127.830 209.125 ;
        RECT 128.095 209.295 128.265 209.465 ;
        RECT 130.405 208.615 130.575 208.785 ;
        RECT 11.265 208.105 11.435 208.275 ;
        RECT 11.725 208.105 11.895 208.275 ;
        RECT 12.185 208.105 12.355 208.275 ;
        RECT 12.645 208.105 12.815 208.275 ;
        RECT 13.105 208.105 13.275 208.275 ;
        RECT 13.565 208.105 13.735 208.275 ;
        RECT 14.025 208.105 14.195 208.275 ;
        RECT 14.485 208.105 14.655 208.275 ;
        RECT 14.945 208.105 15.115 208.275 ;
        RECT 15.405 208.105 15.575 208.275 ;
        RECT 15.865 208.105 16.035 208.275 ;
        RECT 16.325 208.105 16.495 208.275 ;
        RECT 16.785 208.105 16.955 208.275 ;
        RECT 17.245 208.105 17.415 208.275 ;
        RECT 17.705 208.105 17.875 208.275 ;
        RECT 18.165 208.105 18.335 208.275 ;
        RECT 18.625 208.105 18.795 208.275 ;
        RECT 19.085 208.105 19.255 208.275 ;
        RECT 19.545 208.105 19.715 208.275 ;
        RECT 20.005 208.105 20.175 208.275 ;
        RECT 20.465 208.105 20.635 208.275 ;
        RECT 20.925 208.105 21.095 208.275 ;
        RECT 21.385 208.105 21.555 208.275 ;
        RECT 21.845 208.105 22.015 208.275 ;
        RECT 22.305 208.105 22.475 208.275 ;
        RECT 22.765 208.105 22.935 208.275 ;
        RECT 23.225 208.105 23.395 208.275 ;
        RECT 23.685 208.105 23.855 208.275 ;
        RECT 24.145 208.105 24.315 208.275 ;
        RECT 24.605 208.105 24.775 208.275 ;
        RECT 25.065 208.105 25.235 208.275 ;
        RECT 25.525 208.105 25.695 208.275 ;
        RECT 25.985 208.105 26.155 208.275 ;
        RECT 26.445 208.105 26.615 208.275 ;
        RECT 26.905 208.105 27.075 208.275 ;
        RECT 27.365 208.105 27.535 208.275 ;
        RECT 27.825 208.105 27.995 208.275 ;
        RECT 28.285 208.105 28.455 208.275 ;
        RECT 28.745 208.105 28.915 208.275 ;
        RECT 29.205 208.105 29.375 208.275 ;
        RECT 29.665 208.105 29.835 208.275 ;
        RECT 30.125 208.105 30.295 208.275 ;
        RECT 30.585 208.105 30.755 208.275 ;
        RECT 31.045 208.105 31.215 208.275 ;
        RECT 31.505 208.105 31.675 208.275 ;
        RECT 31.965 208.105 32.135 208.275 ;
        RECT 32.425 208.105 32.595 208.275 ;
        RECT 32.885 208.105 33.055 208.275 ;
        RECT 33.345 208.105 33.515 208.275 ;
        RECT 33.805 208.105 33.975 208.275 ;
        RECT 34.265 208.105 34.435 208.275 ;
        RECT 34.725 208.105 34.895 208.275 ;
        RECT 35.185 208.105 35.355 208.275 ;
        RECT 35.645 208.105 35.815 208.275 ;
        RECT 36.105 208.105 36.275 208.275 ;
        RECT 36.565 208.105 36.735 208.275 ;
        RECT 37.025 208.105 37.195 208.275 ;
        RECT 37.485 208.105 37.655 208.275 ;
        RECT 37.945 208.105 38.115 208.275 ;
        RECT 38.405 208.105 38.575 208.275 ;
        RECT 38.865 208.105 39.035 208.275 ;
        RECT 39.325 208.105 39.495 208.275 ;
        RECT 39.785 208.105 39.955 208.275 ;
        RECT 40.245 208.105 40.415 208.275 ;
        RECT 40.705 208.105 40.875 208.275 ;
        RECT 41.165 208.105 41.335 208.275 ;
        RECT 41.625 208.105 41.795 208.275 ;
        RECT 42.085 208.105 42.255 208.275 ;
        RECT 42.545 208.105 42.715 208.275 ;
        RECT 43.005 208.105 43.175 208.275 ;
        RECT 43.465 208.105 43.635 208.275 ;
        RECT 43.925 208.105 44.095 208.275 ;
        RECT 44.385 208.105 44.555 208.275 ;
        RECT 44.845 208.105 45.015 208.275 ;
        RECT 45.305 208.105 45.475 208.275 ;
        RECT 45.765 208.105 45.935 208.275 ;
        RECT 46.225 208.105 46.395 208.275 ;
        RECT 46.685 208.105 46.855 208.275 ;
        RECT 47.145 208.105 47.315 208.275 ;
        RECT 47.605 208.105 47.775 208.275 ;
        RECT 48.065 208.105 48.235 208.275 ;
        RECT 48.525 208.105 48.695 208.275 ;
        RECT 48.985 208.105 49.155 208.275 ;
        RECT 49.445 208.105 49.615 208.275 ;
        RECT 49.905 208.105 50.075 208.275 ;
        RECT 50.365 208.105 50.535 208.275 ;
        RECT 50.825 208.105 50.995 208.275 ;
        RECT 51.285 208.105 51.455 208.275 ;
        RECT 51.745 208.105 51.915 208.275 ;
        RECT 52.205 208.105 52.375 208.275 ;
        RECT 52.665 208.105 52.835 208.275 ;
        RECT 53.125 208.105 53.295 208.275 ;
        RECT 53.585 208.105 53.755 208.275 ;
        RECT 54.045 208.105 54.215 208.275 ;
        RECT 54.505 208.105 54.675 208.275 ;
        RECT 54.965 208.105 55.135 208.275 ;
        RECT 55.425 208.105 55.595 208.275 ;
        RECT 55.885 208.105 56.055 208.275 ;
        RECT 56.345 208.105 56.515 208.275 ;
        RECT 56.805 208.105 56.975 208.275 ;
        RECT 57.265 208.105 57.435 208.275 ;
        RECT 57.725 208.105 57.895 208.275 ;
        RECT 58.185 208.105 58.355 208.275 ;
        RECT 58.645 208.105 58.815 208.275 ;
        RECT 59.105 208.105 59.275 208.275 ;
        RECT 59.565 208.105 59.735 208.275 ;
        RECT 60.025 208.105 60.195 208.275 ;
        RECT 60.485 208.105 60.655 208.275 ;
        RECT 60.945 208.105 61.115 208.275 ;
        RECT 61.405 208.105 61.575 208.275 ;
        RECT 61.865 208.105 62.035 208.275 ;
        RECT 62.325 208.105 62.495 208.275 ;
        RECT 62.785 208.105 62.955 208.275 ;
        RECT 63.245 208.105 63.415 208.275 ;
        RECT 63.705 208.105 63.875 208.275 ;
        RECT 64.165 208.105 64.335 208.275 ;
        RECT 64.625 208.105 64.795 208.275 ;
        RECT 65.085 208.105 65.255 208.275 ;
        RECT 65.545 208.105 65.715 208.275 ;
        RECT 66.005 208.105 66.175 208.275 ;
        RECT 66.465 208.105 66.635 208.275 ;
        RECT 66.925 208.105 67.095 208.275 ;
        RECT 67.385 208.105 67.555 208.275 ;
        RECT 67.845 208.105 68.015 208.275 ;
        RECT 68.305 208.105 68.475 208.275 ;
        RECT 68.765 208.105 68.935 208.275 ;
        RECT 69.225 208.105 69.395 208.275 ;
        RECT 69.685 208.105 69.855 208.275 ;
        RECT 70.145 208.105 70.315 208.275 ;
        RECT 70.605 208.105 70.775 208.275 ;
        RECT 71.065 208.105 71.235 208.275 ;
        RECT 71.525 208.105 71.695 208.275 ;
        RECT 71.985 208.105 72.155 208.275 ;
        RECT 72.445 208.105 72.615 208.275 ;
        RECT 72.905 208.105 73.075 208.275 ;
        RECT 73.365 208.105 73.535 208.275 ;
        RECT 73.825 208.105 73.995 208.275 ;
        RECT 74.285 208.105 74.455 208.275 ;
        RECT 74.745 208.105 74.915 208.275 ;
        RECT 75.205 208.105 75.375 208.275 ;
        RECT 75.665 208.105 75.835 208.275 ;
        RECT 76.125 208.105 76.295 208.275 ;
        RECT 76.585 208.105 76.755 208.275 ;
        RECT 77.045 208.105 77.215 208.275 ;
        RECT 77.505 208.105 77.675 208.275 ;
        RECT 77.965 208.105 78.135 208.275 ;
        RECT 78.425 208.105 78.595 208.275 ;
        RECT 78.885 208.105 79.055 208.275 ;
        RECT 79.345 208.105 79.515 208.275 ;
        RECT 79.805 208.105 79.975 208.275 ;
        RECT 80.265 208.105 80.435 208.275 ;
        RECT 80.725 208.105 80.895 208.275 ;
        RECT 81.185 208.105 81.355 208.275 ;
        RECT 81.645 208.105 81.815 208.275 ;
        RECT 82.105 208.105 82.275 208.275 ;
        RECT 82.565 208.105 82.735 208.275 ;
        RECT 83.025 208.105 83.195 208.275 ;
        RECT 83.485 208.105 83.655 208.275 ;
        RECT 83.945 208.105 84.115 208.275 ;
        RECT 84.405 208.105 84.575 208.275 ;
        RECT 84.865 208.105 85.035 208.275 ;
        RECT 85.325 208.105 85.495 208.275 ;
        RECT 85.785 208.105 85.955 208.275 ;
        RECT 86.245 208.105 86.415 208.275 ;
        RECT 86.705 208.105 86.875 208.275 ;
        RECT 87.165 208.105 87.335 208.275 ;
        RECT 87.625 208.105 87.795 208.275 ;
        RECT 88.085 208.105 88.255 208.275 ;
        RECT 88.545 208.105 88.715 208.275 ;
        RECT 89.005 208.105 89.175 208.275 ;
        RECT 89.465 208.105 89.635 208.275 ;
        RECT 89.925 208.105 90.095 208.275 ;
        RECT 90.385 208.105 90.555 208.275 ;
        RECT 90.845 208.105 91.015 208.275 ;
        RECT 91.305 208.105 91.475 208.275 ;
        RECT 91.765 208.105 91.935 208.275 ;
        RECT 92.225 208.105 92.395 208.275 ;
        RECT 92.685 208.105 92.855 208.275 ;
        RECT 93.145 208.105 93.315 208.275 ;
        RECT 93.605 208.105 93.775 208.275 ;
        RECT 94.065 208.105 94.235 208.275 ;
        RECT 94.525 208.105 94.695 208.275 ;
        RECT 94.985 208.105 95.155 208.275 ;
        RECT 95.445 208.105 95.615 208.275 ;
        RECT 95.905 208.105 96.075 208.275 ;
        RECT 96.365 208.105 96.535 208.275 ;
        RECT 96.825 208.105 96.995 208.275 ;
        RECT 97.285 208.105 97.455 208.275 ;
        RECT 97.745 208.105 97.915 208.275 ;
        RECT 98.205 208.105 98.375 208.275 ;
        RECT 98.665 208.105 98.835 208.275 ;
        RECT 99.125 208.105 99.295 208.275 ;
        RECT 99.585 208.105 99.755 208.275 ;
        RECT 100.045 208.105 100.215 208.275 ;
        RECT 100.505 208.105 100.675 208.275 ;
        RECT 100.965 208.105 101.135 208.275 ;
        RECT 101.425 208.105 101.595 208.275 ;
        RECT 101.885 208.105 102.055 208.275 ;
        RECT 102.345 208.105 102.515 208.275 ;
        RECT 102.805 208.105 102.975 208.275 ;
        RECT 103.265 208.105 103.435 208.275 ;
        RECT 103.725 208.105 103.895 208.275 ;
        RECT 104.185 208.105 104.355 208.275 ;
        RECT 104.645 208.105 104.815 208.275 ;
        RECT 105.105 208.105 105.275 208.275 ;
        RECT 105.565 208.105 105.735 208.275 ;
        RECT 106.025 208.105 106.195 208.275 ;
        RECT 106.485 208.105 106.655 208.275 ;
        RECT 106.945 208.105 107.115 208.275 ;
        RECT 107.405 208.105 107.575 208.275 ;
        RECT 107.865 208.105 108.035 208.275 ;
        RECT 108.325 208.105 108.495 208.275 ;
        RECT 108.785 208.105 108.955 208.275 ;
        RECT 109.245 208.105 109.415 208.275 ;
        RECT 109.705 208.105 109.875 208.275 ;
        RECT 110.165 208.105 110.335 208.275 ;
        RECT 110.625 208.105 110.795 208.275 ;
        RECT 111.085 208.105 111.255 208.275 ;
        RECT 111.545 208.105 111.715 208.275 ;
        RECT 112.005 208.105 112.175 208.275 ;
        RECT 112.465 208.105 112.635 208.275 ;
        RECT 112.925 208.105 113.095 208.275 ;
        RECT 113.385 208.105 113.555 208.275 ;
        RECT 113.845 208.105 114.015 208.275 ;
        RECT 114.305 208.105 114.475 208.275 ;
        RECT 114.765 208.105 114.935 208.275 ;
        RECT 115.225 208.105 115.395 208.275 ;
        RECT 115.685 208.105 115.855 208.275 ;
        RECT 116.145 208.105 116.315 208.275 ;
        RECT 116.605 208.105 116.775 208.275 ;
        RECT 117.065 208.105 117.235 208.275 ;
        RECT 117.525 208.105 117.695 208.275 ;
        RECT 117.985 208.105 118.155 208.275 ;
        RECT 118.445 208.105 118.615 208.275 ;
        RECT 118.905 208.105 119.075 208.275 ;
        RECT 119.365 208.105 119.535 208.275 ;
        RECT 119.825 208.105 119.995 208.275 ;
        RECT 120.285 208.105 120.455 208.275 ;
        RECT 120.745 208.105 120.915 208.275 ;
        RECT 121.205 208.105 121.375 208.275 ;
        RECT 121.665 208.105 121.835 208.275 ;
        RECT 122.125 208.105 122.295 208.275 ;
        RECT 122.585 208.105 122.755 208.275 ;
        RECT 123.045 208.105 123.215 208.275 ;
        RECT 123.505 208.105 123.675 208.275 ;
        RECT 123.965 208.105 124.135 208.275 ;
        RECT 124.425 208.105 124.595 208.275 ;
        RECT 124.885 208.105 125.055 208.275 ;
        RECT 125.345 208.105 125.515 208.275 ;
        RECT 125.805 208.105 125.975 208.275 ;
        RECT 126.265 208.105 126.435 208.275 ;
        RECT 126.725 208.105 126.895 208.275 ;
        RECT 127.185 208.105 127.355 208.275 ;
        RECT 127.645 208.105 127.815 208.275 ;
        RECT 128.105 208.105 128.275 208.275 ;
        RECT 128.565 208.105 128.735 208.275 ;
        RECT 129.025 208.105 129.195 208.275 ;
        RECT 129.485 208.105 129.655 208.275 ;
        RECT 129.945 208.105 130.115 208.275 ;
        RECT 130.405 208.105 130.575 208.275 ;
        RECT 130.865 208.105 131.035 208.275 ;
        RECT 131.325 208.105 131.495 208.275 ;
        RECT 131.785 208.105 131.955 208.275 ;
        RECT 132.245 208.105 132.415 208.275 ;
        RECT 132.705 208.105 132.875 208.275 ;
        RECT 133.165 208.105 133.335 208.275 ;
        RECT 133.625 208.105 133.795 208.275 ;
        RECT 134.085 208.105 134.255 208.275 ;
        RECT 134.545 208.105 134.715 208.275 ;
        RECT 135.005 208.105 135.175 208.275 ;
        RECT 135.465 208.105 135.635 208.275 ;
        RECT 135.925 208.105 136.095 208.275 ;
        RECT 136.385 208.105 136.555 208.275 ;
        RECT 136.845 208.105 137.015 208.275 ;
        RECT 137.305 208.105 137.475 208.275 ;
        RECT 137.765 208.105 137.935 208.275 ;
        RECT 138.225 208.105 138.395 208.275 ;
        RECT 138.685 208.105 138.855 208.275 ;
        RECT 139.145 208.105 139.315 208.275 ;
        RECT 139.605 208.105 139.775 208.275 ;
        RECT 140.065 208.105 140.235 208.275 ;
        RECT 140.525 208.105 140.695 208.275 ;
        RECT 140.985 208.105 141.155 208.275 ;
        RECT 141.445 208.105 141.615 208.275 ;
        RECT 141.905 208.105 142.075 208.275 ;
        RECT 142.365 208.105 142.535 208.275 ;
        RECT 142.825 208.105 142.995 208.275 ;
        RECT 143.285 208.105 143.455 208.275 ;
        RECT 143.745 208.105 143.915 208.275 ;
        RECT 144.205 208.105 144.375 208.275 ;
        RECT 144.665 208.105 144.835 208.275 ;
        RECT 145.125 208.105 145.295 208.275 ;
        RECT 145.585 208.105 145.755 208.275 ;
        RECT 146.045 208.105 146.215 208.275 ;
        RECT 146.505 208.105 146.675 208.275 ;
        RECT 146.965 208.105 147.135 208.275 ;
        RECT 147.425 208.105 147.595 208.275 ;
        RECT 147.885 208.105 148.055 208.275 ;
        RECT 148.345 208.105 148.515 208.275 ;
        RECT 148.805 208.105 148.975 208.275 ;
        RECT 149.265 208.105 149.435 208.275 ;
        RECT 149.725 208.105 149.895 208.275 ;
        RECT 150.185 208.105 150.355 208.275 ;
        RECT 22.305 207.595 22.475 207.765 ;
        RECT 25.525 207.595 25.695 207.765 ;
        RECT 24.605 207.255 24.775 207.425 ;
        RECT 23.225 206.575 23.395 206.745 ;
        RECT 25.525 205.895 25.695 206.065 ;
        RECT 27.365 206.575 27.535 206.745 ;
        RECT 32.885 207.255 33.055 207.425 ;
        RECT 28.745 206.575 28.915 206.745 ;
        RECT 27.825 205.895 27.995 206.065 ;
        RECT 30.125 206.575 30.295 206.745 ;
        RECT 29.665 205.895 29.835 206.065 ;
        RECT 35.195 206.915 35.365 207.085 ;
        RECT 35.630 207.255 35.800 207.425 ;
        RECT 37.200 207.255 37.370 207.425 ;
        RECT 37.715 206.915 37.885 207.085 ;
        RECT 38.450 206.575 38.620 206.745 ;
        RECT 38.905 206.915 39.075 207.085 ;
        RECT 39.300 207.255 39.470 207.425 ;
        RECT 39.785 206.575 39.955 206.745 ;
        RECT 47.605 207.595 47.775 207.765 ;
        RECT 47.145 207.255 47.315 207.425 ;
        RECT 53.125 207.595 53.295 207.765 ;
        RECT 52.205 206.575 52.375 206.745 ;
        RECT 65.085 207.595 65.255 207.765 ;
        RECT 64.625 206.575 64.795 206.745 ;
        RECT 67.385 207.255 67.555 207.425 ;
        RECT 70.145 206.915 70.315 207.085 ;
        RECT 73.825 207.595 73.995 207.765 ;
        RECT 68.305 205.895 68.475 206.065 ;
        RECT 68.765 205.895 68.935 206.065 ;
        RECT 69.225 206.235 69.395 206.405 ;
        RECT 70.605 206.575 70.775 206.745 ;
        RECT 71.525 206.575 71.695 206.745 ;
        RECT 71.985 206.575 72.155 206.745 ;
        RECT 72.445 206.575 72.615 206.745 ;
        RECT 83.485 207.595 83.655 207.765 ;
        RECT 81.645 206.575 81.815 206.745 ;
        RECT 82.565 206.235 82.735 206.405 ;
        RECT 85.810 207.255 85.980 207.425 ;
        RECT 83.945 206.575 84.115 206.745 ;
        RECT 85.325 206.915 85.495 207.085 ;
        RECT 84.865 206.575 85.035 206.745 ;
        RECT 84.405 206.235 84.575 206.405 ;
        RECT 86.205 206.915 86.375 207.085 ;
        RECT 86.550 206.235 86.720 206.405 ;
        RECT 87.910 207.255 88.080 207.425 ;
        RECT 87.395 206.915 87.565 207.085 ;
        RECT 89.480 207.255 89.650 207.425 ;
        RECT 89.915 206.915 90.085 207.085 ;
        RECT 92.225 207.255 92.395 207.425 ;
        RECT 93.145 205.895 93.315 206.065 ;
        RECT 95.905 206.915 96.075 207.085 ;
        RECT 97.745 206.575 97.915 206.745 ;
        RECT 100.045 207.595 100.215 207.765 ;
        RECT 99.585 206.575 99.755 206.745 ;
        RECT 98.665 205.895 98.835 206.065 ;
        RECT 104.210 207.255 104.380 207.425 ;
        RECT 103.725 206.575 103.895 206.745 ;
        RECT 104.605 206.915 104.775 207.085 ;
        RECT 105.060 206.235 105.230 206.405 ;
        RECT 106.310 207.255 106.480 207.425 ;
        RECT 105.795 206.915 105.965 207.085 ;
        RECT 107.880 207.255 108.050 207.425 ;
        RECT 108.315 206.915 108.485 207.085 ;
        RECT 112.030 207.255 112.200 207.425 ;
        RECT 111.545 206.575 111.715 206.745 ;
        RECT 110.625 205.895 110.795 206.065 ;
        RECT 112.425 206.915 112.595 207.085 ;
        RECT 112.880 206.575 113.050 206.745 ;
        RECT 114.130 207.255 114.300 207.425 ;
        RECT 113.615 206.915 113.785 207.085 ;
        RECT 115.700 207.255 115.870 207.425 ;
        RECT 116.135 206.915 116.305 207.085 ;
        RECT 118.445 207.255 118.615 207.425 ;
        RECT 120.285 206.915 120.455 207.085 ;
        RECT 123.505 207.595 123.675 207.765 ;
        RECT 124.425 207.595 124.595 207.765 ;
        RECT 124.885 206.575 125.055 206.745 ;
        RECT 129.945 205.895 130.115 206.065 ;
        RECT 132.705 206.915 132.875 207.085 ;
        RECT 11.265 205.385 11.435 205.555 ;
        RECT 11.725 205.385 11.895 205.555 ;
        RECT 12.185 205.385 12.355 205.555 ;
        RECT 12.645 205.385 12.815 205.555 ;
        RECT 13.105 205.385 13.275 205.555 ;
        RECT 13.565 205.385 13.735 205.555 ;
        RECT 14.025 205.385 14.195 205.555 ;
        RECT 14.485 205.385 14.655 205.555 ;
        RECT 14.945 205.385 15.115 205.555 ;
        RECT 15.405 205.385 15.575 205.555 ;
        RECT 15.865 205.385 16.035 205.555 ;
        RECT 16.325 205.385 16.495 205.555 ;
        RECT 16.785 205.385 16.955 205.555 ;
        RECT 17.245 205.385 17.415 205.555 ;
        RECT 17.705 205.385 17.875 205.555 ;
        RECT 18.165 205.385 18.335 205.555 ;
        RECT 18.625 205.385 18.795 205.555 ;
        RECT 19.085 205.385 19.255 205.555 ;
        RECT 19.545 205.385 19.715 205.555 ;
        RECT 20.005 205.385 20.175 205.555 ;
        RECT 20.465 205.385 20.635 205.555 ;
        RECT 20.925 205.385 21.095 205.555 ;
        RECT 21.385 205.385 21.555 205.555 ;
        RECT 21.845 205.385 22.015 205.555 ;
        RECT 22.305 205.385 22.475 205.555 ;
        RECT 22.765 205.385 22.935 205.555 ;
        RECT 23.225 205.385 23.395 205.555 ;
        RECT 23.685 205.385 23.855 205.555 ;
        RECT 24.145 205.385 24.315 205.555 ;
        RECT 24.605 205.385 24.775 205.555 ;
        RECT 25.065 205.385 25.235 205.555 ;
        RECT 25.525 205.385 25.695 205.555 ;
        RECT 25.985 205.385 26.155 205.555 ;
        RECT 26.445 205.385 26.615 205.555 ;
        RECT 26.905 205.385 27.075 205.555 ;
        RECT 27.365 205.385 27.535 205.555 ;
        RECT 27.825 205.385 27.995 205.555 ;
        RECT 28.285 205.385 28.455 205.555 ;
        RECT 28.745 205.385 28.915 205.555 ;
        RECT 29.205 205.385 29.375 205.555 ;
        RECT 29.665 205.385 29.835 205.555 ;
        RECT 30.125 205.385 30.295 205.555 ;
        RECT 30.585 205.385 30.755 205.555 ;
        RECT 31.045 205.385 31.215 205.555 ;
        RECT 31.505 205.385 31.675 205.555 ;
        RECT 31.965 205.385 32.135 205.555 ;
        RECT 32.425 205.385 32.595 205.555 ;
        RECT 32.885 205.385 33.055 205.555 ;
        RECT 33.345 205.385 33.515 205.555 ;
        RECT 33.805 205.385 33.975 205.555 ;
        RECT 34.265 205.385 34.435 205.555 ;
        RECT 34.725 205.385 34.895 205.555 ;
        RECT 35.185 205.385 35.355 205.555 ;
        RECT 35.645 205.385 35.815 205.555 ;
        RECT 36.105 205.385 36.275 205.555 ;
        RECT 36.565 205.385 36.735 205.555 ;
        RECT 37.025 205.385 37.195 205.555 ;
        RECT 37.485 205.385 37.655 205.555 ;
        RECT 37.945 205.385 38.115 205.555 ;
        RECT 38.405 205.385 38.575 205.555 ;
        RECT 38.865 205.385 39.035 205.555 ;
        RECT 39.325 205.385 39.495 205.555 ;
        RECT 39.785 205.385 39.955 205.555 ;
        RECT 40.245 205.385 40.415 205.555 ;
        RECT 40.705 205.385 40.875 205.555 ;
        RECT 41.165 205.385 41.335 205.555 ;
        RECT 41.625 205.385 41.795 205.555 ;
        RECT 42.085 205.385 42.255 205.555 ;
        RECT 42.545 205.385 42.715 205.555 ;
        RECT 43.005 205.385 43.175 205.555 ;
        RECT 43.465 205.385 43.635 205.555 ;
        RECT 43.925 205.385 44.095 205.555 ;
        RECT 44.385 205.385 44.555 205.555 ;
        RECT 44.845 205.385 45.015 205.555 ;
        RECT 45.305 205.385 45.475 205.555 ;
        RECT 45.765 205.385 45.935 205.555 ;
        RECT 46.225 205.385 46.395 205.555 ;
        RECT 46.685 205.385 46.855 205.555 ;
        RECT 47.145 205.385 47.315 205.555 ;
        RECT 47.605 205.385 47.775 205.555 ;
        RECT 48.065 205.385 48.235 205.555 ;
        RECT 48.525 205.385 48.695 205.555 ;
        RECT 48.985 205.385 49.155 205.555 ;
        RECT 49.445 205.385 49.615 205.555 ;
        RECT 49.905 205.385 50.075 205.555 ;
        RECT 50.365 205.385 50.535 205.555 ;
        RECT 50.825 205.385 50.995 205.555 ;
        RECT 51.285 205.385 51.455 205.555 ;
        RECT 51.745 205.385 51.915 205.555 ;
        RECT 52.205 205.385 52.375 205.555 ;
        RECT 52.665 205.385 52.835 205.555 ;
        RECT 53.125 205.385 53.295 205.555 ;
        RECT 53.585 205.385 53.755 205.555 ;
        RECT 54.045 205.385 54.215 205.555 ;
        RECT 54.505 205.385 54.675 205.555 ;
        RECT 54.965 205.385 55.135 205.555 ;
        RECT 55.425 205.385 55.595 205.555 ;
        RECT 55.885 205.385 56.055 205.555 ;
        RECT 56.345 205.385 56.515 205.555 ;
        RECT 56.805 205.385 56.975 205.555 ;
        RECT 57.265 205.385 57.435 205.555 ;
        RECT 57.725 205.385 57.895 205.555 ;
        RECT 58.185 205.385 58.355 205.555 ;
        RECT 58.645 205.385 58.815 205.555 ;
        RECT 59.105 205.385 59.275 205.555 ;
        RECT 59.565 205.385 59.735 205.555 ;
        RECT 60.025 205.385 60.195 205.555 ;
        RECT 60.485 205.385 60.655 205.555 ;
        RECT 60.945 205.385 61.115 205.555 ;
        RECT 61.405 205.385 61.575 205.555 ;
        RECT 61.865 205.385 62.035 205.555 ;
        RECT 62.325 205.385 62.495 205.555 ;
        RECT 62.785 205.385 62.955 205.555 ;
        RECT 63.245 205.385 63.415 205.555 ;
        RECT 63.705 205.385 63.875 205.555 ;
        RECT 64.165 205.385 64.335 205.555 ;
        RECT 64.625 205.385 64.795 205.555 ;
        RECT 65.085 205.385 65.255 205.555 ;
        RECT 65.545 205.385 65.715 205.555 ;
        RECT 66.005 205.385 66.175 205.555 ;
        RECT 66.465 205.385 66.635 205.555 ;
        RECT 66.925 205.385 67.095 205.555 ;
        RECT 67.385 205.385 67.555 205.555 ;
        RECT 67.845 205.385 68.015 205.555 ;
        RECT 68.305 205.385 68.475 205.555 ;
        RECT 68.765 205.385 68.935 205.555 ;
        RECT 69.225 205.385 69.395 205.555 ;
        RECT 69.685 205.385 69.855 205.555 ;
        RECT 70.145 205.385 70.315 205.555 ;
        RECT 70.605 205.385 70.775 205.555 ;
        RECT 71.065 205.385 71.235 205.555 ;
        RECT 71.525 205.385 71.695 205.555 ;
        RECT 71.985 205.385 72.155 205.555 ;
        RECT 72.445 205.385 72.615 205.555 ;
        RECT 72.905 205.385 73.075 205.555 ;
        RECT 73.365 205.385 73.535 205.555 ;
        RECT 73.825 205.385 73.995 205.555 ;
        RECT 74.285 205.385 74.455 205.555 ;
        RECT 74.745 205.385 74.915 205.555 ;
        RECT 75.205 205.385 75.375 205.555 ;
        RECT 75.665 205.385 75.835 205.555 ;
        RECT 76.125 205.385 76.295 205.555 ;
        RECT 76.585 205.385 76.755 205.555 ;
        RECT 77.045 205.385 77.215 205.555 ;
        RECT 77.505 205.385 77.675 205.555 ;
        RECT 77.965 205.385 78.135 205.555 ;
        RECT 78.425 205.385 78.595 205.555 ;
        RECT 78.885 205.385 79.055 205.555 ;
        RECT 79.345 205.385 79.515 205.555 ;
        RECT 79.805 205.385 79.975 205.555 ;
        RECT 80.265 205.385 80.435 205.555 ;
        RECT 80.725 205.385 80.895 205.555 ;
        RECT 81.185 205.385 81.355 205.555 ;
        RECT 81.645 205.385 81.815 205.555 ;
        RECT 82.105 205.385 82.275 205.555 ;
        RECT 82.565 205.385 82.735 205.555 ;
        RECT 83.025 205.385 83.195 205.555 ;
        RECT 83.485 205.385 83.655 205.555 ;
        RECT 83.945 205.385 84.115 205.555 ;
        RECT 84.405 205.385 84.575 205.555 ;
        RECT 84.865 205.385 85.035 205.555 ;
        RECT 85.325 205.385 85.495 205.555 ;
        RECT 85.785 205.385 85.955 205.555 ;
        RECT 86.245 205.385 86.415 205.555 ;
        RECT 86.705 205.385 86.875 205.555 ;
        RECT 87.165 205.385 87.335 205.555 ;
        RECT 87.625 205.385 87.795 205.555 ;
        RECT 88.085 205.385 88.255 205.555 ;
        RECT 88.545 205.385 88.715 205.555 ;
        RECT 89.005 205.385 89.175 205.555 ;
        RECT 89.465 205.385 89.635 205.555 ;
        RECT 89.925 205.385 90.095 205.555 ;
        RECT 90.385 205.385 90.555 205.555 ;
        RECT 90.845 205.385 91.015 205.555 ;
        RECT 91.305 205.385 91.475 205.555 ;
        RECT 91.765 205.385 91.935 205.555 ;
        RECT 92.225 205.385 92.395 205.555 ;
        RECT 92.685 205.385 92.855 205.555 ;
        RECT 93.145 205.385 93.315 205.555 ;
        RECT 93.605 205.385 93.775 205.555 ;
        RECT 94.065 205.385 94.235 205.555 ;
        RECT 94.525 205.385 94.695 205.555 ;
        RECT 94.985 205.385 95.155 205.555 ;
        RECT 95.445 205.385 95.615 205.555 ;
        RECT 95.905 205.385 96.075 205.555 ;
        RECT 96.365 205.385 96.535 205.555 ;
        RECT 96.825 205.385 96.995 205.555 ;
        RECT 97.285 205.385 97.455 205.555 ;
        RECT 97.745 205.385 97.915 205.555 ;
        RECT 98.205 205.385 98.375 205.555 ;
        RECT 98.665 205.385 98.835 205.555 ;
        RECT 99.125 205.385 99.295 205.555 ;
        RECT 99.585 205.385 99.755 205.555 ;
        RECT 100.045 205.385 100.215 205.555 ;
        RECT 100.505 205.385 100.675 205.555 ;
        RECT 100.965 205.385 101.135 205.555 ;
        RECT 101.425 205.385 101.595 205.555 ;
        RECT 101.885 205.385 102.055 205.555 ;
        RECT 102.345 205.385 102.515 205.555 ;
        RECT 102.805 205.385 102.975 205.555 ;
        RECT 103.265 205.385 103.435 205.555 ;
        RECT 103.725 205.385 103.895 205.555 ;
        RECT 104.185 205.385 104.355 205.555 ;
        RECT 104.645 205.385 104.815 205.555 ;
        RECT 105.105 205.385 105.275 205.555 ;
        RECT 105.565 205.385 105.735 205.555 ;
        RECT 106.025 205.385 106.195 205.555 ;
        RECT 106.485 205.385 106.655 205.555 ;
        RECT 106.945 205.385 107.115 205.555 ;
        RECT 107.405 205.385 107.575 205.555 ;
        RECT 107.865 205.385 108.035 205.555 ;
        RECT 108.325 205.385 108.495 205.555 ;
        RECT 108.785 205.385 108.955 205.555 ;
        RECT 109.245 205.385 109.415 205.555 ;
        RECT 109.705 205.385 109.875 205.555 ;
        RECT 110.165 205.385 110.335 205.555 ;
        RECT 110.625 205.385 110.795 205.555 ;
        RECT 111.085 205.385 111.255 205.555 ;
        RECT 111.545 205.385 111.715 205.555 ;
        RECT 112.005 205.385 112.175 205.555 ;
        RECT 112.465 205.385 112.635 205.555 ;
        RECT 112.925 205.385 113.095 205.555 ;
        RECT 113.385 205.385 113.555 205.555 ;
        RECT 113.845 205.385 114.015 205.555 ;
        RECT 114.305 205.385 114.475 205.555 ;
        RECT 114.765 205.385 114.935 205.555 ;
        RECT 115.225 205.385 115.395 205.555 ;
        RECT 115.685 205.385 115.855 205.555 ;
        RECT 116.145 205.385 116.315 205.555 ;
        RECT 116.605 205.385 116.775 205.555 ;
        RECT 117.065 205.385 117.235 205.555 ;
        RECT 117.525 205.385 117.695 205.555 ;
        RECT 117.985 205.385 118.155 205.555 ;
        RECT 118.445 205.385 118.615 205.555 ;
        RECT 118.905 205.385 119.075 205.555 ;
        RECT 119.365 205.385 119.535 205.555 ;
        RECT 119.825 205.385 119.995 205.555 ;
        RECT 120.285 205.385 120.455 205.555 ;
        RECT 120.745 205.385 120.915 205.555 ;
        RECT 121.205 205.385 121.375 205.555 ;
        RECT 121.665 205.385 121.835 205.555 ;
        RECT 122.125 205.385 122.295 205.555 ;
        RECT 122.585 205.385 122.755 205.555 ;
        RECT 123.045 205.385 123.215 205.555 ;
        RECT 123.505 205.385 123.675 205.555 ;
        RECT 123.965 205.385 124.135 205.555 ;
        RECT 124.425 205.385 124.595 205.555 ;
        RECT 124.885 205.385 125.055 205.555 ;
        RECT 125.345 205.385 125.515 205.555 ;
        RECT 125.805 205.385 125.975 205.555 ;
        RECT 126.265 205.385 126.435 205.555 ;
        RECT 126.725 205.385 126.895 205.555 ;
        RECT 127.185 205.385 127.355 205.555 ;
        RECT 127.645 205.385 127.815 205.555 ;
        RECT 128.105 205.385 128.275 205.555 ;
        RECT 128.565 205.385 128.735 205.555 ;
        RECT 129.025 205.385 129.195 205.555 ;
        RECT 129.485 205.385 129.655 205.555 ;
        RECT 129.945 205.385 130.115 205.555 ;
        RECT 130.405 205.385 130.575 205.555 ;
        RECT 130.865 205.385 131.035 205.555 ;
        RECT 131.325 205.385 131.495 205.555 ;
        RECT 131.785 205.385 131.955 205.555 ;
        RECT 132.245 205.385 132.415 205.555 ;
        RECT 132.705 205.385 132.875 205.555 ;
        RECT 133.165 205.385 133.335 205.555 ;
        RECT 133.625 205.385 133.795 205.555 ;
        RECT 134.085 205.385 134.255 205.555 ;
        RECT 134.545 205.385 134.715 205.555 ;
        RECT 135.005 205.385 135.175 205.555 ;
        RECT 135.465 205.385 135.635 205.555 ;
        RECT 135.925 205.385 136.095 205.555 ;
        RECT 136.385 205.385 136.555 205.555 ;
        RECT 136.845 205.385 137.015 205.555 ;
        RECT 137.305 205.385 137.475 205.555 ;
        RECT 137.765 205.385 137.935 205.555 ;
        RECT 138.225 205.385 138.395 205.555 ;
        RECT 138.685 205.385 138.855 205.555 ;
        RECT 139.145 205.385 139.315 205.555 ;
        RECT 139.605 205.385 139.775 205.555 ;
        RECT 140.065 205.385 140.235 205.555 ;
        RECT 140.525 205.385 140.695 205.555 ;
        RECT 140.985 205.385 141.155 205.555 ;
        RECT 141.445 205.385 141.615 205.555 ;
        RECT 141.905 205.385 142.075 205.555 ;
        RECT 142.365 205.385 142.535 205.555 ;
        RECT 142.825 205.385 142.995 205.555 ;
        RECT 143.285 205.385 143.455 205.555 ;
        RECT 143.745 205.385 143.915 205.555 ;
        RECT 144.205 205.385 144.375 205.555 ;
        RECT 144.665 205.385 144.835 205.555 ;
        RECT 145.125 205.385 145.295 205.555 ;
        RECT 145.585 205.385 145.755 205.555 ;
        RECT 146.045 205.385 146.215 205.555 ;
        RECT 146.505 205.385 146.675 205.555 ;
        RECT 146.965 205.385 147.135 205.555 ;
        RECT 147.425 205.385 147.595 205.555 ;
        RECT 147.885 205.385 148.055 205.555 ;
        RECT 148.345 205.385 148.515 205.555 ;
        RECT 148.805 205.385 148.975 205.555 ;
        RECT 149.265 205.385 149.435 205.555 ;
        RECT 149.725 205.385 149.895 205.555 ;
        RECT 150.185 205.385 150.355 205.555 ;
        RECT 30.125 204.535 30.295 204.705 ;
        RECT 31.175 204.875 31.345 205.045 ;
        RECT 38.865 204.875 39.035 205.045 ;
        RECT 31.965 203.515 32.135 203.685 ;
        RECT 31.045 203.175 31.215 203.345 ;
        RECT 39.785 203.515 39.955 203.685 ;
        RECT 45.305 204.875 45.475 205.045 ;
        RECT 41.165 203.855 41.335 204.025 ;
        RECT 44.845 204.195 45.015 204.365 ;
        RECT 45.765 204.195 45.935 204.365 ;
        RECT 46.225 204.195 46.395 204.365 ;
        RECT 47.145 204.875 47.315 205.045 ;
        RECT 48.525 204.875 48.695 205.045 ;
        RECT 47.605 204.195 47.775 204.365 ;
        RECT 48.065 204.195 48.235 204.365 ;
        RECT 48.985 204.195 49.155 204.365 ;
        RECT 46.225 203.515 46.395 203.685 ;
        RECT 54.965 204.195 55.135 204.365 ;
        RECT 54.505 203.855 54.675 204.025 ;
        RECT 56.805 203.515 56.975 203.685 ;
        RECT 60.485 204.875 60.655 205.045 ;
        RECT 58.645 204.195 58.815 204.365 ;
        RECT 58.185 203.855 58.355 204.025 ;
        RECT 69.225 204.195 69.395 204.365 ;
        RECT 70.605 204.195 70.775 204.365 ;
        RECT 71.065 204.195 71.235 204.365 ;
        RECT 71.985 203.855 72.155 204.025 ;
        RECT 77.505 204.535 77.675 204.705 ;
        RECT 79.345 204.875 79.515 205.045 ;
        RECT 78.655 204.365 78.825 204.535 ;
        RECT 82.105 204.875 82.275 205.045 ;
        RECT 82.565 204.875 82.735 205.045 ;
        RECT 81.185 204.195 81.355 204.365 ;
        RECT 80.265 203.855 80.435 204.025 ;
        RECT 78.425 203.175 78.595 203.345 ;
        RECT 82.565 203.855 82.735 204.025 ;
        RECT 83.945 204.195 84.115 204.365 ;
        RECT 83.485 203.855 83.655 204.025 ;
        RECT 90.845 204.195 91.015 204.365 ;
        RECT 91.330 203.515 91.500 203.685 ;
        RECT 91.725 203.855 91.895 204.025 ;
        RECT 92.125 204.195 92.295 204.365 ;
        RECT 92.915 203.855 93.085 204.025 ;
        RECT 93.430 203.515 93.600 203.685 ;
        RECT 95.000 203.515 95.170 203.685 ;
        RECT 95.435 203.855 95.605 204.025 ;
        RECT 97.745 203.515 97.915 203.685 ;
        RECT 106.945 203.515 107.115 203.685 ;
        RECT 109.255 203.855 109.425 204.025 ;
        RECT 109.690 203.515 109.860 203.685 ;
        RECT 111.775 203.855 111.945 204.025 ;
        RECT 111.260 203.515 111.430 203.685 ;
        RECT 112.510 204.195 112.680 204.365 ;
        RECT 112.965 203.855 113.135 204.025 ;
        RECT 113.845 203.855 114.015 204.025 ;
        RECT 113.360 203.515 113.530 203.685 ;
        RECT 11.265 202.665 11.435 202.835 ;
        RECT 11.725 202.665 11.895 202.835 ;
        RECT 12.185 202.665 12.355 202.835 ;
        RECT 12.645 202.665 12.815 202.835 ;
        RECT 13.105 202.665 13.275 202.835 ;
        RECT 13.565 202.665 13.735 202.835 ;
        RECT 14.025 202.665 14.195 202.835 ;
        RECT 14.485 202.665 14.655 202.835 ;
        RECT 14.945 202.665 15.115 202.835 ;
        RECT 15.405 202.665 15.575 202.835 ;
        RECT 15.865 202.665 16.035 202.835 ;
        RECT 16.325 202.665 16.495 202.835 ;
        RECT 16.785 202.665 16.955 202.835 ;
        RECT 17.245 202.665 17.415 202.835 ;
        RECT 17.705 202.665 17.875 202.835 ;
        RECT 18.165 202.665 18.335 202.835 ;
        RECT 18.625 202.665 18.795 202.835 ;
        RECT 19.085 202.665 19.255 202.835 ;
        RECT 19.545 202.665 19.715 202.835 ;
        RECT 20.005 202.665 20.175 202.835 ;
        RECT 20.465 202.665 20.635 202.835 ;
        RECT 20.925 202.665 21.095 202.835 ;
        RECT 21.385 202.665 21.555 202.835 ;
        RECT 21.845 202.665 22.015 202.835 ;
        RECT 22.305 202.665 22.475 202.835 ;
        RECT 22.765 202.665 22.935 202.835 ;
        RECT 23.225 202.665 23.395 202.835 ;
        RECT 23.685 202.665 23.855 202.835 ;
        RECT 24.145 202.665 24.315 202.835 ;
        RECT 24.605 202.665 24.775 202.835 ;
        RECT 25.065 202.665 25.235 202.835 ;
        RECT 25.525 202.665 25.695 202.835 ;
        RECT 25.985 202.665 26.155 202.835 ;
        RECT 26.445 202.665 26.615 202.835 ;
        RECT 26.905 202.665 27.075 202.835 ;
        RECT 27.365 202.665 27.535 202.835 ;
        RECT 27.825 202.665 27.995 202.835 ;
        RECT 28.285 202.665 28.455 202.835 ;
        RECT 28.745 202.665 28.915 202.835 ;
        RECT 29.205 202.665 29.375 202.835 ;
        RECT 29.665 202.665 29.835 202.835 ;
        RECT 30.125 202.665 30.295 202.835 ;
        RECT 30.585 202.665 30.755 202.835 ;
        RECT 31.045 202.665 31.215 202.835 ;
        RECT 31.505 202.665 31.675 202.835 ;
        RECT 31.965 202.665 32.135 202.835 ;
        RECT 32.425 202.665 32.595 202.835 ;
        RECT 32.885 202.665 33.055 202.835 ;
        RECT 33.345 202.665 33.515 202.835 ;
        RECT 33.805 202.665 33.975 202.835 ;
        RECT 34.265 202.665 34.435 202.835 ;
        RECT 34.725 202.665 34.895 202.835 ;
        RECT 35.185 202.665 35.355 202.835 ;
        RECT 35.645 202.665 35.815 202.835 ;
        RECT 36.105 202.665 36.275 202.835 ;
        RECT 36.565 202.665 36.735 202.835 ;
        RECT 37.025 202.665 37.195 202.835 ;
        RECT 37.485 202.665 37.655 202.835 ;
        RECT 37.945 202.665 38.115 202.835 ;
        RECT 38.405 202.665 38.575 202.835 ;
        RECT 38.865 202.665 39.035 202.835 ;
        RECT 39.325 202.665 39.495 202.835 ;
        RECT 39.785 202.665 39.955 202.835 ;
        RECT 40.245 202.665 40.415 202.835 ;
        RECT 40.705 202.665 40.875 202.835 ;
        RECT 41.165 202.665 41.335 202.835 ;
        RECT 41.625 202.665 41.795 202.835 ;
        RECT 42.085 202.665 42.255 202.835 ;
        RECT 42.545 202.665 42.715 202.835 ;
        RECT 43.005 202.665 43.175 202.835 ;
        RECT 43.465 202.665 43.635 202.835 ;
        RECT 43.925 202.665 44.095 202.835 ;
        RECT 44.385 202.665 44.555 202.835 ;
        RECT 44.845 202.665 45.015 202.835 ;
        RECT 45.305 202.665 45.475 202.835 ;
        RECT 45.765 202.665 45.935 202.835 ;
        RECT 46.225 202.665 46.395 202.835 ;
        RECT 46.685 202.665 46.855 202.835 ;
        RECT 47.145 202.665 47.315 202.835 ;
        RECT 47.605 202.665 47.775 202.835 ;
        RECT 48.065 202.665 48.235 202.835 ;
        RECT 48.525 202.665 48.695 202.835 ;
        RECT 48.985 202.665 49.155 202.835 ;
        RECT 49.445 202.665 49.615 202.835 ;
        RECT 49.905 202.665 50.075 202.835 ;
        RECT 50.365 202.665 50.535 202.835 ;
        RECT 50.825 202.665 50.995 202.835 ;
        RECT 51.285 202.665 51.455 202.835 ;
        RECT 51.745 202.665 51.915 202.835 ;
        RECT 52.205 202.665 52.375 202.835 ;
        RECT 52.665 202.665 52.835 202.835 ;
        RECT 53.125 202.665 53.295 202.835 ;
        RECT 53.585 202.665 53.755 202.835 ;
        RECT 54.045 202.665 54.215 202.835 ;
        RECT 54.505 202.665 54.675 202.835 ;
        RECT 54.965 202.665 55.135 202.835 ;
        RECT 55.425 202.665 55.595 202.835 ;
        RECT 55.885 202.665 56.055 202.835 ;
        RECT 56.345 202.665 56.515 202.835 ;
        RECT 56.805 202.665 56.975 202.835 ;
        RECT 57.265 202.665 57.435 202.835 ;
        RECT 57.725 202.665 57.895 202.835 ;
        RECT 58.185 202.665 58.355 202.835 ;
        RECT 58.645 202.665 58.815 202.835 ;
        RECT 59.105 202.665 59.275 202.835 ;
        RECT 59.565 202.665 59.735 202.835 ;
        RECT 60.025 202.665 60.195 202.835 ;
        RECT 60.485 202.665 60.655 202.835 ;
        RECT 60.945 202.665 61.115 202.835 ;
        RECT 61.405 202.665 61.575 202.835 ;
        RECT 61.865 202.665 62.035 202.835 ;
        RECT 62.325 202.665 62.495 202.835 ;
        RECT 62.785 202.665 62.955 202.835 ;
        RECT 63.245 202.665 63.415 202.835 ;
        RECT 63.705 202.665 63.875 202.835 ;
        RECT 64.165 202.665 64.335 202.835 ;
        RECT 64.625 202.665 64.795 202.835 ;
        RECT 65.085 202.665 65.255 202.835 ;
        RECT 65.545 202.665 65.715 202.835 ;
        RECT 66.005 202.665 66.175 202.835 ;
        RECT 66.465 202.665 66.635 202.835 ;
        RECT 66.925 202.665 67.095 202.835 ;
        RECT 67.385 202.665 67.555 202.835 ;
        RECT 67.845 202.665 68.015 202.835 ;
        RECT 68.305 202.665 68.475 202.835 ;
        RECT 68.765 202.665 68.935 202.835 ;
        RECT 69.225 202.665 69.395 202.835 ;
        RECT 69.685 202.665 69.855 202.835 ;
        RECT 70.145 202.665 70.315 202.835 ;
        RECT 70.605 202.665 70.775 202.835 ;
        RECT 71.065 202.665 71.235 202.835 ;
        RECT 71.525 202.665 71.695 202.835 ;
        RECT 71.985 202.665 72.155 202.835 ;
        RECT 72.445 202.665 72.615 202.835 ;
        RECT 72.905 202.665 73.075 202.835 ;
        RECT 73.365 202.665 73.535 202.835 ;
        RECT 73.825 202.665 73.995 202.835 ;
        RECT 74.285 202.665 74.455 202.835 ;
        RECT 74.745 202.665 74.915 202.835 ;
        RECT 75.205 202.665 75.375 202.835 ;
        RECT 75.665 202.665 75.835 202.835 ;
        RECT 76.125 202.665 76.295 202.835 ;
        RECT 76.585 202.665 76.755 202.835 ;
        RECT 77.045 202.665 77.215 202.835 ;
        RECT 77.505 202.665 77.675 202.835 ;
        RECT 77.965 202.665 78.135 202.835 ;
        RECT 78.425 202.665 78.595 202.835 ;
        RECT 78.885 202.665 79.055 202.835 ;
        RECT 79.345 202.665 79.515 202.835 ;
        RECT 79.805 202.665 79.975 202.835 ;
        RECT 80.265 202.665 80.435 202.835 ;
        RECT 80.725 202.665 80.895 202.835 ;
        RECT 81.185 202.665 81.355 202.835 ;
        RECT 81.645 202.665 81.815 202.835 ;
        RECT 82.105 202.665 82.275 202.835 ;
        RECT 82.565 202.665 82.735 202.835 ;
        RECT 83.025 202.665 83.195 202.835 ;
        RECT 83.485 202.665 83.655 202.835 ;
        RECT 83.945 202.665 84.115 202.835 ;
        RECT 84.405 202.665 84.575 202.835 ;
        RECT 84.865 202.665 85.035 202.835 ;
        RECT 85.325 202.665 85.495 202.835 ;
        RECT 85.785 202.665 85.955 202.835 ;
        RECT 86.245 202.665 86.415 202.835 ;
        RECT 86.705 202.665 86.875 202.835 ;
        RECT 87.165 202.665 87.335 202.835 ;
        RECT 87.625 202.665 87.795 202.835 ;
        RECT 88.085 202.665 88.255 202.835 ;
        RECT 88.545 202.665 88.715 202.835 ;
        RECT 89.005 202.665 89.175 202.835 ;
        RECT 89.465 202.665 89.635 202.835 ;
        RECT 89.925 202.665 90.095 202.835 ;
        RECT 90.385 202.665 90.555 202.835 ;
        RECT 90.845 202.665 91.015 202.835 ;
        RECT 91.305 202.665 91.475 202.835 ;
        RECT 91.765 202.665 91.935 202.835 ;
        RECT 92.225 202.665 92.395 202.835 ;
        RECT 92.685 202.665 92.855 202.835 ;
        RECT 93.145 202.665 93.315 202.835 ;
        RECT 93.605 202.665 93.775 202.835 ;
        RECT 94.065 202.665 94.235 202.835 ;
        RECT 94.525 202.665 94.695 202.835 ;
        RECT 94.985 202.665 95.155 202.835 ;
        RECT 95.445 202.665 95.615 202.835 ;
        RECT 95.905 202.665 96.075 202.835 ;
        RECT 96.365 202.665 96.535 202.835 ;
        RECT 96.825 202.665 96.995 202.835 ;
        RECT 97.285 202.665 97.455 202.835 ;
        RECT 97.745 202.665 97.915 202.835 ;
        RECT 98.205 202.665 98.375 202.835 ;
        RECT 98.665 202.665 98.835 202.835 ;
        RECT 99.125 202.665 99.295 202.835 ;
        RECT 99.585 202.665 99.755 202.835 ;
        RECT 100.045 202.665 100.215 202.835 ;
        RECT 100.505 202.665 100.675 202.835 ;
        RECT 100.965 202.665 101.135 202.835 ;
        RECT 101.425 202.665 101.595 202.835 ;
        RECT 101.885 202.665 102.055 202.835 ;
        RECT 102.345 202.665 102.515 202.835 ;
        RECT 102.805 202.665 102.975 202.835 ;
        RECT 103.265 202.665 103.435 202.835 ;
        RECT 103.725 202.665 103.895 202.835 ;
        RECT 104.185 202.665 104.355 202.835 ;
        RECT 104.645 202.665 104.815 202.835 ;
        RECT 105.105 202.665 105.275 202.835 ;
        RECT 105.565 202.665 105.735 202.835 ;
        RECT 106.025 202.665 106.195 202.835 ;
        RECT 106.485 202.665 106.655 202.835 ;
        RECT 106.945 202.665 107.115 202.835 ;
        RECT 107.405 202.665 107.575 202.835 ;
        RECT 107.865 202.665 108.035 202.835 ;
        RECT 108.325 202.665 108.495 202.835 ;
        RECT 108.785 202.665 108.955 202.835 ;
        RECT 109.245 202.665 109.415 202.835 ;
        RECT 109.705 202.665 109.875 202.835 ;
        RECT 110.165 202.665 110.335 202.835 ;
        RECT 110.625 202.665 110.795 202.835 ;
        RECT 111.085 202.665 111.255 202.835 ;
        RECT 111.545 202.665 111.715 202.835 ;
        RECT 112.005 202.665 112.175 202.835 ;
        RECT 112.465 202.665 112.635 202.835 ;
        RECT 112.925 202.665 113.095 202.835 ;
        RECT 113.385 202.665 113.555 202.835 ;
        RECT 113.845 202.665 114.015 202.835 ;
        RECT 114.305 202.665 114.475 202.835 ;
        RECT 114.765 202.665 114.935 202.835 ;
        RECT 115.225 202.665 115.395 202.835 ;
        RECT 115.685 202.665 115.855 202.835 ;
        RECT 116.145 202.665 116.315 202.835 ;
        RECT 116.605 202.665 116.775 202.835 ;
        RECT 117.065 202.665 117.235 202.835 ;
        RECT 117.525 202.665 117.695 202.835 ;
        RECT 117.985 202.665 118.155 202.835 ;
        RECT 118.445 202.665 118.615 202.835 ;
        RECT 118.905 202.665 119.075 202.835 ;
        RECT 119.365 202.665 119.535 202.835 ;
        RECT 119.825 202.665 119.995 202.835 ;
        RECT 120.285 202.665 120.455 202.835 ;
        RECT 120.745 202.665 120.915 202.835 ;
        RECT 121.205 202.665 121.375 202.835 ;
        RECT 121.665 202.665 121.835 202.835 ;
        RECT 122.125 202.665 122.295 202.835 ;
        RECT 122.585 202.665 122.755 202.835 ;
        RECT 123.045 202.665 123.215 202.835 ;
        RECT 123.505 202.665 123.675 202.835 ;
        RECT 123.965 202.665 124.135 202.835 ;
        RECT 124.425 202.665 124.595 202.835 ;
        RECT 124.885 202.665 125.055 202.835 ;
        RECT 125.345 202.665 125.515 202.835 ;
        RECT 125.805 202.665 125.975 202.835 ;
        RECT 126.265 202.665 126.435 202.835 ;
        RECT 126.725 202.665 126.895 202.835 ;
        RECT 127.185 202.665 127.355 202.835 ;
        RECT 127.645 202.665 127.815 202.835 ;
        RECT 128.105 202.665 128.275 202.835 ;
        RECT 128.565 202.665 128.735 202.835 ;
        RECT 129.025 202.665 129.195 202.835 ;
        RECT 129.485 202.665 129.655 202.835 ;
        RECT 129.945 202.665 130.115 202.835 ;
        RECT 130.405 202.665 130.575 202.835 ;
        RECT 130.865 202.665 131.035 202.835 ;
        RECT 131.325 202.665 131.495 202.835 ;
        RECT 131.785 202.665 131.955 202.835 ;
        RECT 132.245 202.665 132.415 202.835 ;
        RECT 132.705 202.665 132.875 202.835 ;
        RECT 133.165 202.665 133.335 202.835 ;
        RECT 133.625 202.665 133.795 202.835 ;
        RECT 134.085 202.665 134.255 202.835 ;
        RECT 134.545 202.665 134.715 202.835 ;
        RECT 135.005 202.665 135.175 202.835 ;
        RECT 135.465 202.665 135.635 202.835 ;
        RECT 135.925 202.665 136.095 202.835 ;
        RECT 136.385 202.665 136.555 202.835 ;
        RECT 136.845 202.665 137.015 202.835 ;
        RECT 137.305 202.665 137.475 202.835 ;
        RECT 137.765 202.665 137.935 202.835 ;
        RECT 138.225 202.665 138.395 202.835 ;
        RECT 138.685 202.665 138.855 202.835 ;
        RECT 139.145 202.665 139.315 202.835 ;
        RECT 139.605 202.665 139.775 202.835 ;
        RECT 140.065 202.665 140.235 202.835 ;
        RECT 140.525 202.665 140.695 202.835 ;
        RECT 140.985 202.665 141.155 202.835 ;
        RECT 141.445 202.665 141.615 202.835 ;
        RECT 141.905 202.665 142.075 202.835 ;
        RECT 142.365 202.665 142.535 202.835 ;
        RECT 142.825 202.665 142.995 202.835 ;
        RECT 143.285 202.665 143.455 202.835 ;
        RECT 143.745 202.665 143.915 202.835 ;
        RECT 144.205 202.665 144.375 202.835 ;
        RECT 144.665 202.665 144.835 202.835 ;
        RECT 145.125 202.665 145.295 202.835 ;
        RECT 145.585 202.665 145.755 202.835 ;
        RECT 146.045 202.665 146.215 202.835 ;
        RECT 146.505 202.665 146.675 202.835 ;
        RECT 146.965 202.665 147.135 202.835 ;
        RECT 147.425 202.665 147.595 202.835 ;
        RECT 147.885 202.665 148.055 202.835 ;
        RECT 148.345 202.665 148.515 202.835 ;
        RECT 148.805 202.665 148.975 202.835 ;
        RECT 149.265 202.665 149.435 202.835 ;
        RECT 149.725 202.665 149.895 202.835 ;
        RECT 150.185 202.665 150.355 202.835 ;
        RECT 17.270 201.815 17.440 201.985 ;
        RECT 16.785 201.135 16.955 201.305 ;
        RECT 17.665 201.475 17.835 201.645 ;
        RECT 18.120 200.795 18.290 200.965 ;
        RECT 19.370 201.815 19.540 201.985 ;
        RECT 18.855 201.475 19.025 201.645 ;
        RECT 20.940 201.815 21.110 201.985 ;
        RECT 21.375 201.475 21.545 201.645 ;
        RECT 23.685 201.815 23.855 201.985 ;
        RECT 24.605 200.455 24.775 200.625 ;
        RECT 29.690 201.815 29.860 201.985 ;
        RECT 27.365 201.475 27.535 201.645 ;
        RECT 29.205 201.135 29.375 201.305 ;
        RECT 30.085 201.475 30.255 201.645 ;
        RECT 30.540 200.795 30.710 200.965 ;
        RECT 31.790 201.815 31.960 201.985 ;
        RECT 31.275 201.475 31.445 201.645 ;
        RECT 33.360 201.815 33.530 201.985 ;
        RECT 33.795 201.475 33.965 201.645 ;
        RECT 38.405 202.155 38.575 202.325 ;
        RECT 37.485 201.135 37.655 201.305 ;
        RECT 36.105 200.455 36.275 200.625 ;
        RECT 39.785 200.455 39.955 200.625 ;
        RECT 40.245 202.155 40.415 202.325 ;
        RECT 40.705 201.815 40.875 201.985 ;
        RECT 43.005 201.815 43.175 201.985 ;
        RECT 42.545 200.795 42.715 200.965 ;
        RECT 43.005 201.135 43.175 201.305 ;
        RECT 44.385 201.135 44.555 201.305 ;
        RECT 43.925 200.455 44.095 200.625 ;
        RECT 50.365 202.155 50.535 202.325 ;
        RECT 51.285 201.135 51.455 201.305 ;
        RECT 52.665 201.135 52.835 201.305 ;
        RECT 52.205 200.455 52.375 200.625 ;
        RECT 63.245 201.815 63.415 201.985 ;
        RECT 67.845 202.155 68.015 202.325 ;
        RECT 65.085 201.135 65.255 201.305 ;
        RECT 64.165 200.455 64.335 200.625 ;
        RECT 66.465 201.135 66.635 201.305 ;
        RECT 66.005 200.455 66.175 200.625 ;
        RECT 69.225 201.135 69.395 201.305 ;
        RECT 66.925 200.455 67.095 200.625 ;
        RECT 71.065 202.155 71.235 202.325 ;
        RECT 73.825 202.155 73.995 202.325 ;
        RECT 71.985 200.795 72.155 200.965 ;
        RECT 72.905 201.135 73.075 201.305 ;
        RECT 73.365 201.135 73.535 201.305 ;
        RECT 74.285 201.135 74.455 201.305 ;
        RECT 83.025 201.135 83.195 201.305 ;
        RECT 84.865 202.155 85.035 202.325 ;
        RECT 85.785 201.815 85.955 201.985 ;
        RECT 84.865 200.455 85.035 200.625 ;
        RECT 89.925 202.155 90.095 202.325 ;
        RECT 89.005 201.135 89.175 201.305 ;
        RECT 100.045 201.135 100.215 201.305 ;
        RECT 100.965 200.455 101.135 200.625 ;
        RECT 101.885 200.455 102.055 200.625 ;
        RECT 104.195 201.475 104.365 201.645 ;
        RECT 104.630 201.815 104.800 201.985 ;
        RECT 106.200 201.815 106.370 201.985 ;
        RECT 106.715 201.475 106.885 201.645 ;
        RECT 107.450 200.795 107.620 200.965 ;
        RECT 107.905 201.475 108.075 201.645 ;
        RECT 108.300 201.815 108.470 201.985 ;
        RECT 108.785 201.135 108.955 201.305 ;
        RECT 110.165 201.135 110.335 201.305 ;
        RECT 112.925 202.155 113.095 202.325 ;
        RECT 115.250 201.815 115.420 201.985 ;
        RECT 114.765 201.475 114.935 201.645 ;
        RECT 115.645 201.475 115.815 201.645 ;
        RECT 116.100 200.795 116.270 200.965 ;
        RECT 117.350 201.815 117.520 201.985 ;
        RECT 116.835 201.475 117.005 201.645 ;
        RECT 118.920 201.815 119.090 201.985 ;
        RECT 119.355 201.475 119.525 201.645 ;
        RECT 121.665 200.455 121.835 200.625 ;
        RECT 11.265 199.945 11.435 200.115 ;
        RECT 11.725 199.945 11.895 200.115 ;
        RECT 12.185 199.945 12.355 200.115 ;
        RECT 12.645 199.945 12.815 200.115 ;
        RECT 13.105 199.945 13.275 200.115 ;
        RECT 13.565 199.945 13.735 200.115 ;
        RECT 14.025 199.945 14.195 200.115 ;
        RECT 14.485 199.945 14.655 200.115 ;
        RECT 14.945 199.945 15.115 200.115 ;
        RECT 15.405 199.945 15.575 200.115 ;
        RECT 15.865 199.945 16.035 200.115 ;
        RECT 16.325 199.945 16.495 200.115 ;
        RECT 16.785 199.945 16.955 200.115 ;
        RECT 17.245 199.945 17.415 200.115 ;
        RECT 17.705 199.945 17.875 200.115 ;
        RECT 18.165 199.945 18.335 200.115 ;
        RECT 18.625 199.945 18.795 200.115 ;
        RECT 19.085 199.945 19.255 200.115 ;
        RECT 19.545 199.945 19.715 200.115 ;
        RECT 20.005 199.945 20.175 200.115 ;
        RECT 20.465 199.945 20.635 200.115 ;
        RECT 20.925 199.945 21.095 200.115 ;
        RECT 21.385 199.945 21.555 200.115 ;
        RECT 21.845 199.945 22.015 200.115 ;
        RECT 22.305 199.945 22.475 200.115 ;
        RECT 22.765 199.945 22.935 200.115 ;
        RECT 23.225 199.945 23.395 200.115 ;
        RECT 23.685 199.945 23.855 200.115 ;
        RECT 24.145 199.945 24.315 200.115 ;
        RECT 24.605 199.945 24.775 200.115 ;
        RECT 25.065 199.945 25.235 200.115 ;
        RECT 25.525 199.945 25.695 200.115 ;
        RECT 25.985 199.945 26.155 200.115 ;
        RECT 26.445 199.945 26.615 200.115 ;
        RECT 26.905 199.945 27.075 200.115 ;
        RECT 27.365 199.945 27.535 200.115 ;
        RECT 27.825 199.945 27.995 200.115 ;
        RECT 28.285 199.945 28.455 200.115 ;
        RECT 28.745 199.945 28.915 200.115 ;
        RECT 29.205 199.945 29.375 200.115 ;
        RECT 29.665 199.945 29.835 200.115 ;
        RECT 30.125 199.945 30.295 200.115 ;
        RECT 30.585 199.945 30.755 200.115 ;
        RECT 31.045 199.945 31.215 200.115 ;
        RECT 31.505 199.945 31.675 200.115 ;
        RECT 31.965 199.945 32.135 200.115 ;
        RECT 32.425 199.945 32.595 200.115 ;
        RECT 32.885 199.945 33.055 200.115 ;
        RECT 33.345 199.945 33.515 200.115 ;
        RECT 33.805 199.945 33.975 200.115 ;
        RECT 34.265 199.945 34.435 200.115 ;
        RECT 34.725 199.945 34.895 200.115 ;
        RECT 35.185 199.945 35.355 200.115 ;
        RECT 35.645 199.945 35.815 200.115 ;
        RECT 36.105 199.945 36.275 200.115 ;
        RECT 36.565 199.945 36.735 200.115 ;
        RECT 37.025 199.945 37.195 200.115 ;
        RECT 37.485 199.945 37.655 200.115 ;
        RECT 37.945 199.945 38.115 200.115 ;
        RECT 38.405 199.945 38.575 200.115 ;
        RECT 38.865 199.945 39.035 200.115 ;
        RECT 39.325 199.945 39.495 200.115 ;
        RECT 39.785 199.945 39.955 200.115 ;
        RECT 40.245 199.945 40.415 200.115 ;
        RECT 40.705 199.945 40.875 200.115 ;
        RECT 41.165 199.945 41.335 200.115 ;
        RECT 41.625 199.945 41.795 200.115 ;
        RECT 42.085 199.945 42.255 200.115 ;
        RECT 42.545 199.945 42.715 200.115 ;
        RECT 43.005 199.945 43.175 200.115 ;
        RECT 43.465 199.945 43.635 200.115 ;
        RECT 43.925 199.945 44.095 200.115 ;
        RECT 44.385 199.945 44.555 200.115 ;
        RECT 44.845 199.945 45.015 200.115 ;
        RECT 45.305 199.945 45.475 200.115 ;
        RECT 45.765 199.945 45.935 200.115 ;
        RECT 46.225 199.945 46.395 200.115 ;
        RECT 46.685 199.945 46.855 200.115 ;
        RECT 47.145 199.945 47.315 200.115 ;
        RECT 47.605 199.945 47.775 200.115 ;
        RECT 48.065 199.945 48.235 200.115 ;
        RECT 48.525 199.945 48.695 200.115 ;
        RECT 48.985 199.945 49.155 200.115 ;
        RECT 49.445 199.945 49.615 200.115 ;
        RECT 49.905 199.945 50.075 200.115 ;
        RECT 50.365 199.945 50.535 200.115 ;
        RECT 50.825 199.945 50.995 200.115 ;
        RECT 51.285 199.945 51.455 200.115 ;
        RECT 51.745 199.945 51.915 200.115 ;
        RECT 52.205 199.945 52.375 200.115 ;
        RECT 52.665 199.945 52.835 200.115 ;
        RECT 53.125 199.945 53.295 200.115 ;
        RECT 53.585 199.945 53.755 200.115 ;
        RECT 54.045 199.945 54.215 200.115 ;
        RECT 54.505 199.945 54.675 200.115 ;
        RECT 54.965 199.945 55.135 200.115 ;
        RECT 55.425 199.945 55.595 200.115 ;
        RECT 55.885 199.945 56.055 200.115 ;
        RECT 56.345 199.945 56.515 200.115 ;
        RECT 56.805 199.945 56.975 200.115 ;
        RECT 57.265 199.945 57.435 200.115 ;
        RECT 57.725 199.945 57.895 200.115 ;
        RECT 58.185 199.945 58.355 200.115 ;
        RECT 58.645 199.945 58.815 200.115 ;
        RECT 59.105 199.945 59.275 200.115 ;
        RECT 59.565 199.945 59.735 200.115 ;
        RECT 60.025 199.945 60.195 200.115 ;
        RECT 60.485 199.945 60.655 200.115 ;
        RECT 60.945 199.945 61.115 200.115 ;
        RECT 61.405 199.945 61.575 200.115 ;
        RECT 61.865 199.945 62.035 200.115 ;
        RECT 62.325 199.945 62.495 200.115 ;
        RECT 62.785 199.945 62.955 200.115 ;
        RECT 63.245 199.945 63.415 200.115 ;
        RECT 63.705 199.945 63.875 200.115 ;
        RECT 64.165 199.945 64.335 200.115 ;
        RECT 64.625 199.945 64.795 200.115 ;
        RECT 65.085 199.945 65.255 200.115 ;
        RECT 65.545 199.945 65.715 200.115 ;
        RECT 66.005 199.945 66.175 200.115 ;
        RECT 66.465 199.945 66.635 200.115 ;
        RECT 66.925 199.945 67.095 200.115 ;
        RECT 67.385 199.945 67.555 200.115 ;
        RECT 67.845 199.945 68.015 200.115 ;
        RECT 68.305 199.945 68.475 200.115 ;
        RECT 68.765 199.945 68.935 200.115 ;
        RECT 69.225 199.945 69.395 200.115 ;
        RECT 69.685 199.945 69.855 200.115 ;
        RECT 70.145 199.945 70.315 200.115 ;
        RECT 70.605 199.945 70.775 200.115 ;
        RECT 71.065 199.945 71.235 200.115 ;
        RECT 71.525 199.945 71.695 200.115 ;
        RECT 71.985 199.945 72.155 200.115 ;
        RECT 72.445 199.945 72.615 200.115 ;
        RECT 72.905 199.945 73.075 200.115 ;
        RECT 73.365 199.945 73.535 200.115 ;
        RECT 73.825 199.945 73.995 200.115 ;
        RECT 74.285 199.945 74.455 200.115 ;
        RECT 74.745 199.945 74.915 200.115 ;
        RECT 75.205 199.945 75.375 200.115 ;
        RECT 75.665 199.945 75.835 200.115 ;
        RECT 76.125 199.945 76.295 200.115 ;
        RECT 76.585 199.945 76.755 200.115 ;
        RECT 77.045 199.945 77.215 200.115 ;
        RECT 77.505 199.945 77.675 200.115 ;
        RECT 77.965 199.945 78.135 200.115 ;
        RECT 78.425 199.945 78.595 200.115 ;
        RECT 78.885 199.945 79.055 200.115 ;
        RECT 79.345 199.945 79.515 200.115 ;
        RECT 79.805 199.945 79.975 200.115 ;
        RECT 80.265 199.945 80.435 200.115 ;
        RECT 80.725 199.945 80.895 200.115 ;
        RECT 81.185 199.945 81.355 200.115 ;
        RECT 81.645 199.945 81.815 200.115 ;
        RECT 82.105 199.945 82.275 200.115 ;
        RECT 82.565 199.945 82.735 200.115 ;
        RECT 83.025 199.945 83.195 200.115 ;
        RECT 83.485 199.945 83.655 200.115 ;
        RECT 83.945 199.945 84.115 200.115 ;
        RECT 84.405 199.945 84.575 200.115 ;
        RECT 84.865 199.945 85.035 200.115 ;
        RECT 85.325 199.945 85.495 200.115 ;
        RECT 85.785 199.945 85.955 200.115 ;
        RECT 86.245 199.945 86.415 200.115 ;
        RECT 86.705 199.945 86.875 200.115 ;
        RECT 87.165 199.945 87.335 200.115 ;
        RECT 87.625 199.945 87.795 200.115 ;
        RECT 88.085 199.945 88.255 200.115 ;
        RECT 88.545 199.945 88.715 200.115 ;
        RECT 89.005 199.945 89.175 200.115 ;
        RECT 89.465 199.945 89.635 200.115 ;
        RECT 89.925 199.945 90.095 200.115 ;
        RECT 90.385 199.945 90.555 200.115 ;
        RECT 90.845 199.945 91.015 200.115 ;
        RECT 91.305 199.945 91.475 200.115 ;
        RECT 91.765 199.945 91.935 200.115 ;
        RECT 92.225 199.945 92.395 200.115 ;
        RECT 92.685 199.945 92.855 200.115 ;
        RECT 93.145 199.945 93.315 200.115 ;
        RECT 93.605 199.945 93.775 200.115 ;
        RECT 94.065 199.945 94.235 200.115 ;
        RECT 94.525 199.945 94.695 200.115 ;
        RECT 94.985 199.945 95.155 200.115 ;
        RECT 95.445 199.945 95.615 200.115 ;
        RECT 95.905 199.945 96.075 200.115 ;
        RECT 96.365 199.945 96.535 200.115 ;
        RECT 96.825 199.945 96.995 200.115 ;
        RECT 97.285 199.945 97.455 200.115 ;
        RECT 97.745 199.945 97.915 200.115 ;
        RECT 98.205 199.945 98.375 200.115 ;
        RECT 98.665 199.945 98.835 200.115 ;
        RECT 99.125 199.945 99.295 200.115 ;
        RECT 99.585 199.945 99.755 200.115 ;
        RECT 100.045 199.945 100.215 200.115 ;
        RECT 100.505 199.945 100.675 200.115 ;
        RECT 100.965 199.945 101.135 200.115 ;
        RECT 101.425 199.945 101.595 200.115 ;
        RECT 101.885 199.945 102.055 200.115 ;
        RECT 102.345 199.945 102.515 200.115 ;
        RECT 102.805 199.945 102.975 200.115 ;
        RECT 103.265 199.945 103.435 200.115 ;
        RECT 103.725 199.945 103.895 200.115 ;
        RECT 104.185 199.945 104.355 200.115 ;
        RECT 104.645 199.945 104.815 200.115 ;
        RECT 105.105 199.945 105.275 200.115 ;
        RECT 105.565 199.945 105.735 200.115 ;
        RECT 106.025 199.945 106.195 200.115 ;
        RECT 106.485 199.945 106.655 200.115 ;
        RECT 106.945 199.945 107.115 200.115 ;
        RECT 107.405 199.945 107.575 200.115 ;
        RECT 107.865 199.945 108.035 200.115 ;
        RECT 108.325 199.945 108.495 200.115 ;
        RECT 108.785 199.945 108.955 200.115 ;
        RECT 109.245 199.945 109.415 200.115 ;
        RECT 109.705 199.945 109.875 200.115 ;
        RECT 110.165 199.945 110.335 200.115 ;
        RECT 110.625 199.945 110.795 200.115 ;
        RECT 111.085 199.945 111.255 200.115 ;
        RECT 111.545 199.945 111.715 200.115 ;
        RECT 112.005 199.945 112.175 200.115 ;
        RECT 112.465 199.945 112.635 200.115 ;
        RECT 112.925 199.945 113.095 200.115 ;
        RECT 113.385 199.945 113.555 200.115 ;
        RECT 113.845 199.945 114.015 200.115 ;
        RECT 114.305 199.945 114.475 200.115 ;
        RECT 114.765 199.945 114.935 200.115 ;
        RECT 115.225 199.945 115.395 200.115 ;
        RECT 115.685 199.945 115.855 200.115 ;
        RECT 116.145 199.945 116.315 200.115 ;
        RECT 116.605 199.945 116.775 200.115 ;
        RECT 117.065 199.945 117.235 200.115 ;
        RECT 117.525 199.945 117.695 200.115 ;
        RECT 117.985 199.945 118.155 200.115 ;
        RECT 118.445 199.945 118.615 200.115 ;
        RECT 118.905 199.945 119.075 200.115 ;
        RECT 119.365 199.945 119.535 200.115 ;
        RECT 119.825 199.945 119.995 200.115 ;
        RECT 120.285 199.945 120.455 200.115 ;
        RECT 120.745 199.945 120.915 200.115 ;
        RECT 121.205 199.945 121.375 200.115 ;
        RECT 121.665 199.945 121.835 200.115 ;
        RECT 122.125 199.945 122.295 200.115 ;
        RECT 122.585 199.945 122.755 200.115 ;
        RECT 123.045 199.945 123.215 200.115 ;
        RECT 123.505 199.945 123.675 200.115 ;
        RECT 123.965 199.945 124.135 200.115 ;
        RECT 124.425 199.945 124.595 200.115 ;
        RECT 124.885 199.945 125.055 200.115 ;
        RECT 125.345 199.945 125.515 200.115 ;
        RECT 125.805 199.945 125.975 200.115 ;
        RECT 126.265 199.945 126.435 200.115 ;
        RECT 126.725 199.945 126.895 200.115 ;
        RECT 127.185 199.945 127.355 200.115 ;
        RECT 127.645 199.945 127.815 200.115 ;
        RECT 128.105 199.945 128.275 200.115 ;
        RECT 128.565 199.945 128.735 200.115 ;
        RECT 129.025 199.945 129.195 200.115 ;
        RECT 129.485 199.945 129.655 200.115 ;
        RECT 129.945 199.945 130.115 200.115 ;
        RECT 130.405 199.945 130.575 200.115 ;
        RECT 130.865 199.945 131.035 200.115 ;
        RECT 131.325 199.945 131.495 200.115 ;
        RECT 131.785 199.945 131.955 200.115 ;
        RECT 132.245 199.945 132.415 200.115 ;
        RECT 132.705 199.945 132.875 200.115 ;
        RECT 133.165 199.945 133.335 200.115 ;
        RECT 133.625 199.945 133.795 200.115 ;
        RECT 134.085 199.945 134.255 200.115 ;
        RECT 134.545 199.945 134.715 200.115 ;
        RECT 135.005 199.945 135.175 200.115 ;
        RECT 135.465 199.945 135.635 200.115 ;
        RECT 135.925 199.945 136.095 200.115 ;
        RECT 136.385 199.945 136.555 200.115 ;
        RECT 136.845 199.945 137.015 200.115 ;
        RECT 137.305 199.945 137.475 200.115 ;
        RECT 137.765 199.945 137.935 200.115 ;
        RECT 138.225 199.945 138.395 200.115 ;
        RECT 138.685 199.945 138.855 200.115 ;
        RECT 139.145 199.945 139.315 200.115 ;
        RECT 139.605 199.945 139.775 200.115 ;
        RECT 140.065 199.945 140.235 200.115 ;
        RECT 140.525 199.945 140.695 200.115 ;
        RECT 140.985 199.945 141.155 200.115 ;
        RECT 141.445 199.945 141.615 200.115 ;
        RECT 141.905 199.945 142.075 200.115 ;
        RECT 142.365 199.945 142.535 200.115 ;
        RECT 142.825 199.945 142.995 200.115 ;
        RECT 143.285 199.945 143.455 200.115 ;
        RECT 143.745 199.945 143.915 200.115 ;
        RECT 144.205 199.945 144.375 200.115 ;
        RECT 144.665 199.945 144.835 200.115 ;
        RECT 145.125 199.945 145.295 200.115 ;
        RECT 145.585 199.945 145.755 200.115 ;
        RECT 146.045 199.945 146.215 200.115 ;
        RECT 146.505 199.945 146.675 200.115 ;
        RECT 146.965 199.945 147.135 200.115 ;
        RECT 147.425 199.945 147.595 200.115 ;
        RECT 147.885 199.945 148.055 200.115 ;
        RECT 148.345 199.945 148.515 200.115 ;
        RECT 148.805 199.945 148.975 200.115 ;
        RECT 149.265 199.945 149.435 200.115 ;
        RECT 149.725 199.945 149.895 200.115 ;
        RECT 150.185 199.945 150.355 200.115 ;
        RECT 23.225 198.755 23.395 198.925 ;
        RECT 24.145 199.435 24.315 199.605 ;
        RECT 24.605 198.755 24.775 198.925 ;
        RECT 25.525 198.755 25.695 198.925 ;
        RECT 26.905 199.435 27.075 199.605 ;
        RECT 27.745 199.435 27.915 199.605 ;
        RECT 23.225 198.075 23.395 198.245 ;
        RECT 26.445 198.415 26.615 198.585 ;
        RECT 28.745 199.095 28.915 199.265 ;
        RECT 31.965 199.435 32.135 199.605 ;
        RECT 25.985 198.075 26.155 198.245 ;
        RECT 27.825 197.735 27.995 197.905 ;
        RECT 32.885 198.755 33.055 198.925 ;
        RECT 48.065 199.435 48.235 199.605 ;
        RECT 49.905 199.435 50.075 199.605 ;
        RECT 47.605 198.755 47.775 198.925 ;
        RECT 48.525 198.755 48.695 198.925 ;
        RECT 48.985 198.755 49.155 198.925 ;
        RECT 49.905 198.755 50.075 198.925 ;
        RECT 54.045 199.435 54.215 199.605 ;
        RECT 52.205 198.755 52.375 198.925 ;
        RECT 51.745 198.415 51.915 198.585 ;
        RECT 69.685 199.435 69.855 199.605 ;
        RECT 71.985 198.755 72.155 198.925 ;
        RECT 76.585 199.095 76.755 199.265 ;
        RECT 71.525 197.735 71.695 197.905 ;
        RECT 77.665 199.095 77.835 199.265 ;
        RECT 79.345 199.095 79.515 199.265 ;
        RECT 78.425 198.075 78.595 198.245 ;
        RECT 80.345 199.435 80.515 199.605 ;
        RECT 81.185 199.435 81.355 199.605 ;
        RECT 77.505 197.735 77.675 197.905 ;
        RECT 84.865 199.435 85.035 199.605 ;
        RECT 83.025 199.095 83.195 199.265 ;
        RECT 83.945 199.095 84.115 199.265 ;
        RECT 80.265 197.735 80.435 197.905 ;
        RECT 92.225 198.755 92.395 198.925 ;
        RECT 92.685 198.415 92.855 198.585 ;
        RECT 98.665 199.095 98.835 199.265 ;
        RECT 94.065 197.735 94.235 197.905 ;
        RECT 100.505 199.435 100.675 199.605 ;
        RECT 99.745 199.095 99.915 199.265 ;
        RECT 99.585 197.735 99.755 197.905 ;
        RECT 100.965 198.755 101.135 198.925 ;
        RECT 105.105 198.415 105.275 198.585 ;
        RECT 105.590 198.075 105.760 198.245 ;
        RECT 105.985 198.415 106.155 198.585 ;
        RECT 106.440 198.755 106.610 198.925 ;
        RECT 107.175 198.415 107.345 198.585 ;
        RECT 107.690 198.075 107.860 198.245 ;
        RECT 109.260 198.075 109.430 198.245 ;
        RECT 109.695 198.415 109.865 198.585 ;
        RECT 114.765 198.755 114.935 198.925 ;
        RECT 115.685 198.755 115.855 198.925 ;
        RECT 116.605 198.755 116.775 198.925 ;
        RECT 112.005 197.735 112.175 197.905 ;
        RECT 117.065 199.435 117.235 199.605 ;
        RECT 117.985 198.755 118.155 198.925 ;
        RECT 123.045 197.735 123.215 197.905 ;
        RECT 125.355 198.415 125.525 198.585 ;
        RECT 125.790 198.075 125.960 198.245 ;
        RECT 127.875 198.415 128.045 198.585 ;
        RECT 127.360 198.075 127.530 198.245 ;
        RECT 128.665 198.755 128.835 198.925 ;
        RECT 129.065 198.415 129.235 198.585 ;
        RECT 129.945 198.755 130.115 198.925 ;
        RECT 129.460 198.075 129.630 198.245 ;
        RECT 11.265 197.225 11.435 197.395 ;
        RECT 11.725 197.225 11.895 197.395 ;
        RECT 12.185 197.225 12.355 197.395 ;
        RECT 12.645 197.225 12.815 197.395 ;
        RECT 13.105 197.225 13.275 197.395 ;
        RECT 13.565 197.225 13.735 197.395 ;
        RECT 14.025 197.225 14.195 197.395 ;
        RECT 14.485 197.225 14.655 197.395 ;
        RECT 14.945 197.225 15.115 197.395 ;
        RECT 15.405 197.225 15.575 197.395 ;
        RECT 15.865 197.225 16.035 197.395 ;
        RECT 16.325 197.225 16.495 197.395 ;
        RECT 16.785 197.225 16.955 197.395 ;
        RECT 17.245 197.225 17.415 197.395 ;
        RECT 17.705 197.225 17.875 197.395 ;
        RECT 18.165 197.225 18.335 197.395 ;
        RECT 18.625 197.225 18.795 197.395 ;
        RECT 19.085 197.225 19.255 197.395 ;
        RECT 19.545 197.225 19.715 197.395 ;
        RECT 20.005 197.225 20.175 197.395 ;
        RECT 20.465 197.225 20.635 197.395 ;
        RECT 20.925 197.225 21.095 197.395 ;
        RECT 21.385 197.225 21.555 197.395 ;
        RECT 21.845 197.225 22.015 197.395 ;
        RECT 22.305 197.225 22.475 197.395 ;
        RECT 22.765 197.225 22.935 197.395 ;
        RECT 23.225 197.225 23.395 197.395 ;
        RECT 23.685 197.225 23.855 197.395 ;
        RECT 24.145 197.225 24.315 197.395 ;
        RECT 24.605 197.225 24.775 197.395 ;
        RECT 25.065 197.225 25.235 197.395 ;
        RECT 25.525 197.225 25.695 197.395 ;
        RECT 25.985 197.225 26.155 197.395 ;
        RECT 26.445 197.225 26.615 197.395 ;
        RECT 26.905 197.225 27.075 197.395 ;
        RECT 27.365 197.225 27.535 197.395 ;
        RECT 27.825 197.225 27.995 197.395 ;
        RECT 28.285 197.225 28.455 197.395 ;
        RECT 28.745 197.225 28.915 197.395 ;
        RECT 29.205 197.225 29.375 197.395 ;
        RECT 29.665 197.225 29.835 197.395 ;
        RECT 30.125 197.225 30.295 197.395 ;
        RECT 30.585 197.225 30.755 197.395 ;
        RECT 31.045 197.225 31.215 197.395 ;
        RECT 31.505 197.225 31.675 197.395 ;
        RECT 31.965 197.225 32.135 197.395 ;
        RECT 32.425 197.225 32.595 197.395 ;
        RECT 32.885 197.225 33.055 197.395 ;
        RECT 33.345 197.225 33.515 197.395 ;
        RECT 33.805 197.225 33.975 197.395 ;
        RECT 34.265 197.225 34.435 197.395 ;
        RECT 34.725 197.225 34.895 197.395 ;
        RECT 35.185 197.225 35.355 197.395 ;
        RECT 35.645 197.225 35.815 197.395 ;
        RECT 36.105 197.225 36.275 197.395 ;
        RECT 36.565 197.225 36.735 197.395 ;
        RECT 37.025 197.225 37.195 197.395 ;
        RECT 37.485 197.225 37.655 197.395 ;
        RECT 37.945 197.225 38.115 197.395 ;
        RECT 38.405 197.225 38.575 197.395 ;
        RECT 38.865 197.225 39.035 197.395 ;
        RECT 39.325 197.225 39.495 197.395 ;
        RECT 39.785 197.225 39.955 197.395 ;
        RECT 40.245 197.225 40.415 197.395 ;
        RECT 40.705 197.225 40.875 197.395 ;
        RECT 41.165 197.225 41.335 197.395 ;
        RECT 41.625 197.225 41.795 197.395 ;
        RECT 42.085 197.225 42.255 197.395 ;
        RECT 42.545 197.225 42.715 197.395 ;
        RECT 43.005 197.225 43.175 197.395 ;
        RECT 43.465 197.225 43.635 197.395 ;
        RECT 43.925 197.225 44.095 197.395 ;
        RECT 44.385 197.225 44.555 197.395 ;
        RECT 44.845 197.225 45.015 197.395 ;
        RECT 45.305 197.225 45.475 197.395 ;
        RECT 45.765 197.225 45.935 197.395 ;
        RECT 46.225 197.225 46.395 197.395 ;
        RECT 46.685 197.225 46.855 197.395 ;
        RECT 47.145 197.225 47.315 197.395 ;
        RECT 47.605 197.225 47.775 197.395 ;
        RECT 48.065 197.225 48.235 197.395 ;
        RECT 48.525 197.225 48.695 197.395 ;
        RECT 48.985 197.225 49.155 197.395 ;
        RECT 49.445 197.225 49.615 197.395 ;
        RECT 49.905 197.225 50.075 197.395 ;
        RECT 50.365 197.225 50.535 197.395 ;
        RECT 50.825 197.225 50.995 197.395 ;
        RECT 51.285 197.225 51.455 197.395 ;
        RECT 51.745 197.225 51.915 197.395 ;
        RECT 52.205 197.225 52.375 197.395 ;
        RECT 52.665 197.225 52.835 197.395 ;
        RECT 53.125 197.225 53.295 197.395 ;
        RECT 53.585 197.225 53.755 197.395 ;
        RECT 54.045 197.225 54.215 197.395 ;
        RECT 54.505 197.225 54.675 197.395 ;
        RECT 54.965 197.225 55.135 197.395 ;
        RECT 55.425 197.225 55.595 197.395 ;
        RECT 55.885 197.225 56.055 197.395 ;
        RECT 56.345 197.225 56.515 197.395 ;
        RECT 56.805 197.225 56.975 197.395 ;
        RECT 57.265 197.225 57.435 197.395 ;
        RECT 57.725 197.225 57.895 197.395 ;
        RECT 58.185 197.225 58.355 197.395 ;
        RECT 58.645 197.225 58.815 197.395 ;
        RECT 59.105 197.225 59.275 197.395 ;
        RECT 59.565 197.225 59.735 197.395 ;
        RECT 60.025 197.225 60.195 197.395 ;
        RECT 60.485 197.225 60.655 197.395 ;
        RECT 60.945 197.225 61.115 197.395 ;
        RECT 61.405 197.225 61.575 197.395 ;
        RECT 61.865 197.225 62.035 197.395 ;
        RECT 62.325 197.225 62.495 197.395 ;
        RECT 62.785 197.225 62.955 197.395 ;
        RECT 63.245 197.225 63.415 197.395 ;
        RECT 63.705 197.225 63.875 197.395 ;
        RECT 64.165 197.225 64.335 197.395 ;
        RECT 64.625 197.225 64.795 197.395 ;
        RECT 65.085 197.225 65.255 197.395 ;
        RECT 65.545 197.225 65.715 197.395 ;
        RECT 66.005 197.225 66.175 197.395 ;
        RECT 66.465 197.225 66.635 197.395 ;
        RECT 66.925 197.225 67.095 197.395 ;
        RECT 67.385 197.225 67.555 197.395 ;
        RECT 67.845 197.225 68.015 197.395 ;
        RECT 68.305 197.225 68.475 197.395 ;
        RECT 68.765 197.225 68.935 197.395 ;
        RECT 69.225 197.225 69.395 197.395 ;
        RECT 69.685 197.225 69.855 197.395 ;
        RECT 70.145 197.225 70.315 197.395 ;
        RECT 70.605 197.225 70.775 197.395 ;
        RECT 71.065 197.225 71.235 197.395 ;
        RECT 71.525 197.225 71.695 197.395 ;
        RECT 71.985 197.225 72.155 197.395 ;
        RECT 72.445 197.225 72.615 197.395 ;
        RECT 72.905 197.225 73.075 197.395 ;
        RECT 73.365 197.225 73.535 197.395 ;
        RECT 73.825 197.225 73.995 197.395 ;
        RECT 74.285 197.225 74.455 197.395 ;
        RECT 74.745 197.225 74.915 197.395 ;
        RECT 75.205 197.225 75.375 197.395 ;
        RECT 75.665 197.225 75.835 197.395 ;
        RECT 76.125 197.225 76.295 197.395 ;
        RECT 76.585 197.225 76.755 197.395 ;
        RECT 77.045 197.225 77.215 197.395 ;
        RECT 77.505 197.225 77.675 197.395 ;
        RECT 77.965 197.225 78.135 197.395 ;
        RECT 78.425 197.225 78.595 197.395 ;
        RECT 78.885 197.225 79.055 197.395 ;
        RECT 79.345 197.225 79.515 197.395 ;
        RECT 79.805 197.225 79.975 197.395 ;
        RECT 80.265 197.225 80.435 197.395 ;
        RECT 80.725 197.225 80.895 197.395 ;
        RECT 81.185 197.225 81.355 197.395 ;
        RECT 81.645 197.225 81.815 197.395 ;
        RECT 82.105 197.225 82.275 197.395 ;
        RECT 82.565 197.225 82.735 197.395 ;
        RECT 83.025 197.225 83.195 197.395 ;
        RECT 83.485 197.225 83.655 197.395 ;
        RECT 83.945 197.225 84.115 197.395 ;
        RECT 84.405 197.225 84.575 197.395 ;
        RECT 84.865 197.225 85.035 197.395 ;
        RECT 85.325 197.225 85.495 197.395 ;
        RECT 85.785 197.225 85.955 197.395 ;
        RECT 86.245 197.225 86.415 197.395 ;
        RECT 86.705 197.225 86.875 197.395 ;
        RECT 87.165 197.225 87.335 197.395 ;
        RECT 87.625 197.225 87.795 197.395 ;
        RECT 88.085 197.225 88.255 197.395 ;
        RECT 88.545 197.225 88.715 197.395 ;
        RECT 89.005 197.225 89.175 197.395 ;
        RECT 89.465 197.225 89.635 197.395 ;
        RECT 89.925 197.225 90.095 197.395 ;
        RECT 90.385 197.225 90.555 197.395 ;
        RECT 90.845 197.225 91.015 197.395 ;
        RECT 91.305 197.225 91.475 197.395 ;
        RECT 91.765 197.225 91.935 197.395 ;
        RECT 92.225 197.225 92.395 197.395 ;
        RECT 92.685 197.225 92.855 197.395 ;
        RECT 93.145 197.225 93.315 197.395 ;
        RECT 93.605 197.225 93.775 197.395 ;
        RECT 94.065 197.225 94.235 197.395 ;
        RECT 94.525 197.225 94.695 197.395 ;
        RECT 94.985 197.225 95.155 197.395 ;
        RECT 95.445 197.225 95.615 197.395 ;
        RECT 95.905 197.225 96.075 197.395 ;
        RECT 96.365 197.225 96.535 197.395 ;
        RECT 96.825 197.225 96.995 197.395 ;
        RECT 97.285 197.225 97.455 197.395 ;
        RECT 97.745 197.225 97.915 197.395 ;
        RECT 98.205 197.225 98.375 197.395 ;
        RECT 98.665 197.225 98.835 197.395 ;
        RECT 99.125 197.225 99.295 197.395 ;
        RECT 99.585 197.225 99.755 197.395 ;
        RECT 100.045 197.225 100.215 197.395 ;
        RECT 100.505 197.225 100.675 197.395 ;
        RECT 100.965 197.225 101.135 197.395 ;
        RECT 101.425 197.225 101.595 197.395 ;
        RECT 101.885 197.225 102.055 197.395 ;
        RECT 102.345 197.225 102.515 197.395 ;
        RECT 102.805 197.225 102.975 197.395 ;
        RECT 103.265 197.225 103.435 197.395 ;
        RECT 103.725 197.225 103.895 197.395 ;
        RECT 104.185 197.225 104.355 197.395 ;
        RECT 104.645 197.225 104.815 197.395 ;
        RECT 105.105 197.225 105.275 197.395 ;
        RECT 105.565 197.225 105.735 197.395 ;
        RECT 106.025 197.225 106.195 197.395 ;
        RECT 106.485 197.225 106.655 197.395 ;
        RECT 106.945 197.225 107.115 197.395 ;
        RECT 107.405 197.225 107.575 197.395 ;
        RECT 107.865 197.225 108.035 197.395 ;
        RECT 108.325 197.225 108.495 197.395 ;
        RECT 108.785 197.225 108.955 197.395 ;
        RECT 109.245 197.225 109.415 197.395 ;
        RECT 109.705 197.225 109.875 197.395 ;
        RECT 110.165 197.225 110.335 197.395 ;
        RECT 110.625 197.225 110.795 197.395 ;
        RECT 111.085 197.225 111.255 197.395 ;
        RECT 111.545 197.225 111.715 197.395 ;
        RECT 112.005 197.225 112.175 197.395 ;
        RECT 112.465 197.225 112.635 197.395 ;
        RECT 112.925 197.225 113.095 197.395 ;
        RECT 113.385 197.225 113.555 197.395 ;
        RECT 113.845 197.225 114.015 197.395 ;
        RECT 114.305 197.225 114.475 197.395 ;
        RECT 114.765 197.225 114.935 197.395 ;
        RECT 115.225 197.225 115.395 197.395 ;
        RECT 115.685 197.225 115.855 197.395 ;
        RECT 116.145 197.225 116.315 197.395 ;
        RECT 116.605 197.225 116.775 197.395 ;
        RECT 117.065 197.225 117.235 197.395 ;
        RECT 117.525 197.225 117.695 197.395 ;
        RECT 117.985 197.225 118.155 197.395 ;
        RECT 118.445 197.225 118.615 197.395 ;
        RECT 118.905 197.225 119.075 197.395 ;
        RECT 119.365 197.225 119.535 197.395 ;
        RECT 119.825 197.225 119.995 197.395 ;
        RECT 120.285 197.225 120.455 197.395 ;
        RECT 120.745 197.225 120.915 197.395 ;
        RECT 121.205 197.225 121.375 197.395 ;
        RECT 121.665 197.225 121.835 197.395 ;
        RECT 122.125 197.225 122.295 197.395 ;
        RECT 122.585 197.225 122.755 197.395 ;
        RECT 123.045 197.225 123.215 197.395 ;
        RECT 123.505 197.225 123.675 197.395 ;
        RECT 123.965 197.225 124.135 197.395 ;
        RECT 124.425 197.225 124.595 197.395 ;
        RECT 124.885 197.225 125.055 197.395 ;
        RECT 125.345 197.225 125.515 197.395 ;
        RECT 125.805 197.225 125.975 197.395 ;
        RECT 126.265 197.225 126.435 197.395 ;
        RECT 126.725 197.225 126.895 197.395 ;
        RECT 127.185 197.225 127.355 197.395 ;
        RECT 127.645 197.225 127.815 197.395 ;
        RECT 128.105 197.225 128.275 197.395 ;
        RECT 128.565 197.225 128.735 197.395 ;
        RECT 129.025 197.225 129.195 197.395 ;
        RECT 129.485 197.225 129.655 197.395 ;
        RECT 129.945 197.225 130.115 197.395 ;
        RECT 130.405 197.225 130.575 197.395 ;
        RECT 130.865 197.225 131.035 197.395 ;
        RECT 131.325 197.225 131.495 197.395 ;
        RECT 131.785 197.225 131.955 197.395 ;
        RECT 132.245 197.225 132.415 197.395 ;
        RECT 132.705 197.225 132.875 197.395 ;
        RECT 133.165 197.225 133.335 197.395 ;
        RECT 133.625 197.225 133.795 197.395 ;
        RECT 134.085 197.225 134.255 197.395 ;
        RECT 134.545 197.225 134.715 197.395 ;
        RECT 135.005 197.225 135.175 197.395 ;
        RECT 135.465 197.225 135.635 197.395 ;
        RECT 135.925 197.225 136.095 197.395 ;
        RECT 136.385 197.225 136.555 197.395 ;
        RECT 136.845 197.225 137.015 197.395 ;
        RECT 137.305 197.225 137.475 197.395 ;
        RECT 137.765 197.225 137.935 197.395 ;
        RECT 138.225 197.225 138.395 197.395 ;
        RECT 138.685 197.225 138.855 197.395 ;
        RECT 139.145 197.225 139.315 197.395 ;
        RECT 139.605 197.225 139.775 197.395 ;
        RECT 140.065 197.225 140.235 197.395 ;
        RECT 140.525 197.225 140.695 197.395 ;
        RECT 140.985 197.225 141.155 197.395 ;
        RECT 141.445 197.225 141.615 197.395 ;
        RECT 141.905 197.225 142.075 197.395 ;
        RECT 142.365 197.225 142.535 197.395 ;
        RECT 142.825 197.225 142.995 197.395 ;
        RECT 143.285 197.225 143.455 197.395 ;
        RECT 143.745 197.225 143.915 197.395 ;
        RECT 144.205 197.225 144.375 197.395 ;
        RECT 144.665 197.225 144.835 197.395 ;
        RECT 145.125 197.225 145.295 197.395 ;
        RECT 145.585 197.225 145.755 197.395 ;
        RECT 146.045 197.225 146.215 197.395 ;
        RECT 146.505 197.225 146.675 197.395 ;
        RECT 146.965 197.225 147.135 197.395 ;
        RECT 147.425 197.225 147.595 197.395 ;
        RECT 147.885 197.225 148.055 197.395 ;
        RECT 148.345 197.225 148.515 197.395 ;
        RECT 148.805 197.225 148.975 197.395 ;
        RECT 149.265 197.225 149.435 197.395 ;
        RECT 149.725 197.225 149.895 197.395 ;
        RECT 150.185 197.225 150.355 197.395 ;
        RECT 39.785 196.375 39.955 196.545 ;
        RECT 41.625 196.715 41.795 196.885 ;
        RECT 44.385 196.715 44.555 196.885 ;
        RECT 41.165 195.695 41.335 195.865 ;
        RECT 43.925 196.035 44.095 196.205 ;
        RECT 44.845 195.695 45.015 195.865 ;
        RECT 45.305 195.695 45.475 195.865 ;
        RECT 57.725 195.695 57.895 195.865 ;
        RECT 59.565 196.715 59.735 196.885 ;
        RECT 59.565 195.355 59.735 195.525 ;
        RECT 61.430 196.375 61.600 196.545 ;
        RECT 60.945 196.035 61.115 196.205 ;
        RECT 60.485 195.015 60.655 195.185 ;
        RECT 61.825 196.035 61.995 196.205 ;
        RECT 62.280 195.355 62.450 195.525 ;
        RECT 63.530 196.375 63.700 196.545 ;
        RECT 63.015 196.035 63.185 196.205 ;
        RECT 65.100 196.375 65.270 196.545 ;
        RECT 65.535 196.035 65.705 196.205 ;
        RECT 71.065 196.715 71.235 196.885 ;
        RECT 70.145 196.035 70.315 196.205 ;
        RECT 67.845 195.015 68.015 195.185 ;
        RECT 72.445 195.695 72.615 195.865 ;
        RECT 77.965 195.695 78.135 195.865 ;
        RECT 78.885 195.355 79.055 195.525 ;
        RECT 80.265 195.695 80.435 195.865 ;
        RECT 81.185 195.355 81.355 195.525 ;
        RECT 82.565 196.375 82.735 196.545 ;
        RECT 84.405 196.715 84.575 196.885 ;
        RECT 79.805 195.015 79.975 195.185 ;
        RECT 82.105 195.015 82.275 195.185 ;
        RECT 84.405 195.015 84.575 195.185 ;
        RECT 85.325 195.015 85.495 195.185 ;
        RECT 89.950 196.375 90.120 196.545 ;
        RECT 88.085 195.695 88.255 195.865 ;
        RECT 89.465 196.035 89.635 196.205 ;
        RECT 89.005 195.015 89.175 195.185 ;
        RECT 90.345 196.035 90.515 196.205 ;
        RECT 90.690 195.355 90.860 195.525 ;
        RECT 92.050 196.375 92.220 196.545 ;
        RECT 91.535 196.035 91.705 196.205 ;
        RECT 93.620 196.375 93.790 196.545 ;
        RECT 94.055 196.035 94.225 196.205 ;
        RECT 102.805 196.715 102.975 196.885 ;
        RECT 96.365 195.015 96.535 195.185 ;
        RECT 101.885 195.355 102.055 195.525 ;
        RECT 102.885 195.015 103.055 195.185 ;
        RECT 103.725 195.015 103.895 195.185 ;
        RECT 106.485 196.715 106.655 196.885 ;
        RECT 105.105 195.355 105.275 195.525 ;
        RECT 106.025 195.355 106.195 195.525 ;
        RECT 107.405 195.695 107.575 195.865 ;
        RECT 112.925 196.035 113.095 196.205 ;
        RECT 104.185 195.015 104.355 195.185 ;
        RECT 113.845 195.015 114.015 195.185 ;
        RECT 114.305 195.355 114.475 195.525 ;
        RECT 116.145 196.715 116.315 196.885 ;
        RECT 120.745 196.715 120.915 196.885 ;
        RECT 120.285 195.695 120.455 195.865 ;
        RECT 121.665 196.035 121.835 196.205 ;
        RECT 121.665 195.015 121.835 195.185 ;
        RECT 11.265 194.505 11.435 194.675 ;
        RECT 11.725 194.505 11.895 194.675 ;
        RECT 12.185 194.505 12.355 194.675 ;
        RECT 12.645 194.505 12.815 194.675 ;
        RECT 13.105 194.505 13.275 194.675 ;
        RECT 13.565 194.505 13.735 194.675 ;
        RECT 14.025 194.505 14.195 194.675 ;
        RECT 14.485 194.505 14.655 194.675 ;
        RECT 14.945 194.505 15.115 194.675 ;
        RECT 15.405 194.505 15.575 194.675 ;
        RECT 15.865 194.505 16.035 194.675 ;
        RECT 16.325 194.505 16.495 194.675 ;
        RECT 16.785 194.505 16.955 194.675 ;
        RECT 17.245 194.505 17.415 194.675 ;
        RECT 17.705 194.505 17.875 194.675 ;
        RECT 18.165 194.505 18.335 194.675 ;
        RECT 18.625 194.505 18.795 194.675 ;
        RECT 19.085 194.505 19.255 194.675 ;
        RECT 19.545 194.505 19.715 194.675 ;
        RECT 20.005 194.505 20.175 194.675 ;
        RECT 20.465 194.505 20.635 194.675 ;
        RECT 20.925 194.505 21.095 194.675 ;
        RECT 21.385 194.505 21.555 194.675 ;
        RECT 21.845 194.505 22.015 194.675 ;
        RECT 22.305 194.505 22.475 194.675 ;
        RECT 22.765 194.505 22.935 194.675 ;
        RECT 23.225 194.505 23.395 194.675 ;
        RECT 23.685 194.505 23.855 194.675 ;
        RECT 24.145 194.505 24.315 194.675 ;
        RECT 24.605 194.505 24.775 194.675 ;
        RECT 25.065 194.505 25.235 194.675 ;
        RECT 25.525 194.505 25.695 194.675 ;
        RECT 25.985 194.505 26.155 194.675 ;
        RECT 26.445 194.505 26.615 194.675 ;
        RECT 26.905 194.505 27.075 194.675 ;
        RECT 27.365 194.505 27.535 194.675 ;
        RECT 27.825 194.505 27.995 194.675 ;
        RECT 28.285 194.505 28.455 194.675 ;
        RECT 28.745 194.505 28.915 194.675 ;
        RECT 29.205 194.505 29.375 194.675 ;
        RECT 29.665 194.505 29.835 194.675 ;
        RECT 30.125 194.505 30.295 194.675 ;
        RECT 30.585 194.505 30.755 194.675 ;
        RECT 31.045 194.505 31.215 194.675 ;
        RECT 31.505 194.505 31.675 194.675 ;
        RECT 31.965 194.505 32.135 194.675 ;
        RECT 32.425 194.505 32.595 194.675 ;
        RECT 32.885 194.505 33.055 194.675 ;
        RECT 33.345 194.505 33.515 194.675 ;
        RECT 33.805 194.505 33.975 194.675 ;
        RECT 34.265 194.505 34.435 194.675 ;
        RECT 34.725 194.505 34.895 194.675 ;
        RECT 35.185 194.505 35.355 194.675 ;
        RECT 35.645 194.505 35.815 194.675 ;
        RECT 36.105 194.505 36.275 194.675 ;
        RECT 36.565 194.505 36.735 194.675 ;
        RECT 37.025 194.505 37.195 194.675 ;
        RECT 37.485 194.505 37.655 194.675 ;
        RECT 37.945 194.505 38.115 194.675 ;
        RECT 38.405 194.505 38.575 194.675 ;
        RECT 38.865 194.505 39.035 194.675 ;
        RECT 39.325 194.505 39.495 194.675 ;
        RECT 39.785 194.505 39.955 194.675 ;
        RECT 40.245 194.505 40.415 194.675 ;
        RECT 40.705 194.505 40.875 194.675 ;
        RECT 41.165 194.505 41.335 194.675 ;
        RECT 41.625 194.505 41.795 194.675 ;
        RECT 42.085 194.505 42.255 194.675 ;
        RECT 42.545 194.505 42.715 194.675 ;
        RECT 43.005 194.505 43.175 194.675 ;
        RECT 43.465 194.505 43.635 194.675 ;
        RECT 43.925 194.505 44.095 194.675 ;
        RECT 44.385 194.505 44.555 194.675 ;
        RECT 44.845 194.505 45.015 194.675 ;
        RECT 45.305 194.505 45.475 194.675 ;
        RECT 45.765 194.505 45.935 194.675 ;
        RECT 46.225 194.505 46.395 194.675 ;
        RECT 46.685 194.505 46.855 194.675 ;
        RECT 47.145 194.505 47.315 194.675 ;
        RECT 47.605 194.505 47.775 194.675 ;
        RECT 48.065 194.505 48.235 194.675 ;
        RECT 48.525 194.505 48.695 194.675 ;
        RECT 48.985 194.505 49.155 194.675 ;
        RECT 49.445 194.505 49.615 194.675 ;
        RECT 49.905 194.505 50.075 194.675 ;
        RECT 50.365 194.505 50.535 194.675 ;
        RECT 50.825 194.505 50.995 194.675 ;
        RECT 51.285 194.505 51.455 194.675 ;
        RECT 51.745 194.505 51.915 194.675 ;
        RECT 52.205 194.505 52.375 194.675 ;
        RECT 52.665 194.505 52.835 194.675 ;
        RECT 53.125 194.505 53.295 194.675 ;
        RECT 53.585 194.505 53.755 194.675 ;
        RECT 54.045 194.505 54.215 194.675 ;
        RECT 54.505 194.505 54.675 194.675 ;
        RECT 54.965 194.505 55.135 194.675 ;
        RECT 55.425 194.505 55.595 194.675 ;
        RECT 55.885 194.505 56.055 194.675 ;
        RECT 56.345 194.505 56.515 194.675 ;
        RECT 56.805 194.505 56.975 194.675 ;
        RECT 57.265 194.505 57.435 194.675 ;
        RECT 57.725 194.505 57.895 194.675 ;
        RECT 58.185 194.505 58.355 194.675 ;
        RECT 58.645 194.505 58.815 194.675 ;
        RECT 59.105 194.505 59.275 194.675 ;
        RECT 59.565 194.505 59.735 194.675 ;
        RECT 60.025 194.505 60.195 194.675 ;
        RECT 60.485 194.505 60.655 194.675 ;
        RECT 60.945 194.505 61.115 194.675 ;
        RECT 61.405 194.505 61.575 194.675 ;
        RECT 61.865 194.505 62.035 194.675 ;
        RECT 62.325 194.505 62.495 194.675 ;
        RECT 62.785 194.505 62.955 194.675 ;
        RECT 63.245 194.505 63.415 194.675 ;
        RECT 63.705 194.505 63.875 194.675 ;
        RECT 64.165 194.505 64.335 194.675 ;
        RECT 64.625 194.505 64.795 194.675 ;
        RECT 65.085 194.505 65.255 194.675 ;
        RECT 65.545 194.505 65.715 194.675 ;
        RECT 66.005 194.505 66.175 194.675 ;
        RECT 66.465 194.505 66.635 194.675 ;
        RECT 66.925 194.505 67.095 194.675 ;
        RECT 67.385 194.505 67.555 194.675 ;
        RECT 67.845 194.505 68.015 194.675 ;
        RECT 68.305 194.505 68.475 194.675 ;
        RECT 68.765 194.505 68.935 194.675 ;
        RECT 69.225 194.505 69.395 194.675 ;
        RECT 69.685 194.505 69.855 194.675 ;
        RECT 70.145 194.505 70.315 194.675 ;
        RECT 70.605 194.505 70.775 194.675 ;
        RECT 71.065 194.505 71.235 194.675 ;
        RECT 71.525 194.505 71.695 194.675 ;
        RECT 71.985 194.505 72.155 194.675 ;
        RECT 72.445 194.505 72.615 194.675 ;
        RECT 72.905 194.505 73.075 194.675 ;
        RECT 73.365 194.505 73.535 194.675 ;
        RECT 73.825 194.505 73.995 194.675 ;
        RECT 74.285 194.505 74.455 194.675 ;
        RECT 74.745 194.505 74.915 194.675 ;
        RECT 75.205 194.505 75.375 194.675 ;
        RECT 75.665 194.505 75.835 194.675 ;
        RECT 76.125 194.505 76.295 194.675 ;
        RECT 76.585 194.505 76.755 194.675 ;
        RECT 77.045 194.505 77.215 194.675 ;
        RECT 77.505 194.505 77.675 194.675 ;
        RECT 77.965 194.505 78.135 194.675 ;
        RECT 78.425 194.505 78.595 194.675 ;
        RECT 78.885 194.505 79.055 194.675 ;
        RECT 79.345 194.505 79.515 194.675 ;
        RECT 79.805 194.505 79.975 194.675 ;
        RECT 80.265 194.505 80.435 194.675 ;
        RECT 80.725 194.505 80.895 194.675 ;
        RECT 81.185 194.505 81.355 194.675 ;
        RECT 81.645 194.505 81.815 194.675 ;
        RECT 82.105 194.505 82.275 194.675 ;
        RECT 82.565 194.505 82.735 194.675 ;
        RECT 83.025 194.505 83.195 194.675 ;
        RECT 83.485 194.505 83.655 194.675 ;
        RECT 83.945 194.505 84.115 194.675 ;
        RECT 84.405 194.505 84.575 194.675 ;
        RECT 84.865 194.505 85.035 194.675 ;
        RECT 85.325 194.505 85.495 194.675 ;
        RECT 85.785 194.505 85.955 194.675 ;
        RECT 86.245 194.505 86.415 194.675 ;
        RECT 86.705 194.505 86.875 194.675 ;
        RECT 87.165 194.505 87.335 194.675 ;
        RECT 87.625 194.505 87.795 194.675 ;
        RECT 88.085 194.505 88.255 194.675 ;
        RECT 88.545 194.505 88.715 194.675 ;
        RECT 89.005 194.505 89.175 194.675 ;
        RECT 89.465 194.505 89.635 194.675 ;
        RECT 89.925 194.505 90.095 194.675 ;
        RECT 90.385 194.505 90.555 194.675 ;
        RECT 90.845 194.505 91.015 194.675 ;
        RECT 91.305 194.505 91.475 194.675 ;
        RECT 91.765 194.505 91.935 194.675 ;
        RECT 92.225 194.505 92.395 194.675 ;
        RECT 92.685 194.505 92.855 194.675 ;
        RECT 93.145 194.505 93.315 194.675 ;
        RECT 93.605 194.505 93.775 194.675 ;
        RECT 94.065 194.505 94.235 194.675 ;
        RECT 94.525 194.505 94.695 194.675 ;
        RECT 94.985 194.505 95.155 194.675 ;
        RECT 95.445 194.505 95.615 194.675 ;
        RECT 95.905 194.505 96.075 194.675 ;
        RECT 96.365 194.505 96.535 194.675 ;
        RECT 96.825 194.505 96.995 194.675 ;
        RECT 97.285 194.505 97.455 194.675 ;
        RECT 97.745 194.505 97.915 194.675 ;
        RECT 98.205 194.505 98.375 194.675 ;
        RECT 98.665 194.505 98.835 194.675 ;
        RECT 99.125 194.505 99.295 194.675 ;
        RECT 99.585 194.505 99.755 194.675 ;
        RECT 100.045 194.505 100.215 194.675 ;
        RECT 100.505 194.505 100.675 194.675 ;
        RECT 100.965 194.505 101.135 194.675 ;
        RECT 101.425 194.505 101.595 194.675 ;
        RECT 101.885 194.505 102.055 194.675 ;
        RECT 102.345 194.505 102.515 194.675 ;
        RECT 102.805 194.505 102.975 194.675 ;
        RECT 103.265 194.505 103.435 194.675 ;
        RECT 103.725 194.505 103.895 194.675 ;
        RECT 104.185 194.505 104.355 194.675 ;
        RECT 104.645 194.505 104.815 194.675 ;
        RECT 105.105 194.505 105.275 194.675 ;
        RECT 105.565 194.505 105.735 194.675 ;
        RECT 106.025 194.505 106.195 194.675 ;
        RECT 106.485 194.505 106.655 194.675 ;
        RECT 106.945 194.505 107.115 194.675 ;
        RECT 107.405 194.505 107.575 194.675 ;
        RECT 107.865 194.505 108.035 194.675 ;
        RECT 108.325 194.505 108.495 194.675 ;
        RECT 108.785 194.505 108.955 194.675 ;
        RECT 109.245 194.505 109.415 194.675 ;
        RECT 109.705 194.505 109.875 194.675 ;
        RECT 110.165 194.505 110.335 194.675 ;
        RECT 110.625 194.505 110.795 194.675 ;
        RECT 111.085 194.505 111.255 194.675 ;
        RECT 111.545 194.505 111.715 194.675 ;
        RECT 112.005 194.505 112.175 194.675 ;
        RECT 112.465 194.505 112.635 194.675 ;
        RECT 112.925 194.505 113.095 194.675 ;
        RECT 113.385 194.505 113.555 194.675 ;
        RECT 113.845 194.505 114.015 194.675 ;
        RECT 114.305 194.505 114.475 194.675 ;
        RECT 114.765 194.505 114.935 194.675 ;
        RECT 115.225 194.505 115.395 194.675 ;
        RECT 115.685 194.505 115.855 194.675 ;
        RECT 116.145 194.505 116.315 194.675 ;
        RECT 116.605 194.505 116.775 194.675 ;
        RECT 117.065 194.505 117.235 194.675 ;
        RECT 117.525 194.505 117.695 194.675 ;
        RECT 117.985 194.505 118.155 194.675 ;
        RECT 118.445 194.505 118.615 194.675 ;
        RECT 118.905 194.505 119.075 194.675 ;
        RECT 119.365 194.505 119.535 194.675 ;
        RECT 119.825 194.505 119.995 194.675 ;
        RECT 120.285 194.505 120.455 194.675 ;
        RECT 120.745 194.505 120.915 194.675 ;
        RECT 121.205 194.505 121.375 194.675 ;
        RECT 121.665 194.505 121.835 194.675 ;
        RECT 122.125 194.505 122.295 194.675 ;
        RECT 122.585 194.505 122.755 194.675 ;
        RECT 123.045 194.505 123.215 194.675 ;
        RECT 123.505 194.505 123.675 194.675 ;
        RECT 123.965 194.505 124.135 194.675 ;
        RECT 124.425 194.505 124.595 194.675 ;
        RECT 124.885 194.505 125.055 194.675 ;
        RECT 125.345 194.505 125.515 194.675 ;
        RECT 125.805 194.505 125.975 194.675 ;
        RECT 126.265 194.505 126.435 194.675 ;
        RECT 126.725 194.505 126.895 194.675 ;
        RECT 127.185 194.505 127.355 194.675 ;
        RECT 127.645 194.505 127.815 194.675 ;
        RECT 128.105 194.505 128.275 194.675 ;
        RECT 128.565 194.505 128.735 194.675 ;
        RECT 129.025 194.505 129.195 194.675 ;
        RECT 129.485 194.505 129.655 194.675 ;
        RECT 129.945 194.505 130.115 194.675 ;
        RECT 130.405 194.505 130.575 194.675 ;
        RECT 130.865 194.505 131.035 194.675 ;
        RECT 131.325 194.505 131.495 194.675 ;
        RECT 131.785 194.505 131.955 194.675 ;
        RECT 132.245 194.505 132.415 194.675 ;
        RECT 132.705 194.505 132.875 194.675 ;
        RECT 133.165 194.505 133.335 194.675 ;
        RECT 133.625 194.505 133.795 194.675 ;
        RECT 134.085 194.505 134.255 194.675 ;
        RECT 134.545 194.505 134.715 194.675 ;
        RECT 135.005 194.505 135.175 194.675 ;
        RECT 135.465 194.505 135.635 194.675 ;
        RECT 135.925 194.505 136.095 194.675 ;
        RECT 136.385 194.505 136.555 194.675 ;
        RECT 136.845 194.505 137.015 194.675 ;
        RECT 137.305 194.505 137.475 194.675 ;
        RECT 137.765 194.505 137.935 194.675 ;
        RECT 138.225 194.505 138.395 194.675 ;
        RECT 138.685 194.505 138.855 194.675 ;
        RECT 139.145 194.505 139.315 194.675 ;
        RECT 139.605 194.505 139.775 194.675 ;
        RECT 140.065 194.505 140.235 194.675 ;
        RECT 140.525 194.505 140.695 194.675 ;
        RECT 140.985 194.505 141.155 194.675 ;
        RECT 141.445 194.505 141.615 194.675 ;
        RECT 141.905 194.505 142.075 194.675 ;
        RECT 142.365 194.505 142.535 194.675 ;
        RECT 142.825 194.505 142.995 194.675 ;
        RECT 143.285 194.505 143.455 194.675 ;
        RECT 143.745 194.505 143.915 194.675 ;
        RECT 144.205 194.505 144.375 194.675 ;
        RECT 144.665 194.505 144.835 194.675 ;
        RECT 145.125 194.505 145.295 194.675 ;
        RECT 145.585 194.505 145.755 194.675 ;
        RECT 146.045 194.505 146.215 194.675 ;
        RECT 146.505 194.505 146.675 194.675 ;
        RECT 146.965 194.505 147.135 194.675 ;
        RECT 147.425 194.505 147.595 194.675 ;
        RECT 147.885 194.505 148.055 194.675 ;
        RECT 148.345 194.505 148.515 194.675 ;
        RECT 148.805 194.505 148.975 194.675 ;
        RECT 149.265 194.505 149.435 194.675 ;
        RECT 149.725 194.505 149.895 194.675 ;
        RECT 150.185 194.505 150.355 194.675 ;
        RECT 14.945 193.315 15.115 193.485 ;
        RECT 15.865 192.975 16.035 193.145 ;
        RECT 14.025 192.295 14.195 192.465 ;
        RECT 16.350 192.635 16.520 192.805 ;
        RECT 16.745 192.975 16.915 193.145 ;
        RECT 17.200 193.315 17.370 193.485 ;
        RECT 17.935 192.975 18.105 193.145 ;
        RECT 18.450 192.635 18.620 192.805 ;
        RECT 20.020 192.635 20.190 192.805 ;
        RECT 20.455 192.975 20.625 193.145 ;
        RECT 23.225 193.315 23.395 193.485 ;
        RECT 22.765 192.295 22.935 192.465 ;
        RECT 23.710 192.635 23.880 192.805 ;
        RECT 24.105 192.975 24.275 193.145 ;
        RECT 24.560 193.315 24.730 193.485 ;
        RECT 25.295 192.975 25.465 193.145 ;
        RECT 25.810 192.635 25.980 192.805 ;
        RECT 27.380 192.635 27.550 192.805 ;
        RECT 27.815 192.975 27.985 193.145 ;
        RECT 30.125 193.995 30.295 194.165 ;
        RECT 31.505 193.315 31.675 193.485 ;
        RECT 31.965 193.315 32.135 193.485 ;
        RECT 32.425 193.995 32.595 194.165 ;
        RECT 34.265 193.315 34.435 193.485 ;
        RECT 30.585 192.635 30.755 192.805 ;
        RECT 33.345 192.295 33.515 192.465 ;
        RECT 35.185 192.295 35.355 192.465 ;
        RECT 37.485 192.295 37.655 192.465 ;
        RECT 38.405 192.975 38.575 193.145 ;
        RECT 38.865 192.975 39.035 193.145 ;
        RECT 39.325 193.315 39.495 193.485 ;
        RECT 39.785 192.975 39.955 193.145 ;
        RECT 41.625 192.635 41.795 192.805 ;
        RECT 40.705 192.295 40.875 192.465 ;
        RECT 43.005 193.655 43.175 193.825 ;
        RECT 44.845 193.315 45.015 193.485 ;
        RECT 44.385 192.975 44.555 193.145 ;
        RECT 46.685 192.975 46.855 193.145 ;
        RECT 49.905 193.995 50.075 194.165 ;
        RECT 48.065 193.315 48.235 193.485 ;
        RECT 47.605 192.975 47.775 193.145 ;
        RECT 57.135 193.995 57.305 194.165 ;
        RECT 55.885 193.315 56.055 193.485 ;
        RECT 53.585 192.295 53.755 192.465 ;
        RECT 55.425 192.295 55.595 192.465 ;
        RECT 58.185 193.655 58.355 193.825 ;
        RECT 61.865 193.995 62.035 194.165 ;
        RECT 56.345 192.635 56.515 192.805 ;
        RECT 60.945 193.315 61.115 193.485 ;
        RECT 57.265 192.295 57.435 192.465 ;
        RECT 63.245 193.995 63.415 194.165 ;
        RECT 64.165 192.975 64.335 193.145 ;
        RECT 64.630 193.315 64.800 193.485 ;
        RECT 65.085 192.975 65.255 193.145 ;
        RECT 65.545 192.975 65.715 193.145 ;
        RECT 66.465 193.315 66.635 193.485 ;
        RECT 67.385 193.315 67.555 193.485 ;
        RECT 70.605 193.315 70.775 193.485 ;
        RECT 71.065 193.315 71.235 193.485 ;
        RECT 78.885 193.995 79.055 194.165 ;
        RECT 67.385 192.295 67.555 192.465 ;
        RECT 77.965 193.315 78.135 193.485 ;
        RECT 77.045 192.975 77.215 193.145 ;
        RECT 79.805 193.315 79.975 193.485 ;
        RECT 81.645 193.995 81.815 194.165 ;
        RECT 85.325 193.995 85.495 194.165 ;
        RECT 84.405 193.315 84.575 193.485 ;
        RECT 82.565 192.635 82.735 192.805 ;
        RECT 81.645 192.295 81.815 192.465 ;
        RECT 89.005 193.315 89.175 193.485 ;
        RECT 89.490 192.635 89.660 192.805 ;
        RECT 89.885 192.975 90.055 193.145 ;
        RECT 90.230 193.655 90.400 193.825 ;
        RECT 91.075 192.975 91.245 193.145 ;
        RECT 91.590 192.635 91.760 192.805 ;
        RECT 93.160 192.635 93.330 192.805 ;
        RECT 93.595 192.975 93.765 193.145 ;
        RECT 98.205 193.315 98.375 193.485 ;
        RECT 102.345 193.995 102.515 194.165 ;
        RECT 99.125 193.315 99.295 193.485 ;
        RECT 99.585 193.315 99.755 193.485 ;
        RECT 100.965 193.315 101.135 193.485 ;
        RECT 95.905 192.295 96.075 192.465 ;
        RECT 100.045 192.295 100.215 192.465 ;
        RECT 108.325 193.995 108.495 194.165 ;
        RECT 105.565 192.975 105.735 193.145 ;
        RECT 105.105 192.635 105.275 192.805 ;
        RECT 110.625 193.995 110.795 194.165 ;
        RECT 111.085 192.975 111.255 193.145 ;
        RECT 118.445 193.315 118.615 193.485 ;
        RECT 118.905 193.315 119.075 193.485 ;
        RECT 119.825 193.315 119.995 193.485 ;
        RECT 121.205 193.315 121.375 193.485 ;
        RECT 123.965 193.315 124.135 193.485 ;
        RECT 120.745 192.295 120.915 192.465 ;
        RECT 121.205 192.295 121.375 192.465 ;
        RECT 123.045 192.635 123.215 192.805 ;
        RECT 124.885 193.315 125.055 193.485 ;
        RECT 125.345 193.315 125.515 193.485 ;
        RECT 126.265 193.315 126.435 193.485 ;
        RECT 124.425 192.295 124.595 192.465 ;
        RECT 127.645 192.975 127.815 193.145 ;
        RECT 127.185 192.295 127.355 192.465 ;
        RECT 128.130 192.635 128.300 192.805 ;
        RECT 128.525 192.975 128.695 193.145 ;
        RECT 128.980 193.315 129.150 193.485 ;
        RECT 129.715 192.975 129.885 193.145 ;
        RECT 130.230 192.635 130.400 192.805 ;
        RECT 131.800 192.635 131.970 192.805 ;
        RECT 132.235 192.975 132.405 193.145 ;
        RECT 134.545 192.295 134.715 192.465 ;
        RECT 11.265 191.785 11.435 191.955 ;
        RECT 11.725 191.785 11.895 191.955 ;
        RECT 12.185 191.785 12.355 191.955 ;
        RECT 12.645 191.785 12.815 191.955 ;
        RECT 13.105 191.785 13.275 191.955 ;
        RECT 13.565 191.785 13.735 191.955 ;
        RECT 14.025 191.785 14.195 191.955 ;
        RECT 14.485 191.785 14.655 191.955 ;
        RECT 14.945 191.785 15.115 191.955 ;
        RECT 15.405 191.785 15.575 191.955 ;
        RECT 15.865 191.785 16.035 191.955 ;
        RECT 16.325 191.785 16.495 191.955 ;
        RECT 16.785 191.785 16.955 191.955 ;
        RECT 17.245 191.785 17.415 191.955 ;
        RECT 17.705 191.785 17.875 191.955 ;
        RECT 18.165 191.785 18.335 191.955 ;
        RECT 18.625 191.785 18.795 191.955 ;
        RECT 19.085 191.785 19.255 191.955 ;
        RECT 19.545 191.785 19.715 191.955 ;
        RECT 20.005 191.785 20.175 191.955 ;
        RECT 20.465 191.785 20.635 191.955 ;
        RECT 20.925 191.785 21.095 191.955 ;
        RECT 21.385 191.785 21.555 191.955 ;
        RECT 21.845 191.785 22.015 191.955 ;
        RECT 22.305 191.785 22.475 191.955 ;
        RECT 22.765 191.785 22.935 191.955 ;
        RECT 23.225 191.785 23.395 191.955 ;
        RECT 23.685 191.785 23.855 191.955 ;
        RECT 24.145 191.785 24.315 191.955 ;
        RECT 24.605 191.785 24.775 191.955 ;
        RECT 25.065 191.785 25.235 191.955 ;
        RECT 25.525 191.785 25.695 191.955 ;
        RECT 25.985 191.785 26.155 191.955 ;
        RECT 26.445 191.785 26.615 191.955 ;
        RECT 26.905 191.785 27.075 191.955 ;
        RECT 27.365 191.785 27.535 191.955 ;
        RECT 27.825 191.785 27.995 191.955 ;
        RECT 28.285 191.785 28.455 191.955 ;
        RECT 28.745 191.785 28.915 191.955 ;
        RECT 29.205 191.785 29.375 191.955 ;
        RECT 29.665 191.785 29.835 191.955 ;
        RECT 30.125 191.785 30.295 191.955 ;
        RECT 30.585 191.785 30.755 191.955 ;
        RECT 31.045 191.785 31.215 191.955 ;
        RECT 31.505 191.785 31.675 191.955 ;
        RECT 31.965 191.785 32.135 191.955 ;
        RECT 32.425 191.785 32.595 191.955 ;
        RECT 32.885 191.785 33.055 191.955 ;
        RECT 33.345 191.785 33.515 191.955 ;
        RECT 33.805 191.785 33.975 191.955 ;
        RECT 34.265 191.785 34.435 191.955 ;
        RECT 34.725 191.785 34.895 191.955 ;
        RECT 35.185 191.785 35.355 191.955 ;
        RECT 35.645 191.785 35.815 191.955 ;
        RECT 36.105 191.785 36.275 191.955 ;
        RECT 36.565 191.785 36.735 191.955 ;
        RECT 37.025 191.785 37.195 191.955 ;
        RECT 37.485 191.785 37.655 191.955 ;
        RECT 37.945 191.785 38.115 191.955 ;
        RECT 38.405 191.785 38.575 191.955 ;
        RECT 38.865 191.785 39.035 191.955 ;
        RECT 39.325 191.785 39.495 191.955 ;
        RECT 39.785 191.785 39.955 191.955 ;
        RECT 40.245 191.785 40.415 191.955 ;
        RECT 40.705 191.785 40.875 191.955 ;
        RECT 41.165 191.785 41.335 191.955 ;
        RECT 41.625 191.785 41.795 191.955 ;
        RECT 42.085 191.785 42.255 191.955 ;
        RECT 42.545 191.785 42.715 191.955 ;
        RECT 43.005 191.785 43.175 191.955 ;
        RECT 43.465 191.785 43.635 191.955 ;
        RECT 43.925 191.785 44.095 191.955 ;
        RECT 44.385 191.785 44.555 191.955 ;
        RECT 44.845 191.785 45.015 191.955 ;
        RECT 45.305 191.785 45.475 191.955 ;
        RECT 45.765 191.785 45.935 191.955 ;
        RECT 46.225 191.785 46.395 191.955 ;
        RECT 46.685 191.785 46.855 191.955 ;
        RECT 47.145 191.785 47.315 191.955 ;
        RECT 47.605 191.785 47.775 191.955 ;
        RECT 48.065 191.785 48.235 191.955 ;
        RECT 48.525 191.785 48.695 191.955 ;
        RECT 48.985 191.785 49.155 191.955 ;
        RECT 49.445 191.785 49.615 191.955 ;
        RECT 49.905 191.785 50.075 191.955 ;
        RECT 50.365 191.785 50.535 191.955 ;
        RECT 50.825 191.785 50.995 191.955 ;
        RECT 51.285 191.785 51.455 191.955 ;
        RECT 51.745 191.785 51.915 191.955 ;
        RECT 52.205 191.785 52.375 191.955 ;
        RECT 52.665 191.785 52.835 191.955 ;
        RECT 53.125 191.785 53.295 191.955 ;
        RECT 53.585 191.785 53.755 191.955 ;
        RECT 54.045 191.785 54.215 191.955 ;
        RECT 54.505 191.785 54.675 191.955 ;
        RECT 54.965 191.785 55.135 191.955 ;
        RECT 55.425 191.785 55.595 191.955 ;
        RECT 55.885 191.785 56.055 191.955 ;
        RECT 56.345 191.785 56.515 191.955 ;
        RECT 56.805 191.785 56.975 191.955 ;
        RECT 57.265 191.785 57.435 191.955 ;
        RECT 57.725 191.785 57.895 191.955 ;
        RECT 58.185 191.785 58.355 191.955 ;
        RECT 58.645 191.785 58.815 191.955 ;
        RECT 59.105 191.785 59.275 191.955 ;
        RECT 59.565 191.785 59.735 191.955 ;
        RECT 60.025 191.785 60.195 191.955 ;
        RECT 60.485 191.785 60.655 191.955 ;
        RECT 60.945 191.785 61.115 191.955 ;
        RECT 61.405 191.785 61.575 191.955 ;
        RECT 61.865 191.785 62.035 191.955 ;
        RECT 62.325 191.785 62.495 191.955 ;
        RECT 62.785 191.785 62.955 191.955 ;
        RECT 63.245 191.785 63.415 191.955 ;
        RECT 63.705 191.785 63.875 191.955 ;
        RECT 64.165 191.785 64.335 191.955 ;
        RECT 64.625 191.785 64.795 191.955 ;
        RECT 65.085 191.785 65.255 191.955 ;
        RECT 65.545 191.785 65.715 191.955 ;
        RECT 66.005 191.785 66.175 191.955 ;
        RECT 66.465 191.785 66.635 191.955 ;
        RECT 66.925 191.785 67.095 191.955 ;
        RECT 67.385 191.785 67.555 191.955 ;
        RECT 67.845 191.785 68.015 191.955 ;
        RECT 68.305 191.785 68.475 191.955 ;
        RECT 68.765 191.785 68.935 191.955 ;
        RECT 69.225 191.785 69.395 191.955 ;
        RECT 69.685 191.785 69.855 191.955 ;
        RECT 70.145 191.785 70.315 191.955 ;
        RECT 70.605 191.785 70.775 191.955 ;
        RECT 71.065 191.785 71.235 191.955 ;
        RECT 71.525 191.785 71.695 191.955 ;
        RECT 71.985 191.785 72.155 191.955 ;
        RECT 72.445 191.785 72.615 191.955 ;
        RECT 72.905 191.785 73.075 191.955 ;
        RECT 73.365 191.785 73.535 191.955 ;
        RECT 73.825 191.785 73.995 191.955 ;
        RECT 74.285 191.785 74.455 191.955 ;
        RECT 74.745 191.785 74.915 191.955 ;
        RECT 75.205 191.785 75.375 191.955 ;
        RECT 75.665 191.785 75.835 191.955 ;
        RECT 76.125 191.785 76.295 191.955 ;
        RECT 76.585 191.785 76.755 191.955 ;
        RECT 77.045 191.785 77.215 191.955 ;
        RECT 77.505 191.785 77.675 191.955 ;
        RECT 77.965 191.785 78.135 191.955 ;
        RECT 78.425 191.785 78.595 191.955 ;
        RECT 78.885 191.785 79.055 191.955 ;
        RECT 79.345 191.785 79.515 191.955 ;
        RECT 79.805 191.785 79.975 191.955 ;
        RECT 80.265 191.785 80.435 191.955 ;
        RECT 80.725 191.785 80.895 191.955 ;
        RECT 81.185 191.785 81.355 191.955 ;
        RECT 81.645 191.785 81.815 191.955 ;
        RECT 82.105 191.785 82.275 191.955 ;
        RECT 82.565 191.785 82.735 191.955 ;
        RECT 83.025 191.785 83.195 191.955 ;
        RECT 83.485 191.785 83.655 191.955 ;
        RECT 83.945 191.785 84.115 191.955 ;
        RECT 84.405 191.785 84.575 191.955 ;
        RECT 84.865 191.785 85.035 191.955 ;
        RECT 85.325 191.785 85.495 191.955 ;
        RECT 85.785 191.785 85.955 191.955 ;
        RECT 86.245 191.785 86.415 191.955 ;
        RECT 86.705 191.785 86.875 191.955 ;
        RECT 87.165 191.785 87.335 191.955 ;
        RECT 87.625 191.785 87.795 191.955 ;
        RECT 88.085 191.785 88.255 191.955 ;
        RECT 88.545 191.785 88.715 191.955 ;
        RECT 89.005 191.785 89.175 191.955 ;
        RECT 89.465 191.785 89.635 191.955 ;
        RECT 89.925 191.785 90.095 191.955 ;
        RECT 90.385 191.785 90.555 191.955 ;
        RECT 90.845 191.785 91.015 191.955 ;
        RECT 91.305 191.785 91.475 191.955 ;
        RECT 91.765 191.785 91.935 191.955 ;
        RECT 92.225 191.785 92.395 191.955 ;
        RECT 92.685 191.785 92.855 191.955 ;
        RECT 93.145 191.785 93.315 191.955 ;
        RECT 93.605 191.785 93.775 191.955 ;
        RECT 94.065 191.785 94.235 191.955 ;
        RECT 94.525 191.785 94.695 191.955 ;
        RECT 94.985 191.785 95.155 191.955 ;
        RECT 95.445 191.785 95.615 191.955 ;
        RECT 95.905 191.785 96.075 191.955 ;
        RECT 96.365 191.785 96.535 191.955 ;
        RECT 96.825 191.785 96.995 191.955 ;
        RECT 97.285 191.785 97.455 191.955 ;
        RECT 97.745 191.785 97.915 191.955 ;
        RECT 98.205 191.785 98.375 191.955 ;
        RECT 98.665 191.785 98.835 191.955 ;
        RECT 99.125 191.785 99.295 191.955 ;
        RECT 99.585 191.785 99.755 191.955 ;
        RECT 100.045 191.785 100.215 191.955 ;
        RECT 100.505 191.785 100.675 191.955 ;
        RECT 100.965 191.785 101.135 191.955 ;
        RECT 101.425 191.785 101.595 191.955 ;
        RECT 101.885 191.785 102.055 191.955 ;
        RECT 102.345 191.785 102.515 191.955 ;
        RECT 102.805 191.785 102.975 191.955 ;
        RECT 103.265 191.785 103.435 191.955 ;
        RECT 103.725 191.785 103.895 191.955 ;
        RECT 104.185 191.785 104.355 191.955 ;
        RECT 104.645 191.785 104.815 191.955 ;
        RECT 105.105 191.785 105.275 191.955 ;
        RECT 105.565 191.785 105.735 191.955 ;
        RECT 106.025 191.785 106.195 191.955 ;
        RECT 106.485 191.785 106.655 191.955 ;
        RECT 106.945 191.785 107.115 191.955 ;
        RECT 107.405 191.785 107.575 191.955 ;
        RECT 107.865 191.785 108.035 191.955 ;
        RECT 108.325 191.785 108.495 191.955 ;
        RECT 108.785 191.785 108.955 191.955 ;
        RECT 109.245 191.785 109.415 191.955 ;
        RECT 109.705 191.785 109.875 191.955 ;
        RECT 110.165 191.785 110.335 191.955 ;
        RECT 110.625 191.785 110.795 191.955 ;
        RECT 111.085 191.785 111.255 191.955 ;
        RECT 111.545 191.785 111.715 191.955 ;
        RECT 112.005 191.785 112.175 191.955 ;
        RECT 112.465 191.785 112.635 191.955 ;
        RECT 112.925 191.785 113.095 191.955 ;
        RECT 113.385 191.785 113.555 191.955 ;
        RECT 113.845 191.785 114.015 191.955 ;
        RECT 114.305 191.785 114.475 191.955 ;
        RECT 114.765 191.785 114.935 191.955 ;
        RECT 115.225 191.785 115.395 191.955 ;
        RECT 115.685 191.785 115.855 191.955 ;
        RECT 116.145 191.785 116.315 191.955 ;
        RECT 116.605 191.785 116.775 191.955 ;
        RECT 117.065 191.785 117.235 191.955 ;
        RECT 117.525 191.785 117.695 191.955 ;
        RECT 117.985 191.785 118.155 191.955 ;
        RECT 118.445 191.785 118.615 191.955 ;
        RECT 118.905 191.785 119.075 191.955 ;
        RECT 119.365 191.785 119.535 191.955 ;
        RECT 119.825 191.785 119.995 191.955 ;
        RECT 120.285 191.785 120.455 191.955 ;
        RECT 120.745 191.785 120.915 191.955 ;
        RECT 121.205 191.785 121.375 191.955 ;
        RECT 121.665 191.785 121.835 191.955 ;
        RECT 122.125 191.785 122.295 191.955 ;
        RECT 122.585 191.785 122.755 191.955 ;
        RECT 123.045 191.785 123.215 191.955 ;
        RECT 123.505 191.785 123.675 191.955 ;
        RECT 123.965 191.785 124.135 191.955 ;
        RECT 124.425 191.785 124.595 191.955 ;
        RECT 124.885 191.785 125.055 191.955 ;
        RECT 125.345 191.785 125.515 191.955 ;
        RECT 125.805 191.785 125.975 191.955 ;
        RECT 126.265 191.785 126.435 191.955 ;
        RECT 126.725 191.785 126.895 191.955 ;
        RECT 127.185 191.785 127.355 191.955 ;
        RECT 127.645 191.785 127.815 191.955 ;
        RECT 128.105 191.785 128.275 191.955 ;
        RECT 128.565 191.785 128.735 191.955 ;
        RECT 129.025 191.785 129.195 191.955 ;
        RECT 129.485 191.785 129.655 191.955 ;
        RECT 129.945 191.785 130.115 191.955 ;
        RECT 130.405 191.785 130.575 191.955 ;
        RECT 130.865 191.785 131.035 191.955 ;
        RECT 131.325 191.785 131.495 191.955 ;
        RECT 131.785 191.785 131.955 191.955 ;
        RECT 132.245 191.785 132.415 191.955 ;
        RECT 132.705 191.785 132.875 191.955 ;
        RECT 133.165 191.785 133.335 191.955 ;
        RECT 133.625 191.785 133.795 191.955 ;
        RECT 134.085 191.785 134.255 191.955 ;
        RECT 134.545 191.785 134.715 191.955 ;
        RECT 135.005 191.785 135.175 191.955 ;
        RECT 135.465 191.785 135.635 191.955 ;
        RECT 135.925 191.785 136.095 191.955 ;
        RECT 136.385 191.785 136.555 191.955 ;
        RECT 136.845 191.785 137.015 191.955 ;
        RECT 137.305 191.785 137.475 191.955 ;
        RECT 137.765 191.785 137.935 191.955 ;
        RECT 138.225 191.785 138.395 191.955 ;
        RECT 138.685 191.785 138.855 191.955 ;
        RECT 139.145 191.785 139.315 191.955 ;
        RECT 139.605 191.785 139.775 191.955 ;
        RECT 140.065 191.785 140.235 191.955 ;
        RECT 140.525 191.785 140.695 191.955 ;
        RECT 140.985 191.785 141.155 191.955 ;
        RECT 141.445 191.785 141.615 191.955 ;
        RECT 141.905 191.785 142.075 191.955 ;
        RECT 142.365 191.785 142.535 191.955 ;
        RECT 142.825 191.785 142.995 191.955 ;
        RECT 143.285 191.785 143.455 191.955 ;
        RECT 143.745 191.785 143.915 191.955 ;
        RECT 144.205 191.785 144.375 191.955 ;
        RECT 144.665 191.785 144.835 191.955 ;
        RECT 145.125 191.785 145.295 191.955 ;
        RECT 145.585 191.785 145.755 191.955 ;
        RECT 146.045 191.785 146.215 191.955 ;
        RECT 146.505 191.785 146.675 191.955 ;
        RECT 146.965 191.785 147.135 191.955 ;
        RECT 147.425 191.785 147.595 191.955 ;
        RECT 147.885 191.785 148.055 191.955 ;
        RECT 148.345 191.785 148.515 191.955 ;
        RECT 148.805 191.785 148.975 191.955 ;
        RECT 149.265 191.785 149.435 191.955 ;
        RECT 149.725 191.785 149.895 191.955 ;
        RECT 150.185 191.785 150.355 191.955 ;
        RECT 13.130 190.935 13.300 191.105 ;
        RECT 12.645 190.255 12.815 190.425 ;
        RECT 13.525 190.595 13.695 190.765 ;
        RECT 13.980 189.915 14.150 190.085 ;
        RECT 15.230 190.935 15.400 191.105 ;
        RECT 14.715 190.595 14.885 190.765 ;
        RECT 16.800 190.935 16.970 191.105 ;
        RECT 17.235 190.595 17.405 190.765 ;
        RECT 19.545 190.935 19.715 191.105 ;
        RECT 21.845 191.275 22.015 191.445 ;
        RECT 21.385 190.255 21.555 190.425 ;
        RECT 20.465 189.575 20.635 189.745 ;
        RECT 22.765 190.255 22.935 190.425 ;
        RECT 29.665 191.275 29.835 191.445 ;
        RECT 28.745 190.255 28.915 190.425 ;
        RECT 29.205 190.255 29.375 190.425 ;
        RECT 27.825 189.575 27.995 189.745 ;
        RECT 31.505 189.575 31.675 189.745 ;
        RECT 32.425 191.275 32.595 191.445 ;
        RECT 33.345 191.275 33.515 191.445 ;
        RECT 33.345 189.575 33.515 189.745 ;
        RECT 35.185 190.255 35.355 190.425 ;
        RECT 40.705 191.275 40.875 191.445 ;
        RECT 39.325 190.255 39.495 190.425 ;
        RECT 39.785 189.915 39.955 190.085 ;
        RECT 40.705 190.255 40.875 190.425 ;
        RECT 54.045 190.255 54.215 190.425 ;
        RECT 54.965 190.255 55.135 190.425 ;
        RECT 55.425 190.255 55.595 190.425 ;
        RECT 53.125 189.575 53.295 189.745 ;
        RECT 70.145 190.255 70.315 190.425 ;
        RECT 71.105 190.265 71.275 190.435 ;
        RECT 56.345 189.575 56.515 189.745 ;
        RECT 71.065 189.575 71.235 189.745 ;
        RECT 78.425 190.255 78.595 190.425 ;
        RECT 89.005 191.275 89.175 191.445 ;
        RECT 79.345 189.575 79.515 189.745 ;
        RECT 95.905 190.255 96.075 190.425 ;
        RECT 96.370 190.255 96.540 190.425 ;
        RECT 97.285 190.255 97.455 190.425 ;
        RECT 95.445 189.915 95.615 190.085 ;
        RECT 98.435 190.255 98.605 190.425 ;
        RECT 97.745 189.915 97.915 190.085 ;
        RECT 99.125 189.575 99.295 189.745 ;
        RECT 108.325 191.275 108.495 191.445 ;
        RECT 111.085 191.275 111.255 191.445 ;
        RECT 101.885 189.915 102.055 190.085 ;
        RECT 112.465 190.595 112.635 190.765 ;
        RECT 112.925 190.255 113.095 190.425 ;
        RECT 116.605 190.595 116.775 190.765 ;
        RECT 117.525 190.255 117.695 190.425 ;
        RECT 119.365 190.255 119.535 190.425 ;
        RECT 120.285 190.255 120.455 190.425 ;
        RECT 121.205 190.255 121.375 190.425 ;
        RECT 120.745 189.575 120.915 189.745 ;
        RECT 122.125 189.915 122.295 190.085 ;
        RECT 123.045 190.255 123.215 190.425 ;
        RECT 122.585 189.915 122.755 190.085 ;
        RECT 123.965 189.575 124.135 189.745 ;
        RECT 127.645 191.275 127.815 191.445 ;
        RECT 130.865 191.275 131.035 191.445 ;
        RECT 128.565 190.255 128.735 190.425 ;
        RECT 129.025 190.255 129.195 190.425 ;
        RECT 130.405 190.255 130.575 190.425 ;
        RECT 129.485 189.915 129.655 190.085 ;
        RECT 131.785 190.255 131.955 190.425 ;
        RECT 11.265 189.065 11.435 189.235 ;
        RECT 11.725 189.065 11.895 189.235 ;
        RECT 12.185 189.065 12.355 189.235 ;
        RECT 12.645 189.065 12.815 189.235 ;
        RECT 13.105 189.065 13.275 189.235 ;
        RECT 13.565 189.065 13.735 189.235 ;
        RECT 14.025 189.065 14.195 189.235 ;
        RECT 14.485 189.065 14.655 189.235 ;
        RECT 14.945 189.065 15.115 189.235 ;
        RECT 15.405 189.065 15.575 189.235 ;
        RECT 15.865 189.065 16.035 189.235 ;
        RECT 16.325 189.065 16.495 189.235 ;
        RECT 16.785 189.065 16.955 189.235 ;
        RECT 17.245 189.065 17.415 189.235 ;
        RECT 17.705 189.065 17.875 189.235 ;
        RECT 18.165 189.065 18.335 189.235 ;
        RECT 18.625 189.065 18.795 189.235 ;
        RECT 19.085 189.065 19.255 189.235 ;
        RECT 19.545 189.065 19.715 189.235 ;
        RECT 20.005 189.065 20.175 189.235 ;
        RECT 20.465 189.065 20.635 189.235 ;
        RECT 20.925 189.065 21.095 189.235 ;
        RECT 21.385 189.065 21.555 189.235 ;
        RECT 21.845 189.065 22.015 189.235 ;
        RECT 22.305 189.065 22.475 189.235 ;
        RECT 22.765 189.065 22.935 189.235 ;
        RECT 23.225 189.065 23.395 189.235 ;
        RECT 23.685 189.065 23.855 189.235 ;
        RECT 24.145 189.065 24.315 189.235 ;
        RECT 24.605 189.065 24.775 189.235 ;
        RECT 25.065 189.065 25.235 189.235 ;
        RECT 25.525 189.065 25.695 189.235 ;
        RECT 25.985 189.065 26.155 189.235 ;
        RECT 26.445 189.065 26.615 189.235 ;
        RECT 26.905 189.065 27.075 189.235 ;
        RECT 27.365 189.065 27.535 189.235 ;
        RECT 27.825 189.065 27.995 189.235 ;
        RECT 28.285 189.065 28.455 189.235 ;
        RECT 28.745 189.065 28.915 189.235 ;
        RECT 29.205 189.065 29.375 189.235 ;
        RECT 29.665 189.065 29.835 189.235 ;
        RECT 30.125 189.065 30.295 189.235 ;
        RECT 30.585 189.065 30.755 189.235 ;
        RECT 31.045 189.065 31.215 189.235 ;
        RECT 31.505 189.065 31.675 189.235 ;
        RECT 31.965 189.065 32.135 189.235 ;
        RECT 32.425 189.065 32.595 189.235 ;
        RECT 32.885 189.065 33.055 189.235 ;
        RECT 33.345 189.065 33.515 189.235 ;
        RECT 33.805 189.065 33.975 189.235 ;
        RECT 34.265 189.065 34.435 189.235 ;
        RECT 34.725 189.065 34.895 189.235 ;
        RECT 35.185 189.065 35.355 189.235 ;
        RECT 35.645 189.065 35.815 189.235 ;
        RECT 36.105 189.065 36.275 189.235 ;
        RECT 36.565 189.065 36.735 189.235 ;
        RECT 37.025 189.065 37.195 189.235 ;
        RECT 37.485 189.065 37.655 189.235 ;
        RECT 37.945 189.065 38.115 189.235 ;
        RECT 38.405 189.065 38.575 189.235 ;
        RECT 38.865 189.065 39.035 189.235 ;
        RECT 39.325 189.065 39.495 189.235 ;
        RECT 39.785 189.065 39.955 189.235 ;
        RECT 40.245 189.065 40.415 189.235 ;
        RECT 40.705 189.065 40.875 189.235 ;
        RECT 41.165 189.065 41.335 189.235 ;
        RECT 41.625 189.065 41.795 189.235 ;
        RECT 42.085 189.065 42.255 189.235 ;
        RECT 42.545 189.065 42.715 189.235 ;
        RECT 43.005 189.065 43.175 189.235 ;
        RECT 43.465 189.065 43.635 189.235 ;
        RECT 43.925 189.065 44.095 189.235 ;
        RECT 44.385 189.065 44.555 189.235 ;
        RECT 44.845 189.065 45.015 189.235 ;
        RECT 45.305 189.065 45.475 189.235 ;
        RECT 45.765 189.065 45.935 189.235 ;
        RECT 46.225 189.065 46.395 189.235 ;
        RECT 46.685 189.065 46.855 189.235 ;
        RECT 47.145 189.065 47.315 189.235 ;
        RECT 47.605 189.065 47.775 189.235 ;
        RECT 48.065 189.065 48.235 189.235 ;
        RECT 48.525 189.065 48.695 189.235 ;
        RECT 48.985 189.065 49.155 189.235 ;
        RECT 49.445 189.065 49.615 189.235 ;
        RECT 49.905 189.065 50.075 189.235 ;
        RECT 50.365 189.065 50.535 189.235 ;
        RECT 50.825 189.065 50.995 189.235 ;
        RECT 51.285 189.065 51.455 189.235 ;
        RECT 51.745 189.065 51.915 189.235 ;
        RECT 52.205 189.065 52.375 189.235 ;
        RECT 52.665 189.065 52.835 189.235 ;
        RECT 53.125 189.065 53.295 189.235 ;
        RECT 53.585 189.065 53.755 189.235 ;
        RECT 54.045 189.065 54.215 189.235 ;
        RECT 54.505 189.065 54.675 189.235 ;
        RECT 54.965 189.065 55.135 189.235 ;
        RECT 55.425 189.065 55.595 189.235 ;
        RECT 55.885 189.065 56.055 189.235 ;
        RECT 56.345 189.065 56.515 189.235 ;
        RECT 56.805 189.065 56.975 189.235 ;
        RECT 57.265 189.065 57.435 189.235 ;
        RECT 57.725 189.065 57.895 189.235 ;
        RECT 58.185 189.065 58.355 189.235 ;
        RECT 58.645 189.065 58.815 189.235 ;
        RECT 59.105 189.065 59.275 189.235 ;
        RECT 59.565 189.065 59.735 189.235 ;
        RECT 60.025 189.065 60.195 189.235 ;
        RECT 60.485 189.065 60.655 189.235 ;
        RECT 60.945 189.065 61.115 189.235 ;
        RECT 61.405 189.065 61.575 189.235 ;
        RECT 61.865 189.065 62.035 189.235 ;
        RECT 62.325 189.065 62.495 189.235 ;
        RECT 62.785 189.065 62.955 189.235 ;
        RECT 63.245 189.065 63.415 189.235 ;
        RECT 63.705 189.065 63.875 189.235 ;
        RECT 64.165 189.065 64.335 189.235 ;
        RECT 64.625 189.065 64.795 189.235 ;
        RECT 65.085 189.065 65.255 189.235 ;
        RECT 65.545 189.065 65.715 189.235 ;
        RECT 66.005 189.065 66.175 189.235 ;
        RECT 66.465 189.065 66.635 189.235 ;
        RECT 66.925 189.065 67.095 189.235 ;
        RECT 67.385 189.065 67.555 189.235 ;
        RECT 67.845 189.065 68.015 189.235 ;
        RECT 68.305 189.065 68.475 189.235 ;
        RECT 68.765 189.065 68.935 189.235 ;
        RECT 69.225 189.065 69.395 189.235 ;
        RECT 69.685 189.065 69.855 189.235 ;
        RECT 70.145 189.065 70.315 189.235 ;
        RECT 70.605 189.065 70.775 189.235 ;
        RECT 71.065 189.065 71.235 189.235 ;
        RECT 71.525 189.065 71.695 189.235 ;
        RECT 71.985 189.065 72.155 189.235 ;
        RECT 72.445 189.065 72.615 189.235 ;
        RECT 72.905 189.065 73.075 189.235 ;
        RECT 73.365 189.065 73.535 189.235 ;
        RECT 73.825 189.065 73.995 189.235 ;
        RECT 74.285 189.065 74.455 189.235 ;
        RECT 74.745 189.065 74.915 189.235 ;
        RECT 75.205 189.065 75.375 189.235 ;
        RECT 75.665 189.065 75.835 189.235 ;
        RECT 76.125 189.065 76.295 189.235 ;
        RECT 76.585 189.065 76.755 189.235 ;
        RECT 77.045 189.065 77.215 189.235 ;
        RECT 77.505 189.065 77.675 189.235 ;
        RECT 77.965 189.065 78.135 189.235 ;
        RECT 78.425 189.065 78.595 189.235 ;
        RECT 78.885 189.065 79.055 189.235 ;
        RECT 79.345 189.065 79.515 189.235 ;
        RECT 79.805 189.065 79.975 189.235 ;
        RECT 80.265 189.065 80.435 189.235 ;
        RECT 80.725 189.065 80.895 189.235 ;
        RECT 81.185 189.065 81.355 189.235 ;
        RECT 81.645 189.065 81.815 189.235 ;
        RECT 82.105 189.065 82.275 189.235 ;
        RECT 82.565 189.065 82.735 189.235 ;
        RECT 83.025 189.065 83.195 189.235 ;
        RECT 83.485 189.065 83.655 189.235 ;
        RECT 83.945 189.065 84.115 189.235 ;
        RECT 84.405 189.065 84.575 189.235 ;
        RECT 84.865 189.065 85.035 189.235 ;
        RECT 85.325 189.065 85.495 189.235 ;
        RECT 85.785 189.065 85.955 189.235 ;
        RECT 86.245 189.065 86.415 189.235 ;
        RECT 86.705 189.065 86.875 189.235 ;
        RECT 87.165 189.065 87.335 189.235 ;
        RECT 87.625 189.065 87.795 189.235 ;
        RECT 88.085 189.065 88.255 189.235 ;
        RECT 88.545 189.065 88.715 189.235 ;
        RECT 89.005 189.065 89.175 189.235 ;
        RECT 89.465 189.065 89.635 189.235 ;
        RECT 89.925 189.065 90.095 189.235 ;
        RECT 90.385 189.065 90.555 189.235 ;
        RECT 90.845 189.065 91.015 189.235 ;
        RECT 91.305 189.065 91.475 189.235 ;
        RECT 91.765 189.065 91.935 189.235 ;
        RECT 92.225 189.065 92.395 189.235 ;
        RECT 92.685 189.065 92.855 189.235 ;
        RECT 93.145 189.065 93.315 189.235 ;
        RECT 93.605 189.065 93.775 189.235 ;
        RECT 94.065 189.065 94.235 189.235 ;
        RECT 94.525 189.065 94.695 189.235 ;
        RECT 94.985 189.065 95.155 189.235 ;
        RECT 95.445 189.065 95.615 189.235 ;
        RECT 95.905 189.065 96.075 189.235 ;
        RECT 96.365 189.065 96.535 189.235 ;
        RECT 96.825 189.065 96.995 189.235 ;
        RECT 97.285 189.065 97.455 189.235 ;
        RECT 97.745 189.065 97.915 189.235 ;
        RECT 98.205 189.065 98.375 189.235 ;
        RECT 98.665 189.065 98.835 189.235 ;
        RECT 99.125 189.065 99.295 189.235 ;
        RECT 99.585 189.065 99.755 189.235 ;
        RECT 100.045 189.065 100.215 189.235 ;
        RECT 100.505 189.065 100.675 189.235 ;
        RECT 100.965 189.065 101.135 189.235 ;
        RECT 101.425 189.065 101.595 189.235 ;
        RECT 101.885 189.065 102.055 189.235 ;
        RECT 102.345 189.065 102.515 189.235 ;
        RECT 102.805 189.065 102.975 189.235 ;
        RECT 103.265 189.065 103.435 189.235 ;
        RECT 103.725 189.065 103.895 189.235 ;
        RECT 104.185 189.065 104.355 189.235 ;
        RECT 104.645 189.065 104.815 189.235 ;
        RECT 105.105 189.065 105.275 189.235 ;
        RECT 105.565 189.065 105.735 189.235 ;
        RECT 106.025 189.065 106.195 189.235 ;
        RECT 106.485 189.065 106.655 189.235 ;
        RECT 106.945 189.065 107.115 189.235 ;
        RECT 107.405 189.065 107.575 189.235 ;
        RECT 107.865 189.065 108.035 189.235 ;
        RECT 108.325 189.065 108.495 189.235 ;
        RECT 108.785 189.065 108.955 189.235 ;
        RECT 109.245 189.065 109.415 189.235 ;
        RECT 109.705 189.065 109.875 189.235 ;
        RECT 110.165 189.065 110.335 189.235 ;
        RECT 110.625 189.065 110.795 189.235 ;
        RECT 111.085 189.065 111.255 189.235 ;
        RECT 111.545 189.065 111.715 189.235 ;
        RECT 112.005 189.065 112.175 189.235 ;
        RECT 112.465 189.065 112.635 189.235 ;
        RECT 112.925 189.065 113.095 189.235 ;
        RECT 113.385 189.065 113.555 189.235 ;
        RECT 113.845 189.065 114.015 189.235 ;
        RECT 114.305 189.065 114.475 189.235 ;
        RECT 114.765 189.065 114.935 189.235 ;
        RECT 115.225 189.065 115.395 189.235 ;
        RECT 115.685 189.065 115.855 189.235 ;
        RECT 116.145 189.065 116.315 189.235 ;
        RECT 116.605 189.065 116.775 189.235 ;
        RECT 117.065 189.065 117.235 189.235 ;
        RECT 117.525 189.065 117.695 189.235 ;
        RECT 117.985 189.065 118.155 189.235 ;
        RECT 118.445 189.065 118.615 189.235 ;
        RECT 118.905 189.065 119.075 189.235 ;
        RECT 119.365 189.065 119.535 189.235 ;
        RECT 119.825 189.065 119.995 189.235 ;
        RECT 120.285 189.065 120.455 189.235 ;
        RECT 120.745 189.065 120.915 189.235 ;
        RECT 121.205 189.065 121.375 189.235 ;
        RECT 121.665 189.065 121.835 189.235 ;
        RECT 122.125 189.065 122.295 189.235 ;
        RECT 122.585 189.065 122.755 189.235 ;
        RECT 123.045 189.065 123.215 189.235 ;
        RECT 123.505 189.065 123.675 189.235 ;
        RECT 123.965 189.065 124.135 189.235 ;
        RECT 124.425 189.065 124.595 189.235 ;
        RECT 124.885 189.065 125.055 189.235 ;
        RECT 125.345 189.065 125.515 189.235 ;
        RECT 125.805 189.065 125.975 189.235 ;
        RECT 126.265 189.065 126.435 189.235 ;
        RECT 126.725 189.065 126.895 189.235 ;
        RECT 127.185 189.065 127.355 189.235 ;
        RECT 127.645 189.065 127.815 189.235 ;
        RECT 128.105 189.065 128.275 189.235 ;
        RECT 128.565 189.065 128.735 189.235 ;
        RECT 129.025 189.065 129.195 189.235 ;
        RECT 129.485 189.065 129.655 189.235 ;
        RECT 129.945 189.065 130.115 189.235 ;
        RECT 130.405 189.065 130.575 189.235 ;
        RECT 130.865 189.065 131.035 189.235 ;
        RECT 131.325 189.065 131.495 189.235 ;
        RECT 131.785 189.065 131.955 189.235 ;
        RECT 132.245 189.065 132.415 189.235 ;
        RECT 132.705 189.065 132.875 189.235 ;
        RECT 133.165 189.065 133.335 189.235 ;
        RECT 133.625 189.065 133.795 189.235 ;
        RECT 134.085 189.065 134.255 189.235 ;
        RECT 134.545 189.065 134.715 189.235 ;
        RECT 135.005 189.065 135.175 189.235 ;
        RECT 135.465 189.065 135.635 189.235 ;
        RECT 135.925 189.065 136.095 189.235 ;
        RECT 136.385 189.065 136.555 189.235 ;
        RECT 136.845 189.065 137.015 189.235 ;
        RECT 137.305 189.065 137.475 189.235 ;
        RECT 137.765 189.065 137.935 189.235 ;
        RECT 138.225 189.065 138.395 189.235 ;
        RECT 138.685 189.065 138.855 189.235 ;
        RECT 139.145 189.065 139.315 189.235 ;
        RECT 139.605 189.065 139.775 189.235 ;
        RECT 140.065 189.065 140.235 189.235 ;
        RECT 140.525 189.065 140.695 189.235 ;
        RECT 140.985 189.065 141.155 189.235 ;
        RECT 141.445 189.065 141.615 189.235 ;
        RECT 141.905 189.065 142.075 189.235 ;
        RECT 142.365 189.065 142.535 189.235 ;
        RECT 142.825 189.065 142.995 189.235 ;
        RECT 143.285 189.065 143.455 189.235 ;
        RECT 143.745 189.065 143.915 189.235 ;
        RECT 144.205 189.065 144.375 189.235 ;
        RECT 144.665 189.065 144.835 189.235 ;
        RECT 145.125 189.065 145.295 189.235 ;
        RECT 145.585 189.065 145.755 189.235 ;
        RECT 146.045 189.065 146.215 189.235 ;
        RECT 146.505 189.065 146.675 189.235 ;
        RECT 146.965 189.065 147.135 189.235 ;
        RECT 147.425 189.065 147.595 189.235 ;
        RECT 147.885 189.065 148.055 189.235 ;
        RECT 148.345 189.065 148.515 189.235 ;
        RECT 148.805 189.065 148.975 189.235 ;
        RECT 149.265 189.065 149.435 189.235 ;
        RECT 149.725 189.065 149.895 189.235 ;
        RECT 150.185 189.065 150.355 189.235 ;
        RECT 14.025 188.555 14.195 188.725 ;
        RECT 14.945 187.195 15.115 187.365 ;
        RECT 17.245 188.215 17.415 188.385 ;
        RECT 16.325 187.535 16.495 187.705 ;
        RECT 18.325 188.215 18.495 188.385 ;
        RECT 23.685 188.215 23.855 188.385 ;
        RECT 19.085 187.195 19.255 187.365 ;
        RECT 18.165 186.855 18.335 187.025 ;
        RECT 25.525 188.555 25.695 188.725 ;
        RECT 24.685 188.215 24.855 188.385 ;
        RECT 24.605 186.855 24.775 187.025 ;
        RECT 25.985 188.555 26.155 188.725 ;
        RECT 26.905 187.875 27.075 188.045 ;
        RECT 30.585 187.875 30.755 188.045 ;
        RECT 31.505 187.875 31.675 188.045 ;
        RECT 31.045 186.855 31.215 187.025 ;
        RECT 41.625 187.875 41.795 188.045 ;
        RECT 42.085 187.535 42.255 187.705 ;
        RECT 43.465 187.195 43.635 187.365 ;
        RECT 52.665 188.555 52.835 188.725 ;
        RECT 50.365 187.875 50.535 188.045 ;
        RECT 51.745 187.875 51.915 188.045 ;
        RECT 49.905 187.535 50.075 187.705 ;
        RECT 53.125 188.215 53.295 188.385 ;
        RECT 52.665 187.875 52.835 188.045 ;
        RECT 54.125 188.555 54.295 188.725 ;
        RECT 54.965 188.555 55.135 188.725 ;
        RECT 55.425 187.875 55.595 188.045 ;
        RECT 54.045 186.855 54.215 187.025 ;
        RECT 55.910 187.195 56.080 187.365 ;
        RECT 56.305 187.535 56.475 187.705 ;
        RECT 56.760 188.215 56.930 188.385 ;
        RECT 57.495 187.535 57.665 187.705 ;
        RECT 58.010 187.195 58.180 187.365 ;
        RECT 59.580 187.195 59.750 187.365 ;
        RECT 60.015 187.535 60.185 187.705 ;
        RECT 62.325 188.555 62.495 188.725 ;
        RECT 64.040 188.215 64.210 188.385 ;
        RECT 64.625 187.875 64.795 188.045 ;
        RECT 65.085 187.535 65.255 187.705 ;
        RECT 67.845 187.875 68.015 188.045 ;
        RECT 68.585 187.875 68.755 188.045 ;
        RECT 69.225 187.875 69.395 188.045 ;
        RECT 69.685 187.875 69.855 188.045 ;
        RECT 70.365 187.875 70.535 188.045 ;
        RECT 66.465 187.535 66.635 187.705 ;
        RECT 63.245 186.855 63.415 187.025 ;
        RECT 73.825 188.555 73.995 188.725 ;
        RECT 71.525 187.875 71.695 188.045 ;
        RECT 72.870 187.875 73.040 188.045 ;
        RECT 71.065 187.195 71.235 187.365 ;
        RECT 72.445 187.535 72.615 187.705 ;
        RECT 77.505 188.555 77.675 188.725 ;
        RECT 74.315 187.875 74.485 188.045 ;
        RECT 75.205 187.875 75.375 188.045 ;
        RECT 76.125 187.875 76.295 188.045 ;
        RECT 72.905 186.855 73.075 187.025 ;
        RECT 74.285 187.195 74.455 187.365 ;
        RECT 76.585 186.855 76.755 187.025 ;
        RECT 77.965 188.215 78.135 188.385 ;
        RECT 80.265 187.875 80.435 188.045 ;
        RECT 81.185 187.875 81.355 188.045 ;
        RECT 77.045 186.855 77.215 187.025 ;
        RECT 82.565 187.875 82.735 188.045 ;
        RECT 83.025 188.215 83.195 188.385 ;
        RECT 79.345 187.195 79.515 187.365 ;
        RECT 83.945 188.215 84.115 188.385 ;
        RECT 82.105 186.855 82.275 187.025 ;
        RECT 85.325 187.875 85.495 188.045 ;
        RECT 83.945 186.855 84.115 187.025 ;
        RECT 88.085 187.875 88.255 188.045 ;
        RECT 87.625 186.855 87.795 187.025 ;
        RECT 91.305 187.535 91.475 187.705 ;
        RECT 94.985 188.555 95.155 188.725 ;
        RECT 92.225 187.875 92.395 188.045 ;
        RECT 92.690 187.875 92.860 188.045 ;
        RECT 94.065 187.875 94.235 188.045 ;
        RECT 94.525 187.875 94.695 188.045 ;
        RECT 93.605 187.195 93.775 187.365 ;
        RECT 98.665 188.215 98.835 188.385 ;
        RECT 97.285 187.875 97.455 188.045 ;
        RECT 97.745 187.875 97.915 188.045 ;
        RECT 100.505 188.555 100.675 188.725 ;
        RECT 96.365 186.855 96.535 187.025 ;
        RECT 98.665 186.855 98.835 187.025 ;
        RECT 101.885 187.875 102.055 188.045 ;
        RECT 102.345 187.875 102.515 188.045 ;
        RECT 103.725 187.875 103.895 188.045 ;
        RECT 106.025 188.215 106.195 188.385 ;
        RECT 106.485 187.875 106.655 188.045 ;
        RECT 115.685 187.875 115.855 188.045 ;
        RECT 116.145 188.555 116.315 188.725 ;
        RECT 116.605 188.555 116.775 188.725 ;
        RECT 114.765 187.195 114.935 187.365 ;
        RECT 117.525 186.855 117.695 187.025 ;
        RECT 11.265 186.345 11.435 186.515 ;
        RECT 11.725 186.345 11.895 186.515 ;
        RECT 12.185 186.345 12.355 186.515 ;
        RECT 12.645 186.345 12.815 186.515 ;
        RECT 13.105 186.345 13.275 186.515 ;
        RECT 13.565 186.345 13.735 186.515 ;
        RECT 14.025 186.345 14.195 186.515 ;
        RECT 14.485 186.345 14.655 186.515 ;
        RECT 14.945 186.345 15.115 186.515 ;
        RECT 15.405 186.345 15.575 186.515 ;
        RECT 15.865 186.345 16.035 186.515 ;
        RECT 16.325 186.345 16.495 186.515 ;
        RECT 16.785 186.345 16.955 186.515 ;
        RECT 17.245 186.345 17.415 186.515 ;
        RECT 17.705 186.345 17.875 186.515 ;
        RECT 18.165 186.345 18.335 186.515 ;
        RECT 18.625 186.345 18.795 186.515 ;
        RECT 19.085 186.345 19.255 186.515 ;
        RECT 19.545 186.345 19.715 186.515 ;
        RECT 20.005 186.345 20.175 186.515 ;
        RECT 20.465 186.345 20.635 186.515 ;
        RECT 20.925 186.345 21.095 186.515 ;
        RECT 21.385 186.345 21.555 186.515 ;
        RECT 21.845 186.345 22.015 186.515 ;
        RECT 22.305 186.345 22.475 186.515 ;
        RECT 22.765 186.345 22.935 186.515 ;
        RECT 23.225 186.345 23.395 186.515 ;
        RECT 23.685 186.345 23.855 186.515 ;
        RECT 24.145 186.345 24.315 186.515 ;
        RECT 24.605 186.345 24.775 186.515 ;
        RECT 25.065 186.345 25.235 186.515 ;
        RECT 25.525 186.345 25.695 186.515 ;
        RECT 25.985 186.345 26.155 186.515 ;
        RECT 26.445 186.345 26.615 186.515 ;
        RECT 26.905 186.345 27.075 186.515 ;
        RECT 27.365 186.345 27.535 186.515 ;
        RECT 27.825 186.345 27.995 186.515 ;
        RECT 28.285 186.345 28.455 186.515 ;
        RECT 28.745 186.345 28.915 186.515 ;
        RECT 29.205 186.345 29.375 186.515 ;
        RECT 29.665 186.345 29.835 186.515 ;
        RECT 30.125 186.345 30.295 186.515 ;
        RECT 30.585 186.345 30.755 186.515 ;
        RECT 31.045 186.345 31.215 186.515 ;
        RECT 31.505 186.345 31.675 186.515 ;
        RECT 31.965 186.345 32.135 186.515 ;
        RECT 32.425 186.345 32.595 186.515 ;
        RECT 32.885 186.345 33.055 186.515 ;
        RECT 33.345 186.345 33.515 186.515 ;
        RECT 33.805 186.345 33.975 186.515 ;
        RECT 34.265 186.345 34.435 186.515 ;
        RECT 34.725 186.345 34.895 186.515 ;
        RECT 35.185 186.345 35.355 186.515 ;
        RECT 35.645 186.345 35.815 186.515 ;
        RECT 36.105 186.345 36.275 186.515 ;
        RECT 36.565 186.345 36.735 186.515 ;
        RECT 37.025 186.345 37.195 186.515 ;
        RECT 37.485 186.345 37.655 186.515 ;
        RECT 37.945 186.345 38.115 186.515 ;
        RECT 38.405 186.345 38.575 186.515 ;
        RECT 38.865 186.345 39.035 186.515 ;
        RECT 39.325 186.345 39.495 186.515 ;
        RECT 39.785 186.345 39.955 186.515 ;
        RECT 40.245 186.345 40.415 186.515 ;
        RECT 40.705 186.345 40.875 186.515 ;
        RECT 41.165 186.345 41.335 186.515 ;
        RECT 41.625 186.345 41.795 186.515 ;
        RECT 42.085 186.345 42.255 186.515 ;
        RECT 42.545 186.345 42.715 186.515 ;
        RECT 43.005 186.345 43.175 186.515 ;
        RECT 43.465 186.345 43.635 186.515 ;
        RECT 43.925 186.345 44.095 186.515 ;
        RECT 44.385 186.345 44.555 186.515 ;
        RECT 44.845 186.345 45.015 186.515 ;
        RECT 45.305 186.345 45.475 186.515 ;
        RECT 45.765 186.345 45.935 186.515 ;
        RECT 46.225 186.345 46.395 186.515 ;
        RECT 46.685 186.345 46.855 186.515 ;
        RECT 47.145 186.345 47.315 186.515 ;
        RECT 47.605 186.345 47.775 186.515 ;
        RECT 48.065 186.345 48.235 186.515 ;
        RECT 48.525 186.345 48.695 186.515 ;
        RECT 48.985 186.345 49.155 186.515 ;
        RECT 49.445 186.345 49.615 186.515 ;
        RECT 49.905 186.345 50.075 186.515 ;
        RECT 50.365 186.345 50.535 186.515 ;
        RECT 50.825 186.345 50.995 186.515 ;
        RECT 51.285 186.345 51.455 186.515 ;
        RECT 51.745 186.345 51.915 186.515 ;
        RECT 52.205 186.345 52.375 186.515 ;
        RECT 52.665 186.345 52.835 186.515 ;
        RECT 53.125 186.345 53.295 186.515 ;
        RECT 53.585 186.345 53.755 186.515 ;
        RECT 54.045 186.345 54.215 186.515 ;
        RECT 54.505 186.345 54.675 186.515 ;
        RECT 54.965 186.345 55.135 186.515 ;
        RECT 55.425 186.345 55.595 186.515 ;
        RECT 55.885 186.345 56.055 186.515 ;
        RECT 56.345 186.345 56.515 186.515 ;
        RECT 56.805 186.345 56.975 186.515 ;
        RECT 57.265 186.345 57.435 186.515 ;
        RECT 57.725 186.345 57.895 186.515 ;
        RECT 58.185 186.345 58.355 186.515 ;
        RECT 58.645 186.345 58.815 186.515 ;
        RECT 59.105 186.345 59.275 186.515 ;
        RECT 59.565 186.345 59.735 186.515 ;
        RECT 60.025 186.345 60.195 186.515 ;
        RECT 60.485 186.345 60.655 186.515 ;
        RECT 60.945 186.345 61.115 186.515 ;
        RECT 61.405 186.345 61.575 186.515 ;
        RECT 61.865 186.345 62.035 186.515 ;
        RECT 62.325 186.345 62.495 186.515 ;
        RECT 62.785 186.345 62.955 186.515 ;
        RECT 63.245 186.345 63.415 186.515 ;
        RECT 63.705 186.345 63.875 186.515 ;
        RECT 64.165 186.345 64.335 186.515 ;
        RECT 64.625 186.345 64.795 186.515 ;
        RECT 65.085 186.345 65.255 186.515 ;
        RECT 65.545 186.345 65.715 186.515 ;
        RECT 66.005 186.345 66.175 186.515 ;
        RECT 66.465 186.345 66.635 186.515 ;
        RECT 66.925 186.345 67.095 186.515 ;
        RECT 67.385 186.345 67.555 186.515 ;
        RECT 67.845 186.345 68.015 186.515 ;
        RECT 68.305 186.345 68.475 186.515 ;
        RECT 68.765 186.345 68.935 186.515 ;
        RECT 69.225 186.345 69.395 186.515 ;
        RECT 69.685 186.345 69.855 186.515 ;
        RECT 70.145 186.345 70.315 186.515 ;
        RECT 70.605 186.345 70.775 186.515 ;
        RECT 71.065 186.345 71.235 186.515 ;
        RECT 71.525 186.345 71.695 186.515 ;
        RECT 71.985 186.345 72.155 186.515 ;
        RECT 72.445 186.345 72.615 186.515 ;
        RECT 72.905 186.345 73.075 186.515 ;
        RECT 73.365 186.345 73.535 186.515 ;
        RECT 73.825 186.345 73.995 186.515 ;
        RECT 74.285 186.345 74.455 186.515 ;
        RECT 74.745 186.345 74.915 186.515 ;
        RECT 75.205 186.345 75.375 186.515 ;
        RECT 75.665 186.345 75.835 186.515 ;
        RECT 76.125 186.345 76.295 186.515 ;
        RECT 76.585 186.345 76.755 186.515 ;
        RECT 77.045 186.345 77.215 186.515 ;
        RECT 77.505 186.345 77.675 186.515 ;
        RECT 77.965 186.345 78.135 186.515 ;
        RECT 78.425 186.345 78.595 186.515 ;
        RECT 78.885 186.345 79.055 186.515 ;
        RECT 79.345 186.345 79.515 186.515 ;
        RECT 79.805 186.345 79.975 186.515 ;
        RECT 80.265 186.345 80.435 186.515 ;
        RECT 80.725 186.345 80.895 186.515 ;
        RECT 81.185 186.345 81.355 186.515 ;
        RECT 81.645 186.345 81.815 186.515 ;
        RECT 82.105 186.345 82.275 186.515 ;
        RECT 82.565 186.345 82.735 186.515 ;
        RECT 83.025 186.345 83.195 186.515 ;
        RECT 83.485 186.345 83.655 186.515 ;
        RECT 83.945 186.345 84.115 186.515 ;
        RECT 84.405 186.345 84.575 186.515 ;
        RECT 84.865 186.345 85.035 186.515 ;
        RECT 85.325 186.345 85.495 186.515 ;
        RECT 85.785 186.345 85.955 186.515 ;
        RECT 86.245 186.345 86.415 186.515 ;
        RECT 86.705 186.345 86.875 186.515 ;
        RECT 87.165 186.345 87.335 186.515 ;
        RECT 87.625 186.345 87.795 186.515 ;
        RECT 88.085 186.345 88.255 186.515 ;
        RECT 88.545 186.345 88.715 186.515 ;
        RECT 89.005 186.345 89.175 186.515 ;
        RECT 89.465 186.345 89.635 186.515 ;
        RECT 89.925 186.345 90.095 186.515 ;
        RECT 90.385 186.345 90.555 186.515 ;
        RECT 90.845 186.345 91.015 186.515 ;
        RECT 91.305 186.345 91.475 186.515 ;
        RECT 91.765 186.345 91.935 186.515 ;
        RECT 92.225 186.345 92.395 186.515 ;
        RECT 92.685 186.345 92.855 186.515 ;
        RECT 93.145 186.345 93.315 186.515 ;
        RECT 93.605 186.345 93.775 186.515 ;
        RECT 94.065 186.345 94.235 186.515 ;
        RECT 94.525 186.345 94.695 186.515 ;
        RECT 94.985 186.345 95.155 186.515 ;
        RECT 95.445 186.345 95.615 186.515 ;
        RECT 95.905 186.345 96.075 186.515 ;
        RECT 96.365 186.345 96.535 186.515 ;
        RECT 96.825 186.345 96.995 186.515 ;
        RECT 97.285 186.345 97.455 186.515 ;
        RECT 97.745 186.345 97.915 186.515 ;
        RECT 98.205 186.345 98.375 186.515 ;
        RECT 98.665 186.345 98.835 186.515 ;
        RECT 99.125 186.345 99.295 186.515 ;
        RECT 99.585 186.345 99.755 186.515 ;
        RECT 100.045 186.345 100.215 186.515 ;
        RECT 100.505 186.345 100.675 186.515 ;
        RECT 100.965 186.345 101.135 186.515 ;
        RECT 101.425 186.345 101.595 186.515 ;
        RECT 101.885 186.345 102.055 186.515 ;
        RECT 102.345 186.345 102.515 186.515 ;
        RECT 102.805 186.345 102.975 186.515 ;
        RECT 103.265 186.345 103.435 186.515 ;
        RECT 103.725 186.345 103.895 186.515 ;
        RECT 104.185 186.345 104.355 186.515 ;
        RECT 104.645 186.345 104.815 186.515 ;
        RECT 105.105 186.345 105.275 186.515 ;
        RECT 105.565 186.345 105.735 186.515 ;
        RECT 106.025 186.345 106.195 186.515 ;
        RECT 106.485 186.345 106.655 186.515 ;
        RECT 106.945 186.345 107.115 186.515 ;
        RECT 107.405 186.345 107.575 186.515 ;
        RECT 107.865 186.345 108.035 186.515 ;
        RECT 108.325 186.345 108.495 186.515 ;
        RECT 108.785 186.345 108.955 186.515 ;
        RECT 109.245 186.345 109.415 186.515 ;
        RECT 109.705 186.345 109.875 186.515 ;
        RECT 110.165 186.345 110.335 186.515 ;
        RECT 110.625 186.345 110.795 186.515 ;
        RECT 111.085 186.345 111.255 186.515 ;
        RECT 111.545 186.345 111.715 186.515 ;
        RECT 112.005 186.345 112.175 186.515 ;
        RECT 112.465 186.345 112.635 186.515 ;
        RECT 112.925 186.345 113.095 186.515 ;
        RECT 113.385 186.345 113.555 186.515 ;
        RECT 113.845 186.345 114.015 186.515 ;
        RECT 114.305 186.345 114.475 186.515 ;
        RECT 114.765 186.345 114.935 186.515 ;
        RECT 115.225 186.345 115.395 186.515 ;
        RECT 115.685 186.345 115.855 186.515 ;
        RECT 116.145 186.345 116.315 186.515 ;
        RECT 116.605 186.345 116.775 186.515 ;
        RECT 117.065 186.345 117.235 186.515 ;
        RECT 117.525 186.345 117.695 186.515 ;
        RECT 117.985 186.345 118.155 186.515 ;
        RECT 118.445 186.345 118.615 186.515 ;
        RECT 118.905 186.345 119.075 186.515 ;
        RECT 119.365 186.345 119.535 186.515 ;
        RECT 119.825 186.345 119.995 186.515 ;
        RECT 120.285 186.345 120.455 186.515 ;
        RECT 120.745 186.345 120.915 186.515 ;
        RECT 121.205 186.345 121.375 186.515 ;
        RECT 121.665 186.345 121.835 186.515 ;
        RECT 122.125 186.345 122.295 186.515 ;
        RECT 122.585 186.345 122.755 186.515 ;
        RECT 123.045 186.345 123.215 186.515 ;
        RECT 123.505 186.345 123.675 186.515 ;
        RECT 123.965 186.345 124.135 186.515 ;
        RECT 124.425 186.345 124.595 186.515 ;
        RECT 124.885 186.345 125.055 186.515 ;
        RECT 125.345 186.345 125.515 186.515 ;
        RECT 125.805 186.345 125.975 186.515 ;
        RECT 126.265 186.345 126.435 186.515 ;
        RECT 126.725 186.345 126.895 186.515 ;
        RECT 127.185 186.345 127.355 186.515 ;
        RECT 127.645 186.345 127.815 186.515 ;
        RECT 128.105 186.345 128.275 186.515 ;
        RECT 128.565 186.345 128.735 186.515 ;
        RECT 129.025 186.345 129.195 186.515 ;
        RECT 129.485 186.345 129.655 186.515 ;
        RECT 129.945 186.345 130.115 186.515 ;
        RECT 130.405 186.345 130.575 186.515 ;
        RECT 130.865 186.345 131.035 186.515 ;
        RECT 131.325 186.345 131.495 186.515 ;
        RECT 131.785 186.345 131.955 186.515 ;
        RECT 132.245 186.345 132.415 186.515 ;
        RECT 132.705 186.345 132.875 186.515 ;
        RECT 133.165 186.345 133.335 186.515 ;
        RECT 133.625 186.345 133.795 186.515 ;
        RECT 134.085 186.345 134.255 186.515 ;
        RECT 134.545 186.345 134.715 186.515 ;
        RECT 135.005 186.345 135.175 186.515 ;
        RECT 135.465 186.345 135.635 186.515 ;
        RECT 135.925 186.345 136.095 186.515 ;
        RECT 136.385 186.345 136.555 186.515 ;
        RECT 136.845 186.345 137.015 186.515 ;
        RECT 137.305 186.345 137.475 186.515 ;
        RECT 137.765 186.345 137.935 186.515 ;
        RECT 138.225 186.345 138.395 186.515 ;
        RECT 138.685 186.345 138.855 186.515 ;
        RECT 139.145 186.345 139.315 186.515 ;
        RECT 139.605 186.345 139.775 186.515 ;
        RECT 140.065 186.345 140.235 186.515 ;
        RECT 140.525 186.345 140.695 186.515 ;
        RECT 140.985 186.345 141.155 186.515 ;
        RECT 141.445 186.345 141.615 186.515 ;
        RECT 141.905 186.345 142.075 186.515 ;
        RECT 142.365 186.345 142.535 186.515 ;
        RECT 142.825 186.345 142.995 186.515 ;
        RECT 143.285 186.345 143.455 186.515 ;
        RECT 143.745 186.345 143.915 186.515 ;
        RECT 144.205 186.345 144.375 186.515 ;
        RECT 144.665 186.345 144.835 186.515 ;
        RECT 145.125 186.345 145.295 186.515 ;
        RECT 145.585 186.345 145.755 186.515 ;
        RECT 146.045 186.345 146.215 186.515 ;
        RECT 146.505 186.345 146.675 186.515 ;
        RECT 146.965 186.345 147.135 186.515 ;
        RECT 147.425 186.345 147.595 186.515 ;
        RECT 147.885 186.345 148.055 186.515 ;
        RECT 148.345 186.345 148.515 186.515 ;
        RECT 148.805 186.345 148.975 186.515 ;
        RECT 149.265 186.345 149.435 186.515 ;
        RECT 149.725 186.345 149.895 186.515 ;
        RECT 150.185 186.345 150.355 186.515 ;
        RECT 19.085 185.835 19.255 186.005 ;
        RECT 17.245 184.815 17.415 184.985 ;
        RECT 18.165 184.815 18.335 184.985 ;
        RECT 20.005 185.495 20.175 185.665 ;
        RECT 19.545 184.815 19.715 184.985 ;
        RECT 20.465 184.815 20.635 184.985 ;
        RECT 24.605 185.835 24.775 186.005 ;
        RECT 27.365 185.835 27.535 186.005 ;
        RECT 25.525 184.815 25.695 184.985 ;
        RECT 26.905 184.815 27.075 184.985 ;
        RECT 27.365 184.815 27.535 184.985 ;
        RECT 27.825 184.815 27.995 184.985 ;
        RECT 26.445 184.475 26.615 184.645 ;
        RECT 28.745 184.475 28.915 184.645 ;
        RECT 31.965 185.155 32.135 185.325 ;
        RECT 35.185 185.495 35.355 185.665 ;
        RECT 31.045 184.475 31.215 184.645 ;
        RECT 32.425 184.815 32.595 184.985 ;
        RECT 33.345 184.815 33.515 184.985 ;
        RECT 33.805 184.815 33.975 184.985 ;
        RECT 34.265 184.815 34.435 184.985 ;
        RECT 36.105 185.155 36.275 185.325 ;
        RECT 40.245 185.835 40.415 186.005 ;
        RECT 35.645 184.815 35.815 184.985 ;
        RECT 36.565 184.815 36.735 184.985 ;
        RECT 37.485 184.815 37.655 184.985 ;
        RECT 42.545 185.495 42.715 185.665 ;
        RECT 39.325 184.815 39.495 184.985 ;
        RECT 41.625 184.815 41.795 184.985 ;
        RECT 37.945 184.135 38.115 184.305 ;
        RECT 38.405 184.135 38.575 184.305 ;
        RECT 40.245 184.475 40.415 184.645 ;
        RECT 39.325 184.135 39.495 184.305 ;
        RECT 47.145 185.495 47.315 185.665 ;
        RECT 48.065 185.835 48.235 186.005 ;
        RECT 46.685 184.815 46.855 184.985 ;
        RECT 46.225 184.475 46.395 184.645 ;
        RECT 48.065 184.475 48.235 184.645 ;
        RECT 50.825 184.815 50.995 184.985 ;
        RECT 51.285 184.815 51.455 184.985 ;
        RECT 51.745 185.155 51.915 185.325 ;
        RECT 52.205 185.155 52.375 185.325 ;
        RECT 64.625 185.835 64.795 186.005 ;
        RECT 63.245 184.815 63.415 184.985 ;
        RECT 53.125 184.135 53.295 184.305 ;
        RECT 64.165 184.815 64.335 184.985 ;
        RECT 64.625 184.815 64.795 184.985 ;
        RECT 69.225 185.835 69.395 186.005 ;
        RECT 67.385 184.815 67.555 184.985 ;
        RECT 68.305 184.815 68.475 184.985 ;
        RECT 71.065 185.835 71.235 186.005 ;
        RECT 72.905 185.835 73.075 186.005 ;
        RECT 72.445 184.815 72.615 184.985 ;
        RECT 72.905 184.815 73.075 184.985 ;
        RECT 77.045 184.475 77.215 184.645 ;
        RECT 77.965 185.495 78.135 185.665 ;
        RECT 78.425 184.815 78.595 184.985 ;
        RECT 78.885 184.815 79.055 184.985 ;
        RECT 79.805 184.135 79.975 184.305 ;
        RECT 86.245 185.155 86.415 185.325 ;
        RECT 85.785 184.815 85.955 184.985 ;
        RECT 87.625 185.155 87.795 185.325 ;
        RECT 90.385 185.835 90.555 186.005 ;
        RECT 89.465 185.495 89.635 185.665 ;
        RECT 90.305 184.135 90.475 184.305 ;
        RECT 91.305 184.475 91.475 184.645 ;
        RECT 101.885 185.835 102.055 186.005 ;
        RECT 104.185 185.155 104.355 185.325 ;
        RECT 103.725 184.815 103.895 184.985 ;
        RECT 108.785 185.495 108.955 185.665 ;
        RECT 108.205 184.815 108.375 184.985 ;
        RECT 109.245 185.835 109.415 186.005 ;
        RECT 109.705 185.495 109.875 185.665 ;
        RECT 111.545 185.155 111.715 185.325 ;
        RECT 110.290 184.815 110.460 184.985 ;
        RECT 112.005 184.475 112.175 184.645 ;
        RECT 113.385 184.815 113.555 184.985 ;
        RECT 114.305 185.495 114.475 185.665 ;
        RECT 115.225 184.815 115.395 184.985 ;
        RECT 116.145 184.815 116.315 184.985 ;
        RECT 112.465 184.135 112.635 184.305 ;
        RECT 115.685 184.135 115.855 184.305 ;
        RECT 119.825 184.815 119.995 184.985 ;
        RECT 120.285 185.155 120.455 185.325 ;
        RECT 120.745 185.155 120.915 185.325 ;
        RECT 121.205 184.815 121.375 184.985 ;
        RECT 124.885 185.155 125.055 185.325 ;
        RECT 125.805 184.815 125.975 184.985 ;
        RECT 118.905 184.135 119.075 184.305 ;
        RECT 128.130 185.495 128.300 185.665 ;
        RECT 127.645 185.155 127.815 185.325 ;
        RECT 126.725 184.135 126.895 184.305 ;
        RECT 128.525 185.155 128.695 185.325 ;
        RECT 128.980 184.475 129.150 184.645 ;
        RECT 130.230 185.495 130.400 185.665 ;
        RECT 129.715 185.155 129.885 185.325 ;
        RECT 131.800 185.495 131.970 185.665 ;
        RECT 132.235 185.155 132.405 185.325 ;
        RECT 134.545 184.135 134.715 184.305 ;
        RECT 11.265 183.625 11.435 183.795 ;
        RECT 11.725 183.625 11.895 183.795 ;
        RECT 12.185 183.625 12.355 183.795 ;
        RECT 12.645 183.625 12.815 183.795 ;
        RECT 13.105 183.625 13.275 183.795 ;
        RECT 13.565 183.625 13.735 183.795 ;
        RECT 14.025 183.625 14.195 183.795 ;
        RECT 14.485 183.625 14.655 183.795 ;
        RECT 14.945 183.625 15.115 183.795 ;
        RECT 15.405 183.625 15.575 183.795 ;
        RECT 15.865 183.625 16.035 183.795 ;
        RECT 16.325 183.625 16.495 183.795 ;
        RECT 16.785 183.625 16.955 183.795 ;
        RECT 17.245 183.625 17.415 183.795 ;
        RECT 17.705 183.625 17.875 183.795 ;
        RECT 18.165 183.625 18.335 183.795 ;
        RECT 18.625 183.625 18.795 183.795 ;
        RECT 19.085 183.625 19.255 183.795 ;
        RECT 19.545 183.625 19.715 183.795 ;
        RECT 20.005 183.625 20.175 183.795 ;
        RECT 20.465 183.625 20.635 183.795 ;
        RECT 20.925 183.625 21.095 183.795 ;
        RECT 21.385 183.625 21.555 183.795 ;
        RECT 21.845 183.625 22.015 183.795 ;
        RECT 22.305 183.625 22.475 183.795 ;
        RECT 22.765 183.625 22.935 183.795 ;
        RECT 23.225 183.625 23.395 183.795 ;
        RECT 23.685 183.625 23.855 183.795 ;
        RECT 24.145 183.625 24.315 183.795 ;
        RECT 24.605 183.625 24.775 183.795 ;
        RECT 25.065 183.625 25.235 183.795 ;
        RECT 25.525 183.625 25.695 183.795 ;
        RECT 25.985 183.625 26.155 183.795 ;
        RECT 26.445 183.625 26.615 183.795 ;
        RECT 26.905 183.625 27.075 183.795 ;
        RECT 27.365 183.625 27.535 183.795 ;
        RECT 27.825 183.625 27.995 183.795 ;
        RECT 28.285 183.625 28.455 183.795 ;
        RECT 28.745 183.625 28.915 183.795 ;
        RECT 29.205 183.625 29.375 183.795 ;
        RECT 29.665 183.625 29.835 183.795 ;
        RECT 30.125 183.625 30.295 183.795 ;
        RECT 30.585 183.625 30.755 183.795 ;
        RECT 31.045 183.625 31.215 183.795 ;
        RECT 31.505 183.625 31.675 183.795 ;
        RECT 31.965 183.625 32.135 183.795 ;
        RECT 32.425 183.625 32.595 183.795 ;
        RECT 32.885 183.625 33.055 183.795 ;
        RECT 33.345 183.625 33.515 183.795 ;
        RECT 33.805 183.625 33.975 183.795 ;
        RECT 34.265 183.625 34.435 183.795 ;
        RECT 34.725 183.625 34.895 183.795 ;
        RECT 35.185 183.625 35.355 183.795 ;
        RECT 35.645 183.625 35.815 183.795 ;
        RECT 36.105 183.625 36.275 183.795 ;
        RECT 36.565 183.625 36.735 183.795 ;
        RECT 37.025 183.625 37.195 183.795 ;
        RECT 37.485 183.625 37.655 183.795 ;
        RECT 37.945 183.625 38.115 183.795 ;
        RECT 38.405 183.625 38.575 183.795 ;
        RECT 38.865 183.625 39.035 183.795 ;
        RECT 39.325 183.625 39.495 183.795 ;
        RECT 39.785 183.625 39.955 183.795 ;
        RECT 40.245 183.625 40.415 183.795 ;
        RECT 40.705 183.625 40.875 183.795 ;
        RECT 41.165 183.625 41.335 183.795 ;
        RECT 41.625 183.625 41.795 183.795 ;
        RECT 42.085 183.625 42.255 183.795 ;
        RECT 42.545 183.625 42.715 183.795 ;
        RECT 43.005 183.625 43.175 183.795 ;
        RECT 43.465 183.625 43.635 183.795 ;
        RECT 43.925 183.625 44.095 183.795 ;
        RECT 44.385 183.625 44.555 183.795 ;
        RECT 44.845 183.625 45.015 183.795 ;
        RECT 45.305 183.625 45.475 183.795 ;
        RECT 45.765 183.625 45.935 183.795 ;
        RECT 46.225 183.625 46.395 183.795 ;
        RECT 46.685 183.625 46.855 183.795 ;
        RECT 47.145 183.625 47.315 183.795 ;
        RECT 47.605 183.625 47.775 183.795 ;
        RECT 48.065 183.625 48.235 183.795 ;
        RECT 48.525 183.625 48.695 183.795 ;
        RECT 48.985 183.625 49.155 183.795 ;
        RECT 49.445 183.625 49.615 183.795 ;
        RECT 49.905 183.625 50.075 183.795 ;
        RECT 50.365 183.625 50.535 183.795 ;
        RECT 50.825 183.625 50.995 183.795 ;
        RECT 51.285 183.625 51.455 183.795 ;
        RECT 51.745 183.625 51.915 183.795 ;
        RECT 52.205 183.625 52.375 183.795 ;
        RECT 52.665 183.625 52.835 183.795 ;
        RECT 53.125 183.625 53.295 183.795 ;
        RECT 53.585 183.625 53.755 183.795 ;
        RECT 54.045 183.625 54.215 183.795 ;
        RECT 54.505 183.625 54.675 183.795 ;
        RECT 54.965 183.625 55.135 183.795 ;
        RECT 55.425 183.625 55.595 183.795 ;
        RECT 55.885 183.625 56.055 183.795 ;
        RECT 56.345 183.625 56.515 183.795 ;
        RECT 56.805 183.625 56.975 183.795 ;
        RECT 57.265 183.625 57.435 183.795 ;
        RECT 57.725 183.625 57.895 183.795 ;
        RECT 58.185 183.625 58.355 183.795 ;
        RECT 58.645 183.625 58.815 183.795 ;
        RECT 59.105 183.625 59.275 183.795 ;
        RECT 59.565 183.625 59.735 183.795 ;
        RECT 60.025 183.625 60.195 183.795 ;
        RECT 60.485 183.625 60.655 183.795 ;
        RECT 60.945 183.625 61.115 183.795 ;
        RECT 61.405 183.625 61.575 183.795 ;
        RECT 61.865 183.625 62.035 183.795 ;
        RECT 62.325 183.625 62.495 183.795 ;
        RECT 62.785 183.625 62.955 183.795 ;
        RECT 63.245 183.625 63.415 183.795 ;
        RECT 63.705 183.625 63.875 183.795 ;
        RECT 64.165 183.625 64.335 183.795 ;
        RECT 64.625 183.625 64.795 183.795 ;
        RECT 65.085 183.625 65.255 183.795 ;
        RECT 65.545 183.625 65.715 183.795 ;
        RECT 66.005 183.625 66.175 183.795 ;
        RECT 66.465 183.625 66.635 183.795 ;
        RECT 66.925 183.625 67.095 183.795 ;
        RECT 67.385 183.625 67.555 183.795 ;
        RECT 67.845 183.625 68.015 183.795 ;
        RECT 68.305 183.625 68.475 183.795 ;
        RECT 68.765 183.625 68.935 183.795 ;
        RECT 69.225 183.625 69.395 183.795 ;
        RECT 69.685 183.625 69.855 183.795 ;
        RECT 70.145 183.625 70.315 183.795 ;
        RECT 70.605 183.625 70.775 183.795 ;
        RECT 71.065 183.625 71.235 183.795 ;
        RECT 71.525 183.625 71.695 183.795 ;
        RECT 71.985 183.625 72.155 183.795 ;
        RECT 72.445 183.625 72.615 183.795 ;
        RECT 72.905 183.625 73.075 183.795 ;
        RECT 73.365 183.625 73.535 183.795 ;
        RECT 73.825 183.625 73.995 183.795 ;
        RECT 74.285 183.625 74.455 183.795 ;
        RECT 74.745 183.625 74.915 183.795 ;
        RECT 75.205 183.625 75.375 183.795 ;
        RECT 75.665 183.625 75.835 183.795 ;
        RECT 76.125 183.625 76.295 183.795 ;
        RECT 76.585 183.625 76.755 183.795 ;
        RECT 77.045 183.625 77.215 183.795 ;
        RECT 77.505 183.625 77.675 183.795 ;
        RECT 77.965 183.625 78.135 183.795 ;
        RECT 78.425 183.625 78.595 183.795 ;
        RECT 78.885 183.625 79.055 183.795 ;
        RECT 79.345 183.625 79.515 183.795 ;
        RECT 79.805 183.625 79.975 183.795 ;
        RECT 80.265 183.625 80.435 183.795 ;
        RECT 80.725 183.625 80.895 183.795 ;
        RECT 81.185 183.625 81.355 183.795 ;
        RECT 81.645 183.625 81.815 183.795 ;
        RECT 82.105 183.625 82.275 183.795 ;
        RECT 82.565 183.625 82.735 183.795 ;
        RECT 83.025 183.625 83.195 183.795 ;
        RECT 83.485 183.625 83.655 183.795 ;
        RECT 83.945 183.625 84.115 183.795 ;
        RECT 84.405 183.625 84.575 183.795 ;
        RECT 84.865 183.625 85.035 183.795 ;
        RECT 85.325 183.625 85.495 183.795 ;
        RECT 85.785 183.625 85.955 183.795 ;
        RECT 86.245 183.625 86.415 183.795 ;
        RECT 86.705 183.625 86.875 183.795 ;
        RECT 87.165 183.625 87.335 183.795 ;
        RECT 87.625 183.625 87.795 183.795 ;
        RECT 88.085 183.625 88.255 183.795 ;
        RECT 88.545 183.625 88.715 183.795 ;
        RECT 89.005 183.625 89.175 183.795 ;
        RECT 89.465 183.625 89.635 183.795 ;
        RECT 89.925 183.625 90.095 183.795 ;
        RECT 90.385 183.625 90.555 183.795 ;
        RECT 90.845 183.625 91.015 183.795 ;
        RECT 91.305 183.625 91.475 183.795 ;
        RECT 91.765 183.625 91.935 183.795 ;
        RECT 92.225 183.625 92.395 183.795 ;
        RECT 92.685 183.625 92.855 183.795 ;
        RECT 93.145 183.625 93.315 183.795 ;
        RECT 93.605 183.625 93.775 183.795 ;
        RECT 94.065 183.625 94.235 183.795 ;
        RECT 94.525 183.625 94.695 183.795 ;
        RECT 94.985 183.625 95.155 183.795 ;
        RECT 95.445 183.625 95.615 183.795 ;
        RECT 95.905 183.625 96.075 183.795 ;
        RECT 96.365 183.625 96.535 183.795 ;
        RECT 96.825 183.625 96.995 183.795 ;
        RECT 97.285 183.625 97.455 183.795 ;
        RECT 97.745 183.625 97.915 183.795 ;
        RECT 98.205 183.625 98.375 183.795 ;
        RECT 98.665 183.625 98.835 183.795 ;
        RECT 99.125 183.625 99.295 183.795 ;
        RECT 99.585 183.625 99.755 183.795 ;
        RECT 100.045 183.625 100.215 183.795 ;
        RECT 100.505 183.625 100.675 183.795 ;
        RECT 100.965 183.625 101.135 183.795 ;
        RECT 101.425 183.625 101.595 183.795 ;
        RECT 101.885 183.625 102.055 183.795 ;
        RECT 102.345 183.625 102.515 183.795 ;
        RECT 102.805 183.625 102.975 183.795 ;
        RECT 103.265 183.625 103.435 183.795 ;
        RECT 103.725 183.625 103.895 183.795 ;
        RECT 104.185 183.625 104.355 183.795 ;
        RECT 104.645 183.625 104.815 183.795 ;
        RECT 105.105 183.625 105.275 183.795 ;
        RECT 105.565 183.625 105.735 183.795 ;
        RECT 106.025 183.625 106.195 183.795 ;
        RECT 106.485 183.625 106.655 183.795 ;
        RECT 106.945 183.625 107.115 183.795 ;
        RECT 107.405 183.625 107.575 183.795 ;
        RECT 107.865 183.625 108.035 183.795 ;
        RECT 108.325 183.625 108.495 183.795 ;
        RECT 108.785 183.625 108.955 183.795 ;
        RECT 109.245 183.625 109.415 183.795 ;
        RECT 109.705 183.625 109.875 183.795 ;
        RECT 110.165 183.625 110.335 183.795 ;
        RECT 110.625 183.625 110.795 183.795 ;
        RECT 111.085 183.625 111.255 183.795 ;
        RECT 111.545 183.625 111.715 183.795 ;
        RECT 112.005 183.625 112.175 183.795 ;
        RECT 112.465 183.625 112.635 183.795 ;
        RECT 112.925 183.625 113.095 183.795 ;
        RECT 113.385 183.625 113.555 183.795 ;
        RECT 113.845 183.625 114.015 183.795 ;
        RECT 114.305 183.625 114.475 183.795 ;
        RECT 114.765 183.625 114.935 183.795 ;
        RECT 115.225 183.625 115.395 183.795 ;
        RECT 115.685 183.625 115.855 183.795 ;
        RECT 116.145 183.625 116.315 183.795 ;
        RECT 116.605 183.625 116.775 183.795 ;
        RECT 117.065 183.625 117.235 183.795 ;
        RECT 117.525 183.625 117.695 183.795 ;
        RECT 117.985 183.625 118.155 183.795 ;
        RECT 118.445 183.625 118.615 183.795 ;
        RECT 118.905 183.625 119.075 183.795 ;
        RECT 119.365 183.625 119.535 183.795 ;
        RECT 119.825 183.625 119.995 183.795 ;
        RECT 120.285 183.625 120.455 183.795 ;
        RECT 120.745 183.625 120.915 183.795 ;
        RECT 121.205 183.625 121.375 183.795 ;
        RECT 121.665 183.625 121.835 183.795 ;
        RECT 122.125 183.625 122.295 183.795 ;
        RECT 122.585 183.625 122.755 183.795 ;
        RECT 123.045 183.625 123.215 183.795 ;
        RECT 123.505 183.625 123.675 183.795 ;
        RECT 123.965 183.625 124.135 183.795 ;
        RECT 124.425 183.625 124.595 183.795 ;
        RECT 124.885 183.625 125.055 183.795 ;
        RECT 125.345 183.625 125.515 183.795 ;
        RECT 125.805 183.625 125.975 183.795 ;
        RECT 126.265 183.625 126.435 183.795 ;
        RECT 126.725 183.625 126.895 183.795 ;
        RECT 127.185 183.625 127.355 183.795 ;
        RECT 127.645 183.625 127.815 183.795 ;
        RECT 128.105 183.625 128.275 183.795 ;
        RECT 128.565 183.625 128.735 183.795 ;
        RECT 129.025 183.625 129.195 183.795 ;
        RECT 129.485 183.625 129.655 183.795 ;
        RECT 129.945 183.625 130.115 183.795 ;
        RECT 130.405 183.625 130.575 183.795 ;
        RECT 130.865 183.625 131.035 183.795 ;
        RECT 131.325 183.625 131.495 183.795 ;
        RECT 131.785 183.625 131.955 183.795 ;
        RECT 132.245 183.625 132.415 183.795 ;
        RECT 132.705 183.625 132.875 183.795 ;
        RECT 133.165 183.625 133.335 183.795 ;
        RECT 133.625 183.625 133.795 183.795 ;
        RECT 134.085 183.625 134.255 183.795 ;
        RECT 134.545 183.625 134.715 183.795 ;
        RECT 135.005 183.625 135.175 183.795 ;
        RECT 135.465 183.625 135.635 183.795 ;
        RECT 135.925 183.625 136.095 183.795 ;
        RECT 136.385 183.625 136.555 183.795 ;
        RECT 136.845 183.625 137.015 183.795 ;
        RECT 137.305 183.625 137.475 183.795 ;
        RECT 137.765 183.625 137.935 183.795 ;
        RECT 138.225 183.625 138.395 183.795 ;
        RECT 138.685 183.625 138.855 183.795 ;
        RECT 139.145 183.625 139.315 183.795 ;
        RECT 139.605 183.625 139.775 183.795 ;
        RECT 140.065 183.625 140.235 183.795 ;
        RECT 140.525 183.625 140.695 183.795 ;
        RECT 140.985 183.625 141.155 183.795 ;
        RECT 141.445 183.625 141.615 183.795 ;
        RECT 141.905 183.625 142.075 183.795 ;
        RECT 142.365 183.625 142.535 183.795 ;
        RECT 142.825 183.625 142.995 183.795 ;
        RECT 143.285 183.625 143.455 183.795 ;
        RECT 143.745 183.625 143.915 183.795 ;
        RECT 144.205 183.625 144.375 183.795 ;
        RECT 144.665 183.625 144.835 183.795 ;
        RECT 145.125 183.625 145.295 183.795 ;
        RECT 145.585 183.625 145.755 183.795 ;
        RECT 146.045 183.625 146.215 183.795 ;
        RECT 146.505 183.625 146.675 183.795 ;
        RECT 146.965 183.625 147.135 183.795 ;
        RECT 147.425 183.625 147.595 183.795 ;
        RECT 147.885 183.625 148.055 183.795 ;
        RECT 148.345 183.625 148.515 183.795 ;
        RECT 148.805 183.625 148.975 183.795 ;
        RECT 149.265 183.625 149.435 183.795 ;
        RECT 149.725 183.625 149.895 183.795 ;
        RECT 150.185 183.625 150.355 183.795 ;
        RECT 15.865 182.435 16.035 182.605 ;
        RECT 16.325 182.435 16.495 182.605 ;
        RECT 17.245 182.435 17.415 182.605 ;
        RECT 17.245 181.415 17.415 181.585 ;
        RECT 18.625 181.415 18.795 181.585 ;
        RECT 32.425 183.115 32.595 183.285 ;
        RECT 30.585 182.775 30.755 182.945 ;
        RECT 31.505 182.435 31.675 182.605 ;
        RECT 43.925 182.435 44.095 182.605 ;
        RECT 43.005 181.415 43.175 181.585 ;
        RECT 50.825 182.435 50.995 182.605 ;
        RECT 51.745 182.435 51.915 182.605 ;
        RECT 54.965 182.435 55.135 182.605 ;
        RECT 55.425 182.435 55.595 182.605 ;
        RECT 56.345 182.435 56.515 182.605 ;
        RECT 61.405 182.775 61.575 182.945 ;
        RECT 49.905 181.415 50.075 181.585 ;
        RECT 50.825 181.415 50.995 181.585 ;
        RECT 60.945 182.435 61.115 182.605 ;
        RECT 62.325 182.775 62.495 182.945 ;
        RECT 63.245 182.435 63.415 182.605 ;
        RECT 56.345 181.755 56.515 181.925 ;
        RECT 62.325 181.755 62.495 181.925 ;
        RECT 64.165 182.435 64.335 182.605 ;
        RECT 64.625 182.435 64.795 182.605 ;
        RECT 65.085 182.435 65.255 182.605 ;
        RECT 66.465 182.095 66.635 182.265 ;
        RECT 75.205 182.775 75.375 182.945 ;
        RECT 76.125 182.775 76.295 182.945 ;
        RECT 77.045 182.775 77.215 182.945 ;
        RECT 90.385 182.435 90.555 182.605 ;
        RECT 90.845 182.095 91.015 182.265 ;
        RECT 92.225 181.415 92.395 181.585 ;
        RECT 102.345 182.095 102.515 182.265 ;
        RECT 102.830 181.755 103.000 181.925 ;
        RECT 103.225 182.095 103.395 182.265 ;
        RECT 103.570 182.775 103.740 182.945 ;
        RECT 104.415 182.095 104.585 182.265 ;
        RECT 104.930 181.755 105.100 181.925 ;
        RECT 106.500 181.755 106.670 181.925 ;
        RECT 106.935 182.095 107.105 182.265 ;
        RECT 110.165 182.435 110.335 182.605 ;
        RECT 110.625 182.435 110.795 182.605 ;
        RECT 111.545 182.775 111.715 182.945 ;
        RECT 109.245 181.415 109.415 181.585 ;
        RECT 111.545 181.755 111.715 181.925 ;
        RECT 116.605 182.435 116.775 182.605 ;
        RECT 117.065 182.775 117.235 182.945 ;
        RECT 118.445 182.435 118.615 182.605 ;
        RECT 118.905 182.095 119.075 182.265 ;
        RECT 119.825 181.755 119.995 181.925 ;
        RECT 120.285 182.435 120.455 182.605 ;
        RECT 121.205 182.435 121.375 182.605 ;
        RECT 121.665 182.435 121.835 182.605 ;
        RECT 122.585 182.435 122.755 182.605 ;
        RECT 123.045 182.435 123.215 182.605 ;
        RECT 123.965 182.435 124.135 182.605 ;
        RECT 124.885 182.435 125.055 182.605 ;
        RECT 125.325 182.435 125.495 182.605 ;
        RECT 125.805 182.435 125.975 182.605 ;
        RECT 129.945 183.115 130.115 183.285 ;
        RECT 126.725 181.755 126.895 181.925 ;
        RECT 130.865 182.435 131.035 182.605 ;
        RECT 11.265 180.905 11.435 181.075 ;
        RECT 11.725 180.905 11.895 181.075 ;
        RECT 12.185 180.905 12.355 181.075 ;
        RECT 12.645 180.905 12.815 181.075 ;
        RECT 13.105 180.905 13.275 181.075 ;
        RECT 13.565 180.905 13.735 181.075 ;
        RECT 14.025 180.905 14.195 181.075 ;
        RECT 14.485 180.905 14.655 181.075 ;
        RECT 14.945 180.905 15.115 181.075 ;
        RECT 15.405 180.905 15.575 181.075 ;
        RECT 15.865 180.905 16.035 181.075 ;
        RECT 16.325 180.905 16.495 181.075 ;
        RECT 16.785 180.905 16.955 181.075 ;
        RECT 17.245 180.905 17.415 181.075 ;
        RECT 17.705 180.905 17.875 181.075 ;
        RECT 18.165 180.905 18.335 181.075 ;
        RECT 18.625 180.905 18.795 181.075 ;
        RECT 19.085 180.905 19.255 181.075 ;
        RECT 19.545 180.905 19.715 181.075 ;
        RECT 20.005 180.905 20.175 181.075 ;
        RECT 20.465 180.905 20.635 181.075 ;
        RECT 20.925 180.905 21.095 181.075 ;
        RECT 21.385 180.905 21.555 181.075 ;
        RECT 21.845 180.905 22.015 181.075 ;
        RECT 22.305 180.905 22.475 181.075 ;
        RECT 22.765 180.905 22.935 181.075 ;
        RECT 23.225 180.905 23.395 181.075 ;
        RECT 23.685 180.905 23.855 181.075 ;
        RECT 24.145 180.905 24.315 181.075 ;
        RECT 24.605 180.905 24.775 181.075 ;
        RECT 25.065 180.905 25.235 181.075 ;
        RECT 25.525 180.905 25.695 181.075 ;
        RECT 25.985 180.905 26.155 181.075 ;
        RECT 26.445 180.905 26.615 181.075 ;
        RECT 26.905 180.905 27.075 181.075 ;
        RECT 27.365 180.905 27.535 181.075 ;
        RECT 27.825 180.905 27.995 181.075 ;
        RECT 28.285 180.905 28.455 181.075 ;
        RECT 28.745 180.905 28.915 181.075 ;
        RECT 29.205 180.905 29.375 181.075 ;
        RECT 29.665 180.905 29.835 181.075 ;
        RECT 30.125 180.905 30.295 181.075 ;
        RECT 30.585 180.905 30.755 181.075 ;
        RECT 31.045 180.905 31.215 181.075 ;
        RECT 31.505 180.905 31.675 181.075 ;
        RECT 31.965 180.905 32.135 181.075 ;
        RECT 32.425 180.905 32.595 181.075 ;
        RECT 32.885 180.905 33.055 181.075 ;
        RECT 33.345 180.905 33.515 181.075 ;
        RECT 33.805 180.905 33.975 181.075 ;
        RECT 34.265 180.905 34.435 181.075 ;
        RECT 34.725 180.905 34.895 181.075 ;
        RECT 35.185 180.905 35.355 181.075 ;
        RECT 35.645 180.905 35.815 181.075 ;
        RECT 36.105 180.905 36.275 181.075 ;
        RECT 36.565 180.905 36.735 181.075 ;
        RECT 37.025 180.905 37.195 181.075 ;
        RECT 37.485 180.905 37.655 181.075 ;
        RECT 37.945 180.905 38.115 181.075 ;
        RECT 38.405 180.905 38.575 181.075 ;
        RECT 38.865 180.905 39.035 181.075 ;
        RECT 39.325 180.905 39.495 181.075 ;
        RECT 39.785 180.905 39.955 181.075 ;
        RECT 40.245 180.905 40.415 181.075 ;
        RECT 40.705 180.905 40.875 181.075 ;
        RECT 41.165 180.905 41.335 181.075 ;
        RECT 41.625 180.905 41.795 181.075 ;
        RECT 42.085 180.905 42.255 181.075 ;
        RECT 42.545 180.905 42.715 181.075 ;
        RECT 43.005 180.905 43.175 181.075 ;
        RECT 43.465 180.905 43.635 181.075 ;
        RECT 43.925 180.905 44.095 181.075 ;
        RECT 44.385 180.905 44.555 181.075 ;
        RECT 44.845 180.905 45.015 181.075 ;
        RECT 45.305 180.905 45.475 181.075 ;
        RECT 45.765 180.905 45.935 181.075 ;
        RECT 46.225 180.905 46.395 181.075 ;
        RECT 46.685 180.905 46.855 181.075 ;
        RECT 47.145 180.905 47.315 181.075 ;
        RECT 47.605 180.905 47.775 181.075 ;
        RECT 48.065 180.905 48.235 181.075 ;
        RECT 48.525 180.905 48.695 181.075 ;
        RECT 48.985 180.905 49.155 181.075 ;
        RECT 49.445 180.905 49.615 181.075 ;
        RECT 49.905 180.905 50.075 181.075 ;
        RECT 50.365 180.905 50.535 181.075 ;
        RECT 50.825 180.905 50.995 181.075 ;
        RECT 51.285 180.905 51.455 181.075 ;
        RECT 51.745 180.905 51.915 181.075 ;
        RECT 52.205 180.905 52.375 181.075 ;
        RECT 52.665 180.905 52.835 181.075 ;
        RECT 53.125 180.905 53.295 181.075 ;
        RECT 53.585 180.905 53.755 181.075 ;
        RECT 54.045 180.905 54.215 181.075 ;
        RECT 54.505 180.905 54.675 181.075 ;
        RECT 54.965 180.905 55.135 181.075 ;
        RECT 55.425 180.905 55.595 181.075 ;
        RECT 55.885 180.905 56.055 181.075 ;
        RECT 56.345 180.905 56.515 181.075 ;
        RECT 56.805 180.905 56.975 181.075 ;
        RECT 57.265 180.905 57.435 181.075 ;
        RECT 57.725 180.905 57.895 181.075 ;
        RECT 58.185 180.905 58.355 181.075 ;
        RECT 58.645 180.905 58.815 181.075 ;
        RECT 59.105 180.905 59.275 181.075 ;
        RECT 59.565 180.905 59.735 181.075 ;
        RECT 60.025 180.905 60.195 181.075 ;
        RECT 60.485 180.905 60.655 181.075 ;
        RECT 60.945 180.905 61.115 181.075 ;
        RECT 61.405 180.905 61.575 181.075 ;
        RECT 61.865 180.905 62.035 181.075 ;
        RECT 62.325 180.905 62.495 181.075 ;
        RECT 62.785 180.905 62.955 181.075 ;
        RECT 63.245 180.905 63.415 181.075 ;
        RECT 63.705 180.905 63.875 181.075 ;
        RECT 64.165 180.905 64.335 181.075 ;
        RECT 64.625 180.905 64.795 181.075 ;
        RECT 65.085 180.905 65.255 181.075 ;
        RECT 65.545 180.905 65.715 181.075 ;
        RECT 66.005 180.905 66.175 181.075 ;
        RECT 66.465 180.905 66.635 181.075 ;
        RECT 66.925 180.905 67.095 181.075 ;
        RECT 67.385 180.905 67.555 181.075 ;
        RECT 67.845 180.905 68.015 181.075 ;
        RECT 68.305 180.905 68.475 181.075 ;
        RECT 68.765 180.905 68.935 181.075 ;
        RECT 69.225 180.905 69.395 181.075 ;
        RECT 69.685 180.905 69.855 181.075 ;
        RECT 70.145 180.905 70.315 181.075 ;
        RECT 70.605 180.905 70.775 181.075 ;
        RECT 71.065 180.905 71.235 181.075 ;
        RECT 71.525 180.905 71.695 181.075 ;
        RECT 71.985 180.905 72.155 181.075 ;
        RECT 72.445 180.905 72.615 181.075 ;
        RECT 72.905 180.905 73.075 181.075 ;
        RECT 73.365 180.905 73.535 181.075 ;
        RECT 73.825 180.905 73.995 181.075 ;
        RECT 74.285 180.905 74.455 181.075 ;
        RECT 74.745 180.905 74.915 181.075 ;
        RECT 75.205 180.905 75.375 181.075 ;
        RECT 75.665 180.905 75.835 181.075 ;
        RECT 76.125 180.905 76.295 181.075 ;
        RECT 76.585 180.905 76.755 181.075 ;
        RECT 77.045 180.905 77.215 181.075 ;
        RECT 77.505 180.905 77.675 181.075 ;
        RECT 77.965 180.905 78.135 181.075 ;
        RECT 78.425 180.905 78.595 181.075 ;
        RECT 78.885 180.905 79.055 181.075 ;
        RECT 79.345 180.905 79.515 181.075 ;
        RECT 79.805 180.905 79.975 181.075 ;
        RECT 80.265 180.905 80.435 181.075 ;
        RECT 80.725 180.905 80.895 181.075 ;
        RECT 81.185 180.905 81.355 181.075 ;
        RECT 81.645 180.905 81.815 181.075 ;
        RECT 82.105 180.905 82.275 181.075 ;
        RECT 82.565 180.905 82.735 181.075 ;
        RECT 83.025 180.905 83.195 181.075 ;
        RECT 83.485 180.905 83.655 181.075 ;
        RECT 83.945 180.905 84.115 181.075 ;
        RECT 84.405 180.905 84.575 181.075 ;
        RECT 84.865 180.905 85.035 181.075 ;
        RECT 85.325 180.905 85.495 181.075 ;
        RECT 85.785 180.905 85.955 181.075 ;
        RECT 86.245 180.905 86.415 181.075 ;
        RECT 86.705 180.905 86.875 181.075 ;
        RECT 87.165 180.905 87.335 181.075 ;
        RECT 87.625 180.905 87.795 181.075 ;
        RECT 88.085 180.905 88.255 181.075 ;
        RECT 88.545 180.905 88.715 181.075 ;
        RECT 89.005 180.905 89.175 181.075 ;
        RECT 89.465 180.905 89.635 181.075 ;
        RECT 89.925 180.905 90.095 181.075 ;
        RECT 90.385 180.905 90.555 181.075 ;
        RECT 90.845 180.905 91.015 181.075 ;
        RECT 91.305 180.905 91.475 181.075 ;
        RECT 91.765 180.905 91.935 181.075 ;
        RECT 92.225 180.905 92.395 181.075 ;
        RECT 92.685 180.905 92.855 181.075 ;
        RECT 93.145 180.905 93.315 181.075 ;
        RECT 93.605 180.905 93.775 181.075 ;
        RECT 94.065 180.905 94.235 181.075 ;
        RECT 94.525 180.905 94.695 181.075 ;
        RECT 94.985 180.905 95.155 181.075 ;
        RECT 95.445 180.905 95.615 181.075 ;
        RECT 95.905 180.905 96.075 181.075 ;
        RECT 96.365 180.905 96.535 181.075 ;
        RECT 96.825 180.905 96.995 181.075 ;
        RECT 97.285 180.905 97.455 181.075 ;
        RECT 97.745 180.905 97.915 181.075 ;
        RECT 98.205 180.905 98.375 181.075 ;
        RECT 98.665 180.905 98.835 181.075 ;
        RECT 99.125 180.905 99.295 181.075 ;
        RECT 99.585 180.905 99.755 181.075 ;
        RECT 100.045 180.905 100.215 181.075 ;
        RECT 100.505 180.905 100.675 181.075 ;
        RECT 100.965 180.905 101.135 181.075 ;
        RECT 101.425 180.905 101.595 181.075 ;
        RECT 101.885 180.905 102.055 181.075 ;
        RECT 102.345 180.905 102.515 181.075 ;
        RECT 102.805 180.905 102.975 181.075 ;
        RECT 103.265 180.905 103.435 181.075 ;
        RECT 103.725 180.905 103.895 181.075 ;
        RECT 104.185 180.905 104.355 181.075 ;
        RECT 104.645 180.905 104.815 181.075 ;
        RECT 105.105 180.905 105.275 181.075 ;
        RECT 105.565 180.905 105.735 181.075 ;
        RECT 106.025 180.905 106.195 181.075 ;
        RECT 106.485 180.905 106.655 181.075 ;
        RECT 106.945 180.905 107.115 181.075 ;
        RECT 107.405 180.905 107.575 181.075 ;
        RECT 107.865 180.905 108.035 181.075 ;
        RECT 108.325 180.905 108.495 181.075 ;
        RECT 108.785 180.905 108.955 181.075 ;
        RECT 109.245 180.905 109.415 181.075 ;
        RECT 109.705 180.905 109.875 181.075 ;
        RECT 110.165 180.905 110.335 181.075 ;
        RECT 110.625 180.905 110.795 181.075 ;
        RECT 111.085 180.905 111.255 181.075 ;
        RECT 111.545 180.905 111.715 181.075 ;
        RECT 112.005 180.905 112.175 181.075 ;
        RECT 112.465 180.905 112.635 181.075 ;
        RECT 112.925 180.905 113.095 181.075 ;
        RECT 113.385 180.905 113.555 181.075 ;
        RECT 113.845 180.905 114.015 181.075 ;
        RECT 114.305 180.905 114.475 181.075 ;
        RECT 114.765 180.905 114.935 181.075 ;
        RECT 115.225 180.905 115.395 181.075 ;
        RECT 115.685 180.905 115.855 181.075 ;
        RECT 116.145 180.905 116.315 181.075 ;
        RECT 116.605 180.905 116.775 181.075 ;
        RECT 117.065 180.905 117.235 181.075 ;
        RECT 117.525 180.905 117.695 181.075 ;
        RECT 117.985 180.905 118.155 181.075 ;
        RECT 118.445 180.905 118.615 181.075 ;
        RECT 118.905 180.905 119.075 181.075 ;
        RECT 119.365 180.905 119.535 181.075 ;
        RECT 119.825 180.905 119.995 181.075 ;
        RECT 120.285 180.905 120.455 181.075 ;
        RECT 120.745 180.905 120.915 181.075 ;
        RECT 121.205 180.905 121.375 181.075 ;
        RECT 121.665 180.905 121.835 181.075 ;
        RECT 122.125 180.905 122.295 181.075 ;
        RECT 122.585 180.905 122.755 181.075 ;
        RECT 123.045 180.905 123.215 181.075 ;
        RECT 123.505 180.905 123.675 181.075 ;
        RECT 123.965 180.905 124.135 181.075 ;
        RECT 124.425 180.905 124.595 181.075 ;
        RECT 124.885 180.905 125.055 181.075 ;
        RECT 125.345 180.905 125.515 181.075 ;
        RECT 125.805 180.905 125.975 181.075 ;
        RECT 126.265 180.905 126.435 181.075 ;
        RECT 126.725 180.905 126.895 181.075 ;
        RECT 127.185 180.905 127.355 181.075 ;
        RECT 127.645 180.905 127.815 181.075 ;
        RECT 128.105 180.905 128.275 181.075 ;
        RECT 128.565 180.905 128.735 181.075 ;
        RECT 129.025 180.905 129.195 181.075 ;
        RECT 129.485 180.905 129.655 181.075 ;
        RECT 129.945 180.905 130.115 181.075 ;
        RECT 130.405 180.905 130.575 181.075 ;
        RECT 130.865 180.905 131.035 181.075 ;
        RECT 131.325 180.905 131.495 181.075 ;
        RECT 131.785 180.905 131.955 181.075 ;
        RECT 132.245 180.905 132.415 181.075 ;
        RECT 132.705 180.905 132.875 181.075 ;
        RECT 133.165 180.905 133.335 181.075 ;
        RECT 133.625 180.905 133.795 181.075 ;
        RECT 134.085 180.905 134.255 181.075 ;
        RECT 134.545 180.905 134.715 181.075 ;
        RECT 135.005 180.905 135.175 181.075 ;
        RECT 135.465 180.905 135.635 181.075 ;
        RECT 135.925 180.905 136.095 181.075 ;
        RECT 136.385 180.905 136.555 181.075 ;
        RECT 136.845 180.905 137.015 181.075 ;
        RECT 137.305 180.905 137.475 181.075 ;
        RECT 137.765 180.905 137.935 181.075 ;
        RECT 138.225 180.905 138.395 181.075 ;
        RECT 138.685 180.905 138.855 181.075 ;
        RECT 139.145 180.905 139.315 181.075 ;
        RECT 139.605 180.905 139.775 181.075 ;
        RECT 140.065 180.905 140.235 181.075 ;
        RECT 140.525 180.905 140.695 181.075 ;
        RECT 140.985 180.905 141.155 181.075 ;
        RECT 141.445 180.905 141.615 181.075 ;
        RECT 141.905 180.905 142.075 181.075 ;
        RECT 142.365 180.905 142.535 181.075 ;
        RECT 142.825 180.905 142.995 181.075 ;
        RECT 143.285 180.905 143.455 181.075 ;
        RECT 143.745 180.905 143.915 181.075 ;
        RECT 144.205 180.905 144.375 181.075 ;
        RECT 144.665 180.905 144.835 181.075 ;
        RECT 145.125 180.905 145.295 181.075 ;
        RECT 145.585 180.905 145.755 181.075 ;
        RECT 146.045 180.905 146.215 181.075 ;
        RECT 146.505 180.905 146.675 181.075 ;
        RECT 146.965 180.905 147.135 181.075 ;
        RECT 147.425 180.905 147.595 181.075 ;
        RECT 147.885 180.905 148.055 181.075 ;
        RECT 148.345 180.905 148.515 181.075 ;
        RECT 148.805 180.905 148.975 181.075 ;
        RECT 149.265 180.905 149.435 181.075 ;
        RECT 149.725 180.905 149.895 181.075 ;
        RECT 150.185 180.905 150.355 181.075 ;
        RECT 14.050 180.055 14.220 180.225 ;
        RECT 13.565 179.375 13.735 179.545 ;
        RECT 14.445 179.715 14.615 179.885 ;
        RECT 14.900 179.375 15.070 179.545 ;
        RECT 16.150 180.055 16.320 180.225 ;
        RECT 15.635 179.715 15.805 179.885 ;
        RECT 17.720 180.055 17.890 180.225 ;
        RECT 18.155 179.715 18.325 179.885 ;
        RECT 20.465 180.395 20.635 180.565 ;
        RECT 23.685 180.055 23.855 180.225 ;
        RECT 22.305 179.375 22.475 179.545 ;
        RECT 25.090 180.055 25.260 180.225 ;
        RECT 22.765 178.695 22.935 178.865 ;
        RECT 24.605 179.375 24.775 179.545 ;
        RECT 23.685 179.035 23.855 179.205 ;
        RECT 25.485 179.715 25.655 179.885 ;
        RECT 25.830 179.035 26.000 179.205 ;
        RECT 27.190 180.055 27.360 180.225 ;
        RECT 26.675 179.715 26.845 179.885 ;
        RECT 28.760 180.055 28.930 180.225 ;
        RECT 29.195 179.715 29.365 179.885 ;
        RECT 31.505 178.695 31.675 178.865 ;
        RECT 35.645 180.395 35.815 180.565 ;
        RECT 36.590 180.055 36.760 180.225 ;
        RECT 33.345 179.375 33.515 179.545 ;
        RECT 34.725 179.375 34.895 179.545 ;
        RECT 36.105 179.715 36.275 179.885 ;
        RECT 35.645 179.375 35.815 179.545 ;
        RECT 32.425 178.695 32.595 178.865 ;
        RECT 36.985 179.715 37.155 179.885 ;
        RECT 37.440 179.035 37.610 179.205 ;
        RECT 38.690 180.055 38.860 180.225 ;
        RECT 38.175 179.715 38.345 179.885 ;
        RECT 40.260 180.055 40.430 180.225 ;
        RECT 40.695 179.715 40.865 179.885 ;
        RECT 43.925 179.375 44.095 179.545 ;
        RECT 45.765 179.375 45.935 179.545 ;
        RECT 47.145 179.375 47.315 179.545 ;
        RECT 47.605 179.375 47.775 179.545 ;
        RECT 43.005 178.695 43.175 178.865 ;
        RECT 50.365 180.055 50.535 180.225 ;
        RECT 51.285 180.395 51.455 180.565 ;
        RECT 51.285 179.375 51.455 179.545 ;
        RECT 53.125 179.375 53.295 179.545 ;
        RECT 55.425 180.395 55.595 180.565 ;
        RECT 67.845 180.055 68.015 180.225 ;
        RECT 56.115 179.375 56.285 179.545 ;
        RECT 56.805 179.035 56.975 179.205 ;
        RECT 58.180 179.375 58.350 179.545 ;
        RECT 58.645 179.375 58.815 179.545 ;
        RECT 60.025 179.375 60.195 179.545 ;
        RECT 57.265 179.035 57.435 179.205 ;
        RECT 60.945 179.375 61.115 179.545 ;
        RECT 60.485 179.035 60.655 179.205 ;
        RECT 67.385 179.375 67.555 179.545 ;
        RECT 68.305 179.375 68.475 179.545 ;
        RECT 79.345 180.395 79.515 180.565 ;
        RECT 80.750 180.055 80.920 180.225 ;
        RECT 78.425 179.375 78.595 179.545 ;
        RECT 80.265 179.715 80.435 179.885 ;
        RECT 79.345 179.375 79.515 179.545 ;
        RECT 81.145 179.715 81.315 179.885 ;
        RECT 81.600 179.035 81.770 179.205 ;
        RECT 82.850 180.055 83.020 180.225 ;
        RECT 82.335 179.715 82.505 179.885 ;
        RECT 84.420 180.055 84.590 180.225 ;
        RECT 84.855 179.715 85.025 179.885 ;
        RECT 89.465 180.395 89.635 180.565 ;
        RECT 89.005 179.375 89.175 179.545 ;
        RECT 89.925 179.375 90.095 179.545 ;
        RECT 90.385 180.055 90.555 180.225 ;
        RECT 91.305 179.375 91.475 179.545 ;
        RECT 87.165 178.695 87.335 178.865 ;
        RECT 87.625 178.695 87.795 178.865 ;
        RECT 91.765 179.035 91.935 179.205 ;
        RECT 95.445 180.055 95.615 180.225 ;
        RECT 94.525 179.375 94.695 179.545 ;
        RECT 96.825 179.715 96.995 179.885 ;
        RECT 97.285 179.375 97.455 179.545 ;
        RECT 98.665 179.375 98.835 179.545 ;
        RECT 99.585 179.375 99.755 179.545 ;
        RECT 99.125 179.035 99.295 179.205 ;
        RECT 104.185 180.395 104.355 180.565 ;
        RECT 103.265 179.375 103.435 179.545 ;
        RECT 112.925 179.715 113.095 179.885 ;
        RECT 114.765 180.395 114.935 180.565 ;
        RECT 112.465 179.375 112.635 179.545 ;
        RECT 113.845 179.375 114.015 179.545 ;
        RECT 118.445 180.395 118.615 180.565 ;
        RECT 115.225 179.375 115.395 179.545 ;
        RECT 116.145 179.375 116.315 179.545 ;
        RECT 116.605 178.695 116.775 178.865 ;
        RECT 120.285 179.715 120.455 179.885 ;
        RECT 119.365 179.375 119.535 179.545 ;
        RECT 124.425 180.395 124.595 180.565 ;
        RECT 124.885 179.715 125.055 179.885 ;
        RECT 125.345 179.375 125.515 179.545 ;
        RECT 127.645 179.715 127.815 179.885 ;
        RECT 128.565 180.055 128.735 180.225 ;
        RECT 129.025 179.375 129.195 179.545 ;
        RECT 123.505 178.695 123.675 178.865 ;
        RECT 11.265 178.185 11.435 178.355 ;
        RECT 11.725 178.185 11.895 178.355 ;
        RECT 12.185 178.185 12.355 178.355 ;
        RECT 12.645 178.185 12.815 178.355 ;
        RECT 13.105 178.185 13.275 178.355 ;
        RECT 13.565 178.185 13.735 178.355 ;
        RECT 14.025 178.185 14.195 178.355 ;
        RECT 14.485 178.185 14.655 178.355 ;
        RECT 14.945 178.185 15.115 178.355 ;
        RECT 15.405 178.185 15.575 178.355 ;
        RECT 15.865 178.185 16.035 178.355 ;
        RECT 16.325 178.185 16.495 178.355 ;
        RECT 16.785 178.185 16.955 178.355 ;
        RECT 17.245 178.185 17.415 178.355 ;
        RECT 17.705 178.185 17.875 178.355 ;
        RECT 18.165 178.185 18.335 178.355 ;
        RECT 18.625 178.185 18.795 178.355 ;
        RECT 19.085 178.185 19.255 178.355 ;
        RECT 19.545 178.185 19.715 178.355 ;
        RECT 20.005 178.185 20.175 178.355 ;
        RECT 20.465 178.185 20.635 178.355 ;
        RECT 20.925 178.185 21.095 178.355 ;
        RECT 21.385 178.185 21.555 178.355 ;
        RECT 21.845 178.185 22.015 178.355 ;
        RECT 22.305 178.185 22.475 178.355 ;
        RECT 22.765 178.185 22.935 178.355 ;
        RECT 23.225 178.185 23.395 178.355 ;
        RECT 23.685 178.185 23.855 178.355 ;
        RECT 24.145 178.185 24.315 178.355 ;
        RECT 24.605 178.185 24.775 178.355 ;
        RECT 25.065 178.185 25.235 178.355 ;
        RECT 25.525 178.185 25.695 178.355 ;
        RECT 25.985 178.185 26.155 178.355 ;
        RECT 26.445 178.185 26.615 178.355 ;
        RECT 26.905 178.185 27.075 178.355 ;
        RECT 27.365 178.185 27.535 178.355 ;
        RECT 27.825 178.185 27.995 178.355 ;
        RECT 28.285 178.185 28.455 178.355 ;
        RECT 28.745 178.185 28.915 178.355 ;
        RECT 29.205 178.185 29.375 178.355 ;
        RECT 29.665 178.185 29.835 178.355 ;
        RECT 30.125 178.185 30.295 178.355 ;
        RECT 30.585 178.185 30.755 178.355 ;
        RECT 31.045 178.185 31.215 178.355 ;
        RECT 31.505 178.185 31.675 178.355 ;
        RECT 31.965 178.185 32.135 178.355 ;
        RECT 32.425 178.185 32.595 178.355 ;
        RECT 32.885 178.185 33.055 178.355 ;
        RECT 33.345 178.185 33.515 178.355 ;
        RECT 33.805 178.185 33.975 178.355 ;
        RECT 34.265 178.185 34.435 178.355 ;
        RECT 34.725 178.185 34.895 178.355 ;
        RECT 35.185 178.185 35.355 178.355 ;
        RECT 35.645 178.185 35.815 178.355 ;
        RECT 36.105 178.185 36.275 178.355 ;
        RECT 36.565 178.185 36.735 178.355 ;
        RECT 37.025 178.185 37.195 178.355 ;
        RECT 37.485 178.185 37.655 178.355 ;
        RECT 37.945 178.185 38.115 178.355 ;
        RECT 38.405 178.185 38.575 178.355 ;
        RECT 38.865 178.185 39.035 178.355 ;
        RECT 39.325 178.185 39.495 178.355 ;
        RECT 39.785 178.185 39.955 178.355 ;
        RECT 40.245 178.185 40.415 178.355 ;
        RECT 40.705 178.185 40.875 178.355 ;
        RECT 41.165 178.185 41.335 178.355 ;
        RECT 41.625 178.185 41.795 178.355 ;
        RECT 42.085 178.185 42.255 178.355 ;
        RECT 42.545 178.185 42.715 178.355 ;
        RECT 43.005 178.185 43.175 178.355 ;
        RECT 43.465 178.185 43.635 178.355 ;
        RECT 43.925 178.185 44.095 178.355 ;
        RECT 44.385 178.185 44.555 178.355 ;
        RECT 44.845 178.185 45.015 178.355 ;
        RECT 45.305 178.185 45.475 178.355 ;
        RECT 45.765 178.185 45.935 178.355 ;
        RECT 46.225 178.185 46.395 178.355 ;
        RECT 46.685 178.185 46.855 178.355 ;
        RECT 47.145 178.185 47.315 178.355 ;
        RECT 47.605 178.185 47.775 178.355 ;
        RECT 48.065 178.185 48.235 178.355 ;
        RECT 48.525 178.185 48.695 178.355 ;
        RECT 48.985 178.185 49.155 178.355 ;
        RECT 49.445 178.185 49.615 178.355 ;
        RECT 49.905 178.185 50.075 178.355 ;
        RECT 50.365 178.185 50.535 178.355 ;
        RECT 50.825 178.185 50.995 178.355 ;
        RECT 51.285 178.185 51.455 178.355 ;
        RECT 51.745 178.185 51.915 178.355 ;
        RECT 52.205 178.185 52.375 178.355 ;
        RECT 52.665 178.185 52.835 178.355 ;
        RECT 53.125 178.185 53.295 178.355 ;
        RECT 53.585 178.185 53.755 178.355 ;
        RECT 54.045 178.185 54.215 178.355 ;
        RECT 54.505 178.185 54.675 178.355 ;
        RECT 54.965 178.185 55.135 178.355 ;
        RECT 55.425 178.185 55.595 178.355 ;
        RECT 55.885 178.185 56.055 178.355 ;
        RECT 56.345 178.185 56.515 178.355 ;
        RECT 56.805 178.185 56.975 178.355 ;
        RECT 57.265 178.185 57.435 178.355 ;
        RECT 57.725 178.185 57.895 178.355 ;
        RECT 58.185 178.185 58.355 178.355 ;
        RECT 58.645 178.185 58.815 178.355 ;
        RECT 59.105 178.185 59.275 178.355 ;
        RECT 59.565 178.185 59.735 178.355 ;
        RECT 60.025 178.185 60.195 178.355 ;
        RECT 60.485 178.185 60.655 178.355 ;
        RECT 60.945 178.185 61.115 178.355 ;
        RECT 61.405 178.185 61.575 178.355 ;
        RECT 61.865 178.185 62.035 178.355 ;
        RECT 62.325 178.185 62.495 178.355 ;
        RECT 62.785 178.185 62.955 178.355 ;
        RECT 63.245 178.185 63.415 178.355 ;
        RECT 63.705 178.185 63.875 178.355 ;
        RECT 64.165 178.185 64.335 178.355 ;
        RECT 64.625 178.185 64.795 178.355 ;
        RECT 65.085 178.185 65.255 178.355 ;
        RECT 65.545 178.185 65.715 178.355 ;
        RECT 66.005 178.185 66.175 178.355 ;
        RECT 66.465 178.185 66.635 178.355 ;
        RECT 66.925 178.185 67.095 178.355 ;
        RECT 67.385 178.185 67.555 178.355 ;
        RECT 67.845 178.185 68.015 178.355 ;
        RECT 68.305 178.185 68.475 178.355 ;
        RECT 68.765 178.185 68.935 178.355 ;
        RECT 69.225 178.185 69.395 178.355 ;
        RECT 69.685 178.185 69.855 178.355 ;
        RECT 70.145 178.185 70.315 178.355 ;
        RECT 70.605 178.185 70.775 178.355 ;
        RECT 71.065 178.185 71.235 178.355 ;
        RECT 71.525 178.185 71.695 178.355 ;
        RECT 71.985 178.185 72.155 178.355 ;
        RECT 72.445 178.185 72.615 178.355 ;
        RECT 72.905 178.185 73.075 178.355 ;
        RECT 73.365 178.185 73.535 178.355 ;
        RECT 73.825 178.185 73.995 178.355 ;
        RECT 74.285 178.185 74.455 178.355 ;
        RECT 74.745 178.185 74.915 178.355 ;
        RECT 75.205 178.185 75.375 178.355 ;
        RECT 75.665 178.185 75.835 178.355 ;
        RECT 76.125 178.185 76.295 178.355 ;
        RECT 76.585 178.185 76.755 178.355 ;
        RECT 77.045 178.185 77.215 178.355 ;
        RECT 77.505 178.185 77.675 178.355 ;
        RECT 77.965 178.185 78.135 178.355 ;
        RECT 78.425 178.185 78.595 178.355 ;
        RECT 78.885 178.185 79.055 178.355 ;
        RECT 79.345 178.185 79.515 178.355 ;
        RECT 79.805 178.185 79.975 178.355 ;
        RECT 80.265 178.185 80.435 178.355 ;
        RECT 80.725 178.185 80.895 178.355 ;
        RECT 81.185 178.185 81.355 178.355 ;
        RECT 81.645 178.185 81.815 178.355 ;
        RECT 82.105 178.185 82.275 178.355 ;
        RECT 82.565 178.185 82.735 178.355 ;
        RECT 83.025 178.185 83.195 178.355 ;
        RECT 83.485 178.185 83.655 178.355 ;
        RECT 83.945 178.185 84.115 178.355 ;
        RECT 84.405 178.185 84.575 178.355 ;
        RECT 84.865 178.185 85.035 178.355 ;
        RECT 85.325 178.185 85.495 178.355 ;
        RECT 85.785 178.185 85.955 178.355 ;
        RECT 86.245 178.185 86.415 178.355 ;
        RECT 86.705 178.185 86.875 178.355 ;
        RECT 87.165 178.185 87.335 178.355 ;
        RECT 87.625 178.185 87.795 178.355 ;
        RECT 88.085 178.185 88.255 178.355 ;
        RECT 88.545 178.185 88.715 178.355 ;
        RECT 89.005 178.185 89.175 178.355 ;
        RECT 89.465 178.185 89.635 178.355 ;
        RECT 89.925 178.185 90.095 178.355 ;
        RECT 90.385 178.185 90.555 178.355 ;
        RECT 90.845 178.185 91.015 178.355 ;
        RECT 91.305 178.185 91.475 178.355 ;
        RECT 91.765 178.185 91.935 178.355 ;
        RECT 92.225 178.185 92.395 178.355 ;
        RECT 92.685 178.185 92.855 178.355 ;
        RECT 93.145 178.185 93.315 178.355 ;
        RECT 93.605 178.185 93.775 178.355 ;
        RECT 94.065 178.185 94.235 178.355 ;
        RECT 94.525 178.185 94.695 178.355 ;
        RECT 94.985 178.185 95.155 178.355 ;
        RECT 95.445 178.185 95.615 178.355 ;
        RECT 95.905 178.185 96.075 178.355 ;
        RECT 96.365 178.185 96.535 178.355 ;
        RECT 96.825 178.185 96.995 178.355 ;
        RECT 97.285 178.185 97.455 178.355 ;
        RECT 97.745 178.185 97.915 178.355 ;
        RECT 98.205 178.185 98.375 178.355 ;
        RECT 98.665 178.185 98.835 178.355 ;
        RECT 99.125 178.185 99.295 178.355 ;
        RECT 99.585 178.185 99.755 178.355 ;
        RECT 100.045 178.185 100.215 178.355 ;
        RECT 100.505 178.185 100.675 178.355 ;
        RECT 100.965 178.185 101.135 178.355 ;
        RECT 101.425 178.185 101.595 178.355 ;
        RECT 101.885 178.185 102.055 178.355 ;
        RECT 102.345 178.185 102.515 178.355 ;
        RECT 102.805 178.185 102.975 178.355 ;
        RECT 103.265 178.185 103.435 178.355 ;
        RECT 103.725 178.185 103.895 178.355 ;
        RECT 104.185 178.185 104.355 178.355 ;
        RECT 104.645 178.185 104.815 178.355 ;
        RECT 105.105 178.185 105.275 178.355 ;
        RECT 105.565 178.185 105.735 178.355 ;
        RECT 106.025 178.185 106.195 178.355 ;
        RECT 106.485 178.185 106.655 178.355 ;
        RECT 106.945 178.185 107.115 178.355 ;
        RECT 107.405 178.185 107.575 178.355 ;
        RECT 107.865 178.185 108.035 178.355 ;
        RECT 108.325 178.185 108.495 178.355 ;
        RECT 108.785 178.185 108.955 178.355 ;
        RECT 109.245 178.185 109.415 178.355 ;
        RECT 109.705 178.185 109.875 178.355 ;
        RECT 110.165 178.185 110.335 178.355 ;
        RECT 110.625 178.185 110.795 178.355 ;
        RECT 111.085 178.185 111.255 178.355 ;
        RECT 111.545 178.185 111.715 178.355 ;
        RECT 112.005 178.185 112.175 178.355 ;
        RECT 112.465 178.185 112.635 178.355 ;
        RECT 112.925 178.185 113.095 178.355 ;
        RECT 113.385 178.185 113.555 178.355 ;
        RECT 113.845 178.185 114.015 178.355 ;
        RECT 114.305 178.185 114.475 178.355 ;
        RECT 114.765 178.185 114.935 178.355 ;
        RECT 115.225 178.185 115.395 178.355 ;
        RECT 115.685 178.185 115.855 178.355 ;
        RECT 116.145 178.185 116.315 178.355 ;
        RECT 116.605 178.185 116.775 178.355 ;
        RECT 117.065 178.185 117.235 178.355 ;
        RECT 117.525 178.185 117.695 178.355 ;
        RECT 117.985 178.185 118.155 178.355 ;
        RECT 118.445 178.185 118.615 178.355 ;
        RECT 118.905 178.185 119.075 178.355 ;
        RECT 119.365 178.185 119.535 178.355 ;
        RECT 119.825 178.185 119.995 178.355 ;
        RECT 120.285 178.185 120.455 178.355 ;
        RECT 120.745 178.185 120.915 178.355 ;
        RECT 121.205 178.185 121.375 178.355 ;
        RECT 121.665 178.185 121.835 178.355 ;
        RECT 122.125 178.185 122.295 178.355 ;
        RECT 122.585 178.185 122.755 178.355 ;
        RECT 123.045 178.185 123.215 178.355 ;
        RECT 123.505 178.185 123.675 178.355 ;
        RECT 123.965 178.185 124.135 178.355 ;
        RECT 124.425 178.185 124.595 178.355 ;
        RECT 124.885 178.185 125.055 178.355 ;
        RECT 125.345 178.185 125.515 178.355 ;
        RECT 125.805 178.185 125.975 178.355 ;
        RECT 126.265 178.185 126.435 178.355 ;
        RECT 126.725 178.185 126.895 178.355 ;
        RECT 127.185 178.185 127.355 178.355 ;
        RECT 127.645 178.185 127.815 178.355 ;
        RECT 128.105 178.185 128.275 178.355 ;
        RECT 128.565 178.185 128.735 178.355 ;
        RECT 129.025 178.185 129.195 178.355 ;
        RECT 129.485 178.185 129.655 178.355 ;
        RECT 129.945 178.185 130.115 178.355 ;
        RECT 130.405 178.185 130.575 178.355 ;
        RECT 130.865 178.185 131.035 178.355 ;
        RECT 131.325 178.185 131.495 178.355 ;
        RECT 131.785 178.185 131.955 178.355 ;
        RECT 132.245 178.185 132.415 178.355 ;
        RECT 132.705 178.185 132.875 178.355 ;
        RECT 133.165 178.185 133.335 178.355 ;
        RECT 133.625 178.185 133.795 178.355 ;
        RECT 134.085 178.185 134.255 178.355 ;
        RECT 134.545 178.185 134.715 178.355 ;
        RECT 135.005 178.185 135.175 178.355 ;
        RECT 135.465 178.185 135.635 178.355 ;
        RECT 135.925 178.185 136.095 178.355 ;
        RECT 136.385 178.185 136.555 178.355 ;
        RECT 136.845 178.185 137.015 178.355 ;
        RECT 137.305 178.185 137.475 178.355 ;
        RECT 137.765 178.185 137.935 178.355 ;
        RECT 138.225 178.185 138.395 178.355 ;
        RECT 138.685 178.185 138.855 178.355 ;
        RECT 139.145 178.185 139.315 178.355 ;
        RECT 139.605 178.185 139.775 178.355 ;
        RECT 140.065 178.185 140.235 178.355 ;
        RECT 140.525 178.185 140.695 178.355 ;
        RECT 140.985 178.185 141.155 178.355 ;
        RECT 141.445 178.185 141.615 178.355 ;
        RECT 141.905 178.185 142.075 178.355 ;
        RECT 142.365 178.185 142.535 178.355 ;
        RECT 142.825 178.185 142.995 178.355 ;
        RECT 143.285 178.185 143.455 178.355 ;
        RECT 143.745 178.185 143.915 178.355 ;
        RECT 144.205 178.185 144.375 178.355 ;
        RECT 144.665 178.185 144.835 178.355 ;
        RECT 145.125 178.185 145.295 178.355 ;
        RECT 145.585 178.185 145.755 178.355 ;
        RECT 146.045 178.185 146.215 178.355 ;
        RECT 146.505 178.185 146.675 178.355 ;
        RECT 146.965 178.185 147.135 178.355 ;
        RECT 147.425 178.185 147.595 178.355 ;
        RECT 147.885 178.185 148.055 178.355 ;
        RECT 148.345 178.185 148.515 178.355 ;
        RECT 148.805 178.185 148.975 178.355 ;
        RECT 149.265 178.185 149.435 178.355 ;
        RECT 149.725 178.185 149.895 178.355 ;
        RECT 150.185 178.185 150.355 178.355 ;
        RECT 17.245 177.675 17.415 177.845 ;
        RECT 24.605 177.675 24.775 177.845 ;
        RECT 17.245 176.655 17.415 176.825 ;
        RECT 18.625 176.995 18.795 177.165 ;
        RECT 18.165 175.975 18.335 176.145 ;
        RECT 24.605 176.655 24.775 176.825 ;
        RECT 25.985 176.995 26.155 177.165 ;
        RECT 25.525 176.315 25.695 176.485 ;
        RECT 33.345 176.995 33.515 177.165 ;
        RECT 35.185 176.995 35.355 177.165 ;
        RECT 34.265 176.655 34.435 176.825 ;
        RECT 32.425 176.315 32.595 176.485 ;
        RECT 36.105 176.655 36.275 176.825 ;
        RECT 35.645 175.975 35.815 176.145 ;
        RECT 46.225 176.995 46.395 177.165 ;
        RECT 47.605 176.995 47.775 177.165 ;
        RECT 54.045 177.675 54.215 177.845 ;
        RECT 56.805 177.335 56.975 177.505 ;
        RECT 57.725 176.655 57.895 176.825 ;
        RECT 58.185 176.655 58.355 176.825 ;
        RECT 60.485 177.335 60.655 177.505 ;
        RECT 64.165 177.335 64.335 177.505 ;
        RECT 63.245 176.315 63.415 176.485 ;
        RECT 64.165 175.975 64.335 176.145 ;
        RECT 66.005 176.315 66.175 176.485 ;
        RECT 68.305 177.335 68.475 177.505 ;
        RECT 67.385 176.995 67.555 177.165 ;
        RECT 68.765 176.995 68.935 177.165 ;
        RECT 66.465 175.975 66.635 176.145 ;
        RECT 71.065 176.995 71.235 177.165 ;
        RECT 71.550 176.315 71.720 176.485 ;
        RECT 71.945 176.655 72.115 176.825 ;
        RECT 72.400 176.995 72.570 177.165 ;
        RECT 73.135 176.655 73.305 176.825 ;
        RECT 73.650 176.315 73.820 176.485 ;
        RECT 75.220 176.315 75.390 176.485 ;
        RECT 75.655 176.655 75.825 176.825 ;
        RECT 82.565 177.675 82.735 177.845 ;
        RECT 79.345 176.995 79.515 177.165 ;
        RECT 80.265 176.995 80.435 177.165 ;
        RECT 77.965 176.315 78.135 176.485 ;
        RECT 78.425 175.975 78.595 176.145 ;
        RECT 80.265 175.975 80.435 176.145 ;
        RECT 83.485 176.995 83.655 177.165 ;
        RECT 84.405 176.995 84.575 177.165 ;
        RECT 92.100 177.335 92.270 177.505 ;
        RECT 91.305 176.315 91.475 176.485 ;
        RECT 92.685 176.655 92.855 176.825 ;
        RECT 93.145 176.655 93.315 176.825 ;
        RECT 95.445 177.335 95.615 177.505 ;
        RECT 94.985 176.995 95.155 177.165 ;
        RECT 94.525 176.655 94.695 176.825 ;
        RECT 95.905 176.995 96.075 177.165 ;
        RECT 102.345 177.675 102.515 177.845 ;
        RECT 101.885 176.315 102.055 176.485 ;
        RECT 104.645 177.675 104.815 177.845 ;
        RECT 102.805 176.655 102.975 176.825 ;
        RECT 103.725 176.655 103.895 176.825 ;
        RECT 105.565 177.335 105.735 177.505 ;
        RECT 106.025 176.655 106.195 176.825 ;
        RECT 108.330 177.335 108.500 177.505 ;
        RECT 108.915 176.995 109.085 177.165 ;
        RECT 109.705 176.995 109.875 177.165 ;
        RECT 122.125 177.675 122.295 177.845 ;
        RECT 106.485 176.315 106.655 176.485 ;
        RECT 117.525 176.995 117.695 177.165 ;
        RECT 118.445 176.995 118.615 177.165 ;
        RECT 117.525 175.975 117.695 176.145 ;
        RECT 123.965 176.995 124.135 177.165 ;
        RECT 124.425 176.995 124.595 177.165 ;
        RECT 125.345 175.975 125.515 176.145 ;
        RECT 11.265 175.465 11.435 175.635 ;
        RECT 11.725 175.465 11.895 175.635 ;
        RECT 12.185 175.465 12.355 175.635 ;
        RECT 12.645 175.465 12.815 175.635 ;
        RECT 13.105 175.465 13.275 175.635 ;
        RECT 13.565 175.465 13.735 175.635 ;
        RECT 14.025 175.465 14.195 175.635 ;
        RECT 14.485 175.465 14.655 175.635 ;
        RECT 14.945 175.465 15.115 175.635 ;
        RECT 15.405 175.465 15.575 175.635 ;
        RECT 15.865 175.465 16.035 175.635 ;
        RECT 16.325 175.465 16.495 175.635 ;
        RECT 16.785 175.465 16.955 175.635 ;
        RECT 17.245 175.465 17.415 175.635 ;
        RECT 17.705 175.465 17.875 175.635 ;
        RECT 18.165 175.465 18.335 175.635 ;
        RECT 18.625 175.465 18.795 175.635 ;
        RECT 19.085 175.465 19.255 175.635 ;
        RECT 19.545 175.465 19.715 175.635 ;
        RECT 20.005 175.465 20.175 175.635 ;
        RECT 20.465 175.465 20.635 175.635 ;
        RECT 20.925 175.465 21.095 175.635 ;
        RECT 21.385 175.465 21.555 175.635 ;
        RECT 21.845 175.465 22.015 175.635 ;
        RECT 22.305 175.465 22.475 175.635 ;
        RECT 22.765 175.465 22.935 175.635 ;
        RECT 23.225 175.465 23.395 175.635 ;
        RECT 23.685 175.465 23.855 175.635 ;
        RECT 24.145 175.465 24.315 175.635 ;
        RECT 24.605 175.465 24.775 175.635 ;
        RECT 25.065 175.465 25.235 175.635 ;
        RECT 25.525 175.465 25.695 175.635 ;
        RECT 25.985 175.465 26.155 175.635 ;
        RECT 26.445 175.465 26.615 175.635 ;
        RECT 26.905 175.465 27.075 175.635 ;
        RECT 27.365 175.465 27.535 175.635 ;
        RECT 27.825 175.465 27.995 175.635 ;
        RECT 28.285 175.465 28.455 175.635 ;
        RECT 28.745 175.465 28.915 175.635 ;
        RECT 29.205 175.465 29.375 175.635 ;
        RECT 29.665 175.465 29.835 175.635 ;
        RECT 30.125 175.465 30.295 175.635 ;
        RECT 30.585 175.465 30.755 175.635 ;
        RECT 31.045 175.465 31.215 175.635 ;
        RECT 31.505 175.465 31.675 175.635 ;
        RECT 31.965 175.465 32.135 175.635 ;
        RECT 32.425 175.465 32.595 175.635 ;
        RECT 32.885 175.465 33.055 175.635 ;
        RECT 33.345 175.465 33.515 175.635 ;
        RECT 33.805 175.465 33.975 175.635 ;
        RECT 34.265 175.465 34.435 175.635 ;
        RECT 34.725 175.465 34.895 175.635 ;
        RECT 35.185 175.465 35.355 175.635 ;
        RECT 35.645 175.465 35.815 175.635 ;
        RECT 36.105 175.465 36.275 175.635 ;
        RECT 36.565 175.465 36.735 175.635 ;
        RECT 37.025 175.465 37.195 175.635 ;
        RECT 37.485 175.465 37.655 175.635 ;
        RECT 37.945 175.465 38.115 175.635 ;
        RECT 38.405 175.465 38.575 175.635 ;
        RECT 38.865 175.465 39.035 175.635 ;
        RECT 39.325 175.465 39.495 175.635 ;
        RECT 39.785 175.465 39.955 175.635 ;
        RECT 40.245 175.465 40.415 175.635 ;
        RECT 40.705 175.465 40.875 175.635 ;
        RECT 41.165 175.465 41.335 175.635 ;
        RECT 41.625 175.465 41.795 175.635 ;
        RECT 42.085 175.465 42.255 175.635 ;
        RECT 42.545 175.465 42.715 175.635 ;
        RECT 43.005 175.465 43.175 175.635 ;
        RECT 43.465 175.465 43.635 175.635 ;
        RECT 43.925 175.465 44.095 175.635 ;
        RECT 44.385 175.465 44.555 175.635 ;
        RECT 44.845 175.465 45.015 175.635 ;
        RECT 45.305 175.465 45.475 175.635 ;
        RECT 45.765 175.465 45.935 175.635 ;
        RECT 46.225 175.465 46.395 175.635 ;
        RECT 46.685 175.465 46.855 175.635 ;
        RECT 47.145 175.465 47.315 175.635 ;
        RECT 47.605 175.465 47.775 175.635 ;
        RECT 48.065 175.465 48.235 175.635 ;
        RECT 48.525 175.465 48.695 175.635 ;
        RECT 48.985 175.465 49.155 175.635 ;
        RECT 49.445 175.465 49.615 175.635 ;
        RECT 49.905 175.465 50.075 175.635 ;
        RECT 50.365 175.465 50.535 175.635 ;
        RECT 50.825 175.465 50.995 175.635 ;
        RECT 51.285 175.465 51.455 175.635 ;
        RECT 51.745 175.465 51.915 175.635 ;
        RECT 52.205 175.465 52.375 175.635 ;
        RECT 52.665 175.465 52.835 175.635 ;
        RECT 53.125 175.465 53.295 175.635 ;
        RECT 53.585 175.465 53.755 175.635 ;
        RECT 54.045 175.465 54.215 175.635 ;
        RECT 54.505 175.465 54.675 175.635 ;
        RECT 54.965 175.465 55.135 175.635 ;
        RECT 55.425 175.465 55.595 175.635 ;
        RECT 55.885 175.465 56.055 175.635 ;
        RECT 56.345 175.465 56.515 175.635 ;
        RECT 56.805 175.465 56.975 175.635 ;
        RECT 57.265 175.465 57.435 175.635 ;
        RECT 57.725 175.465 57.895 175.635 ;
        RECT 58.185 175.465 58.355 175.635 ;
        RECT 58.645 175.465 58.815 175.635 ;
        RECT 59.105 175.465 59.275 175.635 ;
        RECT 59.565 175.465 59.735 175.635 ;
        RECT 60.025 175.465 60.195 175.635 ;
        RECT 60.485 175.465 60.655 175.635 ;
        RECT 60.945 175.465 61.115 175.635 ;
        RECT 61.405 175.465 61.575 175.635 ;
        RECT 61.865 175.465 62.035 175.635 ;
        RECT 62.325 175.465 62.495 175.635 ;
        RECT 62.785 175.465 62.955 175.635 ;
        RECT 63.245 175.465 63.415 175.635 ;
        RECT 63.705 175.465 63.875 175.635 ;
        RECT 64.165 175.465 64.335 175.635 ;
        RECT 64.625 175.465 64.795 175.635 ;
        RECT 65.085 175.465 65.255 175.635 ;
        RECT 65.545 175.465 65.715 175.635 ;
        RECT 66.005 175.465 66.175 175.635 ;
        RECT 66.465 175.465 66.635 175.635 ;
        RECT 66.925 175.465 67.095 175.635 ;
        RECT 67.385 175.465 67.555 175.635 ;
        RECT 67.845 175.465 68.015 175.635 ;
        RECT 68.305 175.465 68.475 175.635 ;
        RECT 68.765 175.465 68.935 175.635 ;
        RECT 69.225 175.465 69.395 175.635 ;
        RECT 69.685 175.465 69.855 175.635 ;
        RECT 70.145 175.465 70.315 175.635 ;
        RECT 70.605 175.465 70.775 175.635 ;
        RECT 71.065 175.465 71.235 175.635 ;
        RECT 71.525 175.465 71.695 175.635 ;
        RECT 71.985 175.465 72.155 175.635 ;
        RECT 72.445 175.465 72.615 175.635 ;
        RECT 72.905 175.465 73.075 175.635 ;
        RECT 73.365 175.465 73.535 175.635 ;
        RECT 73.825 175.465 73.995 175.635 ;
        RECT 74.285 175.465 74.455 175.635 ;
        RECT 74.745 175.465 74.915 175.635 ;
        RECT 75.205 175.465 75.375 175.635 ;
        RECT 75.665 175.465 75.835 175.635 ;
        RECT 76.125 175.465 76.295 175.635 ;
        RECT 76.585 175.465 76.755 175.635 ;
        RECT 77.045 175.465 77.215 175.635 ;
        RECT 77.505 175.465 77.675 175.635 ;
        RECT 77.965 175.465 78.135 175.635 ;
        RECT 78.425 175.465 78.595 175.635 ;
        RECT 78.885 175.465 79.055 175.635 ;
        RECT 79.345 175.465 79.515 175.635 ;
        RECT 79.805 175.465 79.975 175.635 ;
        RECT 80.265 175.465 80.435 175.635 ;
        RECT 80.725 175.465 80.895 175.635 ;
        RECT 81.185 175.465 81.355 175.635 ;
        RECT 81.645 175.465 81.815 175.635 ;
        RECT 82.105 175.465 82.275 175.635 ;
        RECT 82.565 175.465 82.735 175.635 ;
        RECT 83.025 175.465 83.195 175.635 ;
        RECT 83.485 175.465 83.655 175.635 ;
        RECT 83.945 175.465 84.115 175.635 ;
        RECT 84.405 175.465 84.575 175.635 ;
        RECT 84.865 175.465 85.035 175.635 ;
        RECT 85.325 175.465 85.495 175.635 ;
        RECT 85.785 175.465 85.955 175.635 ;
        RECT 86.245 175.465 86.415 175.635 ;
        RECT 86.705 175.465 86.875 175.635 ;
        RECT 87.165 175.465 87.335 175.635 ;
        RECT 87.625 175.465 87.795 175.635 ;
        RECT 88.085 175.465 88.255 175.635 ;
        RECT 88.545 175.465 88.715 175.635 ;
        RECT 89.005 175.465 89.175 175.635 ;
        RECT 89.465 175.465 89.635 175.635 ;
        RECT 89.925 175.465 90.095 175.635 ;
        RECT 90.385 175.465 90.555 175.635 ;
        RECT 90.845 175.465 91.015 175.635 ;
        RECT 91.305 175.465 91.475 175.635 ;
        RECT 91.765 175.465 91.935 175.635 ;
        RECT 92.225 175.465 92.395 175.635 ;
        RECT 92.685 175.465 92.855 175.635 ;
        RECT 93.145 175.465 93.315 175.635 ;
        RECT 93.605 175.465 93.775 175.635 ;
        RECT 94.065 175.465 94.235 175.635 ;
        RECT 94.525 175.465 94.695 175.635 ;
        RECT 94.985 175.465 95.155 175.635 ;
        RECT 95.445 175.465 95.615 175.635 ;
        RECT 95.905 175.465 96.075 175.635 ;
        RECT 96.365 175.465 96.535 175.635 ;
        RECT 96.825 175.465 96.995 175.635 ;
        RECT 97.285 175.465 97.455 175.635 ;
        RECT 97.745 175.465 97.915 175.635 ;
        RECT 98.205 175.465 98.375 175.635 ;
        RECT 98.665 175.465 98.835 175.635 ;
        RECT 99.125 175.465 99.295 175.635 ;
        RECT 99.585 175.465 99.755 175.635 ;
        RECT 100.045 175.465 100.215 175.635 ;
        RECT 100.505 175.465 100.675 175.635 ;
        RECT 100.965 175.465 101.135 175.635 ;
        RECT 101.425 175.465 101.595 175.635 ;
        RECT 101.885 175.465 102.055 175.635 ;
        RECT 102.345 175.465 102.515 175.635 ;
        RECT 102.805 175.465 102.975 175.635 ;
        RECT 103.265 175.465 103.435 175.635 ;
        RECT 103.725 175.465 103.895 175.635 ;
        RECT 104.185 175.465 104.355 175.635 ;
        RECT 104.645 175.465 104.815 175.635 ;
        RECT 105.105 175.465 105.275 175.635 ;
        RECT 105.565 175.465 105.735 175.635 ;
        RECT 106.025 175.465 106.195 175.635 ;
        RECT 106.485 175.465 106.655 175.635 ;
        RECT 106.945 175.465 107.115 175.635 ;
        RECT 107.405 175.465 107.575 175.635 ;
        RECT 107.865 175.465 108.035 175.635 ;
        RECT 108.325 175.465 108.495 175.635 ;
        RECT 108.785 175.465 108.955 175.635 ;
        RECT 109.245 175.465 109.415 175.635 ;
        RECT 109.705 175.465 109.875 175.635 ;
        RECT 110.165 175.465 110.335 175.635 ;
        RECT 110.625 175.465 110.795 175.635 ;
        RECT 111.085 175.465 111.255 175.635 ;
        RECT 111.545 175.465 111.715 175.635 ;
        RECT 112.005 175.465 112.175 175.635 ;
        RECT 112.465 175.465 112.635 175.635 ;
        RECT 112.925 175.465 113.095 175.635 ;
        RECT 113.385 175.465 113.555 175.635 ;
        RECT 113.845 175.465 114.015 175.635 ;
        RECT 114.305 175.465 114.475 175.635 ;
        RECT 114.765 175.465 114.935 175.635 ;
        RECT 115.225 175.465 115.395 175.635 ;
        RECT 115.685 175.465 115.855 175.635 ;
        RECT 116.145 175.465 116.315 175.635 ;
        RECT 116.605 175.465 116.775 175.635 ;
        RECT 117.065 175.465 117.235 175.635 ;
        RECT 117.525 175.465 117.695 175.635 ;
        RECT 117.985 175.465 118.155 175.635 ;
        RECT 118.445 175.465 118.615 175.635 ;
        RECT 118.905 175.465 119.075 175.635 ;
        RECT 119.365 175.465 119.535 175.635 ;
        RECT 119.825 175.465 119.995 175.635 ;
        RECT 120.285 175.465 120.455 175.635 ;
        RECT 120.745 175.465 120.915 175.635 ;
        RECT 121.205 175.465 121.375 175.635 ;
        RECT 121.665 175.465 121.835 175.635 ;
        RECT 122.125 175.465 122.295 175.635 ;
        RECT 122.585 175.465 122.755 175.635 ;
        RECT 123.045 175.465 123.215 175.635 ;
        RECT 123.505 175.465 123.675 175.635 ;
        RECT 123.965 175.465 124.135 175.635 ;
        RECT 124.425 175.465 124.595 175.635 ;
        RECT 124.885 175.465 125.055 175.635 ;
        RECT 125.345 175.465 125.515 175.635 ;
        RECT 125.805 175.465 125.975 175.635 ;
        RECT 126.265 175.465 126.435 175.635 ;
        RECT 126.725 175.465 126.895 175.635 ;
        RECT 127.185 175.465 127.355 175.635 ;
        RECT 127.645 175.465 127.815 175.635 ;
        RECT 128.105 175.465 128.275 175.635 ;
        RECT 128.565 175.465 128.735 175.635 ;
        RECT 129.025 175.465 129.195 175.635 ;
        RECT 129.485 175.465 129.655 175.635 ;
        RECT 129.945 175.465 130.115 175.635 ;
        RECT 130.405 175.465 130.575 175.635 ;
        RECT 130.865 175.465 131.035 175.635 ;
        RECT 131.325 175.465 131.495 175.635 ;
        RECT 131.785 175.465 131.955 175.635 ;
        RECT 132.245 175.465 132.415 175.635 ;
        RECT 132.705 175.465 132.875 175.635 ;
        RECT 133.165 175.465 133.335 175.635 ;
        RECT 133.625 175.465 133.795 175.635 ;
        RECT 134.085 175.465 134.255 175.635 ;
        RECT 134.545 175.465 134.715 175.635 ;
        RECT 135.005 175.465 135.175 175.635 ;
        RECT 135.465 175.465 135.635 175.635 ;
        RECT 135.925 175.465 136.095 175.635 ;
        RECT 136.385 175.465 136.555 175.635 ;
        RECT 136.845 175.465 137.015 175.635 ;
        RECT 137.305 175.465 137.475 175.635 ;
        RECT 137.765 175.465 137.935 175.635 ;
        RECT 138.225 175.465 138.395 175.635 ;
        RECT 138.685 175.465 138.855 175.635 ;
        RECT 139.145 175.465 139.315 175.635 ;
        RECT 139.605 175.465 139.775 175.635 ;
        RECT 140.065 175.465 140.235 175.635 ;
        RECT 140.525 175.465 140.695 175.635 ;
        RECT 140.985 175.465 141.155 175.635 ;
        RECT 141.445 175.465 141.615 175.635 ;
        RECT 141.905 175.465 142.075 175.635 ;
        RECT 142.365 175.465 142.535 175.635 ;
        RECT 142.825 175.465 142.995 175.635 ;
        RECT 143.285 175.465 143.455 175.635 ;
        RECT 143.745 175.465 143.915 175.635 ;
        RECT 144.205 175.465 144.375 175.635 ;
        RECT 144.665 175.465 144.835 175.635 ;
        RECT 145.125 175.465 145.295 175.635 ;
        RECT 145.585 175.465 145.755 175.635 ;
        RECT 146.045 175.465 146.215 175.635 ;
        RECT 146.505 175.465 146.675 175.635 ;
        RECT 146.965 175.465 147.135 175.635 ;
        RECT 147.425 175.465 147.595 175.635 ;
        RECT 147.885 175.465 148.055 175.635 ;
        RECT 148.345 175.465 148.515 175.635 ;
        RECT 148.805 175.465 148.975 175.635 ;
        RECT 149.265 175.465 149.435 175.635 ;
        RECT 149.725 175.465 149.895 175.635 ;
        RECT 150.185 175.465 150.355 175.635 ;
        RECT 17.245 173.935 17.415 174.105 ;
        RECT 16.325 173.255 16.495 173.425 ;
        RECT 37.485 174.955 37.655 175.125 ;
        RECT 37.485 173.935 37.655 174.105 ;
        RECT 38.405 173.935 38.575 174.105 ;
        RECT 42.085 174.615 42.255 174.785 ;
        RECT 43.005 173.935 43.175 174.105 ;
        RECT 43.465 173.255 43.635 173.425 ;
        RECT 43.925 173.935 44.095 174.105 ;
        RECT 44.845 173.595 45.015 173.765 ;
        RECT 52.205 174.955 52.375 175.125 ;
        RECT 50.365 174.275 50.535 174.445 ;
        RECT 51.285 173.935 51.455 174.105 ;
        RECT 55.425 174.955 55.595 175.125 ;
        RECT 55.885 174.955 56.055 175.125 ;
        RECT 53.585 173.935 53.755 174.105 ;
        RECT 54.505 173.935 54.675 174.105 ;
        RECT 54.965 173.935 55.135 174.105 ;
        RECT 56.345 174.275 56.515 174.445 ;
        RECT 53.125 173.255 53.295 173.425 ;
        RECT 64.165 173.935 64.335 174.105 ;
        RECT 65.085 173.255 65.255 173.425 ;
        RECT 67.385 174.955 67.555 175.125 ;
        RECT 68.305 173.935 68.475 174.105 ;
        RECT 68.765 173.595 68.935 173.765 ;
        RECT 70.145 173.935 70.315 174.105 ;
        RECT 69.225 173.595 69.395 173.765 ;
        RECT 72.445 174.955 72.615 175.125 ;
        RECT 72.445 173.595 72.615 173.765 ;
        RECT 73.825 173.935 73.995 174.105 ;
        RECT 76.125 173.935 76.295 174.105 ;
        RECT 76.585 173.935 76.755 174.105 ;
        RECT 77.505 174.275 77.675 174.445 ;
        RECT 73.365 173.255 73.535 173.425 ;
        RECT 77.505 173.595 77.675 173.765 ;
        RECT 82.565 173.255 82.735 173.425 ;
        RECT 85.325 174.275 85.495 174.445 ;
        RECT 89.925 174.955 90.095 175.125 ;
        RECT 92.225 174.275 92.395 174.445 ;
        RECT 93.145 174.275 93.315 174.445 ;
        RECT 100.045 173.595 100.215 173.765 ;
        RECT 98.665 173.255 98.835 173.425 ;
        RECT 101.885 173.935 102.055 174.105 ;
        RECT 102.345 173.595 102.515 173.765 ;
        RECT 109.245 174.955 109.415 175.125 ;
        RECT 112.925 174.955 113.095 175.125 ;
        RECT 110.165 173.935 110.335 174.105 ;
        RECT 110.625 174.275 110.795 174.445 ;
        RECT 111.085 173.935 111.255 174.105 ;
        RECT 111.545 174.275 111.715 174.445 ;
        RECT 112.465 174.275 112.635 174.445 ;
        RECT 113.385 173.935 113.555 174.105 ;
        RECT 113.845 173.935 114.015 174.105 ;
        RECT 119.365 174.955 119.535 175.125 ;
        RECT 116.605 173.935 116.775 174.105 ;
        RECT 117.065 173.935 117.235 174.105 ;
        RECT 118.905 173.935 119.075 174.105 ;
        RECT 120.285 174.275 120.455 174.445 ;
        RECT 115.685 173.595 115.855 173.765 ;
        RECT 120.745 173.935 120.915 174.105 ;
        RECT 120.285 173.595 120.455 173.765 ;
        RECT 121.665 173.595 121.835 173.765 ;
        RECT 122.585 173.935 122.755 174.105 ;
        RECT 122.125 173.595 122.295 173.765 ;
        RECT 123.505 173.255 123.675 173.425 ;
        RECT 11.265 172.745 11.435 172.915 ;
        RECT 11.725 172.745 11.895 172.915 ;
        RECT 12.185 172.745 12.355 172.915 ;
        RECT 12.645 172.745 12.815 172.915 ;
        RECT 13.105 172.745 13.275 172.915 ;
        RECT 13.565 172.745 13.735 172.915 ;
        RECT 14.025 172.745 14.195 172.915 ;
        RECT 14.485 172.745 14.655 172.915 ;
        RECT 14.945 172.745 15.115 172.915 ;
        RECT 15.405 172.745 15.575 172.915 ;
        RECT 15.865 172.745 16.035 172.915 ;
        RECT 16.325 172.745 16.495 172.915 ;
        RECT 16.785 172.745 16.955 172.915 ;
        RECT 17.245 172.745 17.415 172.915 ;
        RECT 17.705 172.745 17.875 172.915 ;
        RECT 18.165 172.745 18.335 172.915 ;
        RECT 18.625 172.745 18.795 172.915 ;
        RECT 19.085 172.745 19.255 172.915 ;
        RECT 19.545 172.745 19.715 172.915 ;
        RECT 20.005 172.745 20.175 172.915 ;
        RECT 20.465 172.745 20.635 172.915 ;
        RECT 20.925 172.745 21.095 172.915 ;
        RECT 21.385 172.745 21.555 172.915 ;
        RECT 21.845 172.745 22.015 172.915 ;
        RECT 22.305 172.745 22.475 172.915 ;
        RECT 22.765 172.745 22.935 172.915 ;
        RECT 23.225 172.745 23.395 172.915 ;
        RECT 23.685 172.745 23.855 172.915 ;
        RECT 24.145 172.745 24.315 172.915 ;
        RECT 24.605 172.745 24.775 172.915 ;
        RECT 25.065 172.745 25.235 172.915 ;
        RECT 25.525 172.745 25.695 172.915 ;
        RECT 25.985 172.745 26.155 172.915 ;
        RECT 26.445 172.745 26.615 172.915 ;
        RECT 26.905 172.745 27.075 172.915 ;
        RECT 27.365 172.745 27.535 172.915 ;
        RECT 27.825 172.745 27.995 172.915 ;
        RECT 28.285 172.745 28.455 172.915 ;
        RECT 28.745 172.745 28.915 172.915 ;
        RECT 29.205 172.745 29.375 172.915 ;
        RECT 29.665 172.745 29.835 172.915 ;
        RECT 30.125 172.745 30.295 172.915 ;
        RECT 30.585 172.745 30.755 172.915 ;
        RECT 31.045 172.745 31.215 172.915 ;
        RECT 31.505 172.745 31.675 172.915 ;
        RECT 31.965 172.745 32.135 172.915 ;
        RECT 32.425 172.745 32.595 172.915 ;
        RECT 32.885 172.745 33.055 172.915 ;
        RECT 33.345 172.745 33.515 172.915 ;
        RECT 33.805 172.745 33.975 172.915 ;
        RECT 34.265 172.745 34.435 172.915 ;
        RECT 34.725 172.745 34.895 172.915 ;
        RECT 35.185 172.745 35.355 172.915 ;
        RECT 35.645 172.745 35.815 172.915 ;
        RECT 36.105 172.745 36.275 172.915 ;
        RECT 36.565 172.745 36.735 172.915 ;
        RECT 37.025 172.745 37.195 172.915 ;
        RECT 37.485 172.745 37.655 172.915 ;
        RECT 37.945 172.745 38.115 172.915 ;
        RECT 38.405 172.745 38.575 172.915 ;
        RECT 38.865 172.745 39.035 172.915 ;
        RECT 39.325 172.745 39.495 172.915 ;
        RECT 39.785 172.745 39.955 172.915 ;
        RECT 40.245 172.745 40.415 172.915 ;
        RECT 40.705 172.745 40.875 172.915 ;
        RECT 41.165 172.745 41.335 172.915 ;
        RECT 41.625 172.745 41.795 172.915 ;
        RECT 42.085 172.745 42.255 172.915 ;
        RECT 42.545 172.745 42.715 172.915 ;
        RECT 43.005 172.745 43.175 172.915 ;
        RECT 43.465 172.745 43.635 172.915 ;
        RECT 43.925 172.745 44.095 172.915 ;
        RECT 44.385 172.745 44.555 172.915 ;
        RECT 44.845 172.745 45.015 172.915 ;
        RECT 45.305 172.745 45.475 172.915 ;
        RECT 45.765 172.745 45.935 172.915 ;
        RECT 46.225 172.745 46.395 172.915 ;
        RECT 46.685 172.745 46.855 172.915 ;
        RECT 47.145 172.745 47.315 172.915 ;
        RECT 47.605 172.745 47.775 172.915 ;
        RECT 48.065 172.745 48.235 172.915 ;
        RECT 48.525 172.745 48.695 172.915 ;
        RECT 48.985 172.745 49.155 172.915 ;
        RECT 49.445 172.745 49.615 172.915 ;
        RECT 49.905 172.745 50.075 172.915 ;
        RECT 50.365 172.745 50.535 172.915 ;
        RECT 50.825 172.745 50.995 172.915 ;
        RECT 51.285 172.745 51.455 172.915 ;
        RECT 51.745 172.745 51.915 172.915 ;
        RECT 52.205 172.745 52.375 172.915 ;
        RECT 52.665 172.745 52.835 172.915 ;
        RECT 53.125 172.745 53.295 172.915 ;
        RECT 53.585 172.745 53.755 172.915 ;
        RECT 54.045 172.745 54.215 172.915 ;
        RECT 54.505 172.745 54.675 172.915 ;
        RECT 54.965 172.745 55.135 172.915 ;
        RECT 55.425 172.745 55.595 172.915 ;
        RECT 55.885 172.745 56.055 172.915 ;
        RECT 56.345 172.745 56.515 172.915 ;
        RECT 56.805 172.745 56.975 172.915 ;
        RECT 57.265 172.745 57.435 172.915 ;
        RECT 57.725 172.745 57.895 172.915 ;
        RECT 58.185 172.745 58.355 172.915 ;
        RECT 58.645 172.745 58.815 172.915 ;
        RECT 59.105 172.745 59.275 172.915 ;
        RECT 59.565 172.745 59.735 172.915 ;
        RECT 60.025 172.745 60.195 172.915 ;
        RECT 60.485 172.745 60.655 172.915 ;
        RECT 60.945 172.745 61.115 172.915 ;
        RECT 61.405 172.745 61.575 172.915 ;
        RECT 61.865 172.745 62.035 172.915 ;
        RECT 62.325 172.745 62.495 172.915 ;
        RECT 62.785 172.745 62.955 172.915 ;
        RECT 63.245 172.745 63.415 172.915 ;
        RECT 63.705 172.745 63.875 172.915 ;
        RECT 64.165 172.745 64.335 172.915 ;
        RECT 64.625 172.745 64.795 172.915 ;
        RECT 65.085 172.745 65.255 172.915 ;
        RECT 65.545 172.745 65.715 172.915 ;
        RECT 66.005 172.745 66.175 172.915 ;
        RECT 66.465 172.745 66.635 172.915 ;
        RECT 66.925 172.745 67.095 172.915 ;
        RECT 67.385 172.745 67.555 172.915 ;
        RECT 67.845 172.745 68.015 172.915 ;
        RECT 68.305 172.745 68.475 172.915 ;
        RECT 68.765 172.745 68.935 172.915 ;
        RECT 69.225 172.745 69.395 172.915 ;
        RECT 69.685 172.745 69.855 172.915 ;
        RECT 70.145 172.745 70.315 172.915 ;
        RECT 70.605 172.745 70.775 172.915 ;
        RECT 71.065 172.745 71.235 172.915 ;
        RECT 71.525 172.745 71.695 172.915 ;
        RECT 71.985 172.745 72.155 172.915 ;
        RECT 72.445 172.745 72.615 172.915 ;
        RECT 72.905 172.745 73.075 172.915 ;
        RECT 73.365 172.745 73.535 172.915 ;
        RECT 73.825 172.745 73.995 172.915 ;
        RECT 74.285 172.745 74.455 172.915 ;
        RECT 74.745 172.745 74.915 172.915 ;
        RECT 75.205 172.745 75.375 172.915 ;
        RECT 75.665 172.745 75.835 172.915 ;
        RECT 76.125 172.745 76.295 172.915 ;
        RECT 76.585 172.745 76.755 172.915 ;
        RECT 77.045 172.745 77.215 172.915 ;
        RECT 77.505 172.745 77.675 172.915 ;
        RECT 77.965 172.745 78.135 172.915 ;
        RECT 78.425 172.745 78.595 172.915 ;
        RECT 78.885 172.745 79.055 172.915 ;
        RECT 79.345 172.745 79.515 172.915 ;
        RECT 79.805 172.745 79.975 172.915 ;
        RECT 80.265 172.745 80.435 172.915 ;
        RECT 80.725 172.745 80.895 172.915 ;
        RECT 81.185 172.745 81.355 172.915 ;
        RECT 81.645 172.745 81.815 172.915 ;
        RECT 82.105 172.745 82.275 172.915 ;
        RECT 82.565 172.745 82.735 172.915 ;
        RECT 83.025 172.745 83.195 172.915 ;
        RECT 83.485 172.745 83.655 172.915 ;
        RECT 83.945 172.745 84.115 172.915 ;
        RECT 84.405 172.745 84.575 172.915 ;
        RECT 84.865 172.745 85.035 172.915 ;
        RECT 85.325 172.745 85.495 172.915 ;
        RECT 85.785 172.745 85.955 172.915 ;
        RECT 86.245 172.745 86.415 172.915 ;
        RECT 86.705 172.745 86.875 172.915 ;
        RECT 87.165 172.745 87.335 172.915 ;
        RECT 87.625 172.745 87.795 172.915 ;
        RECT 88.085 172.745 88.255 172.915 ;
        RECT 88.545 172.745 88.715 172.915 ;
        RECT 89.005 172.745 89.175 172.915 ;
        RECT 89.465 172.745 89.635 172.915 ;
        RECT 89.925 172.745 90.095 172.915 ;
        RECT 90.385 172.745 90.555 172.915 ;
        RECT 90.845 172.745 91.015 172.915 ;
        RECT 91.305 172.745 91.475 172.915 ;
        RECT 91.765 172.745 91.935 172.915 ;
        RECT 92.225 172.745 92.395 172.915 ;
        RECT 92.685 172.745 92.855 172.915 ;
        RECT 93.145 172.745 93.315 172.915 ;
        RECT 93.605 172.745 93.775 172.915 ;
        RECT 94.065 172.745 94.235 172.915 ;
        RECT 94.525 172.745 94.695 172.915 ;
        RECT 94.985 172.745 95.155 172.915 ;
        RECT 95.445 172.745 95.615 172.915 ;
        RECT 95.905 172.745 96.075 172.915 ;
        RECT 96.365 172.745 96.535 172.915 ;
        RECT 96.825 172.745 96.995 172.915 ;
        RECT 97.285 172.745 97.455 172.915 ;
        RECT 97.745 172.745 97.915 172.915 ;
        RECT 98.205 172.745 98.375 172.915 ;
        RECT 98.665 172.745 98.835 172.915 ;
        RECT 99.125 172.745 99.295 172.915 ;
        RECT 99.585 172.745 99.755 172.915 ;
        RECT 100.045 172.745 100.215 172.915 ;
        RECT 100.505 172.745 100.675 172.915 ;
        RECT 100.965 172.745 101.135 172.915 ;
        RECT 101.425 172.745 101.595 172.915 ;
        RECT 101.885 172.745 102.055 172.915 ;
        RECT 102.345 172.745 102.515 172.915 ;
        RECT 102.805 172.745 102.975 172.915 ;
        RECT 103.265 172.745 103.435 172.915 ;
        RECT 103.725 172.745 103.895 172.915 ;
        RECT 104.185 172.745 104.355 172.915 ;
        RECT 104.645 172.745 104.815 172.915 ;
        RECT 105.105 172.745 105.275 172.915 ;
        RECT 105.565 172.745 105.735 172.915 ;
        RECT 106.025 172.745 106.195 172.915 ;
        RECT 106.485 172.745 106.655 172.915 ;
        RECT 106.945 172.745 107.115 172.915 ;
        RECT 107.405 172.745 107.575 172.915 ;
        RECT 107.865 172.745 108.035 172.915 ;
        RECT 108.325 172.745 108.495 172.915 ;
        RECT 108.785 172.745 108.955 172.915 ;
        RECT 109.245 172.745 109.415 172.915 ;
        RECT 109.705 172.745 109.875 172.915 ;
        RECT 110.165 172.745 110.335 172.915 ;
        RECT 110.625 172.745 110.795 172.915 ;
        RECT 111.085 172.745 111.255 172.915 ;
        RECT 111.545 172.745 111.715 172.915 ;
        RECT 112.005 172.745 112.175 172.915 ;
        RECT 112.465 172.745 112.635 172.915 ;
        RECT 112.925 172.745 113.095 172.915 ;
        RECT 113.385 172.745 113.555 172.915 ;
        RECT 113.845 172.745 114.015 172.915 ;
        RECT 114.305 172.745 114.475 172.915 ;
        RECT 114.765 172.745 114.935 172.915 ;
        RECT 115.225 172.745 115.395 172.915 ;
        RECT 115.685 172.745 115.855 172.915 ;
        RECT 116.145 172.745 116.315 172.915 ;
        RECT 116.605 172.745 116.775 172.915 ;
        RECT 117.065 172.745 117.235 172.915 ;
        RECT 117.525 172.745 117.695 172.915 ;
        RECT 117.985 172.745 118.155 172.915 ;
        RECT 118.445 172.745 118.615 172.915 ;
        RECT 118.905 172.745 119.075 172.915 ;
        RECT 119.365 172.745 119.535 172.915 ;
        RECT 119.825 172.745 119.995 172.915 ;
        RECT 120.285 172.745 120.455 172.915 ;
        RECT 120.745 172.745 120.915 172.915 ;
        RECT 121.205 172.745 121.375 172.915 ;
        RECT 121.665 172.745 121.835 172.915 ;
        RECT 122.125 172.745 122.295 172.915 ;
        RECT 122.585 172.745 122.755 172.915 ;
        RECT 123.045 172.745 123.215 172.915 ;
        RECT 123.505 172.745 123.675 172.915 ;
        RECT 123.965 172.745 124.135 172.915 ;
        RECT 124.425 172.745 124.595 172.915 ;
        RECT 124.885 172.745 125.055 172.915 ;
        RECT 125.345 172.745 125.515 172.915 ;
        RECT 125.805 172.745 125.975 172.915 ;
        RECT 126.265 172.745 126.435 172.915 ;
        RECT 126.725 172.745 126.895 172.915 ;
        RECT 127.185 172.745 127.355 172.915 ;
        RECT 127.645 172.745 127.815 172.915 ;
        RECT 128.105 172.745 128.275 172.915 ;
        RECT 128.565 172.745 128.735 172.915 ;
        RECT 129.025 172.745 129.195 172.915 ;
        RECT 129.485 172.745 129.655 172.915 ;
        RECT 129.945 172.745 130.115 172.915 ;
        RECT 130.405 172.745 130.575 172.915 ;
        RECT 130.865 172.745 131.035 172.915 ;
        RECT 131.325 172.745 131.495 172.915 ;
        RECT 131.785 172.745 131.955 172.915 ;
        RECT 132.245 172.745 132.415 172.915 ;
        RECT 132.705 172.745 132.875 172.915 ;
        RECT 133.165 172.745 133.335 172.915 ;
        RECT 133.625 172.745 133.795 172.915 ;
        RECT 134.085 172.745 134.255 172.915 ;
        RECT 134.545 172.745 134.715 172.915 ;
        RECT 135.005 172.745 135.175 172.915 ;
        RECT 135.465 172.745 135.635 172.915 ;
        RECT 135.925 172.745 136.095 172.915 ;
        RECT 136.385 172.745 136.555 172.915 ;
        RECT 136.845 172.745 137.015 172.915 ;
        RECT 137.305 172.745 137.475 172.915 ;
        RECT 137.765 172.745 137.935 172.915 ;
        RECT 138.225 172.745 138.395 172.915 ;
        RECT 138.685 172.745 138.855 172.915 ;
        RECT 139.145 172.745 139.315 172.915 ;
        RECT 139.605 172.745 139.775 172.915 ;
        RECT 140.065 172.745 140.235 172.915 ;
        RECT 140.525 172.745 140.695 172.915 ;
        RECT 140.985 172.745 141.155 172.915 ;
        RECT 141.445 172.745 141.615 172.915 ;
        RECT 141.905 172.745 142.075 172.915 ;
        RECT 142.365 172.745 142.535 172.915 ;
        RECT 142.825 172.745 142.995 172.915 ;
        RECT 143.285 172.745 143.455 172.915 ;
        RECT 143.745 172.745 143.915 172.915 ;
        RECT 144.205 172.745 144.375 172.915 ;
        RECT 144.665 172.745 144.835 172.915 ;
        RECT 145.125 172.745 145.295 172.915 ;
        RECT 145.585 172.745 145.755 172.915 ;
        RECT 146.045 172.745 146.215 172.915 ;
        RECT 146.505 172.745 146.675 172.915 ;
        RECT 146.965 172.745 147.135 172.915 ;
        RECT 147.425 172.745 147.595 172.915 ;
        RECT 147.885 172.745 148.055 172.915 ;
        RECT 148.345 172.745 148.515 172.915 ;
        RECT 148.805 172.745 148.975 172.915 ;
        RECT 149.265 172.745 149.435 172.915 ;
        RECT 149.725 172.745 149.895 172.915 ;
        RECT 150.185 172.745 150.355 172.915 ;
        RECT 14.945 171.555 15.115 171.725 ;
        RECT 15.430 170.875 15.600 171.045 ;
        RECT 15.825 171.215 15.995 171.385 ;
        RECT 16.280 171.895 16.450 172.065 ;
        RECT 17.015 171.215 17.185 171.385 ;
        RECT 17.530 170.875 17.700 171.045 ;
        RECT 19.100 170.875 19.270 171.045 ;
        RECT 19.535 171.215 19.705 171.385 ;
        RECT 21.845 170.535 22.015 170.705 ;
        RECT 24.065 171.895 24.235 172.065 ;
        RECT 25.065 171.895 25.235 172.065 ;
        RECT 23.225 170.875 23.395 171.045 ;
        RECT 24.145 170.535 24.315 170.705 ;
        RECT 28.285 170.875 28.455 171.045 ;
        RECT 30.125 172.235 30.295 172.405 ;
        RECT 30.125 170.535 30.295 170.705 ;
        RECT 31.045 170.535 31.215 170.705 ;
        RECT 32.425 172.235 32.595 172.405 ;
        RECT 33.345 171.215 33.515 171.385 ;
        RECT 33.805 171.215 33.975 171.385 ;
        RECT 34.265 171.555 34.435 171.725 ;
        RECT 34.725 171.215 34.895 171.385 ;
        RECT 38.865 171.555 39.035 171.725 ;
        RECT 41.625 172.235 41.795 172.405 ;
        RECT 40.705 171.895 40.875 172.065 ;
        RECT 43.925 172.235 44.095 172.405 ;
        RECT 42.085 171.555 42.255 171.725 ;
        RECT 40.705 170.535 40.875 170.705 ;
        RECT 42.545 171.215 42.715 171.385 ;
        RECT 44.845 172.235 45.015 172.405 ;
        RECT 45.400 171.895 45.570 172.065 ;
        RECT 46.225 172.235 46.395 172.405 ;
        RECT 44.385 171.555 44.555 171.725 ;
        RECT 50.365 172.235 50.535 172.405 ;
        RECT 42.545 170.535 42.715 170.705 ;
        RECT 46.225 171.215 46.395 171.385 ;
        RECT 48.525 171.555 48.695 171.725 ;
        RECT 49.445 171.555 49.615 171.725 ;
        RECT 58.185 171.555 58.355 171.725 ;
        RECT 58.645 171.555 58.815 171.725 ;
        RECT 59.105 170.535 59.275 170.705 ;
        RECT 60.025 170.535 60.195 170.705 ;
        RECT 63.245 171.215 63.415 171.385 ;
        RECT 63.730 170.875 63.900 171.045 ;
        RECT 64.125 171.215 64.295 171.385 ;
        RECT 64.580 171.895 64.750 172.065 ;
        RECT 65.315 171.215 65.485 171.385 ;
        RECT 65.830 170.875 66.000 171.045 ;
        RECT 67.400 170.875 67.570 171.045 ;
        RECT 67.835 171.215 68.005 171.385 ;
        RECT 70.145 172.235 70.315 172.405 ;
        RECT 76.125 172.235 76.295 172.405 ;
        RECT 73.825 171.555 73.995 171.725 ;
        RECT 74.285 171.555 74.455 171.725 ;
        RECT 73.365 170.535 73.535 170.705 ;
        RECT 74.745 171.215 74.915 171.385 ;
        RECT 74.745 170.535 74.915 170.705 ;
        RECT 76.585 172.235 76.755 172.405 ;
        RECT 77.425 172.235 77.595 172.405 ;
        RECT 78.425 171.895 78.595 172.065 ;
        RECT 78.885 171.555 79.055 171.725 ;
        RECT 79.370 170.875 79.540 171.045 ;
        RECT 79.765 171.215 79.935 171.385 ;
        RECT 77.505 170.535 77.675 170.705 ;
        RECT 80.165 171.555 80.335 171.725 ;
        RECT 80.955 171.215 81.125 171.385 ;
        RECT 81.470 170.875 81.640 171.045 ;
        RECT 83.040 170.875 83.210 171.045 ;
        RECT 83.475 171.215 83.645 171.385 ;
        RECT 85.785 172.235 85.955 172.405 ;
        RECT 91.765 172.235 91.935 172.405 ;
        RECT 89.465 171.555 89.635 171.725 ;
        RECT 94.525 172.235 94.695 172.405 ;
        RECT 92.225 171.555 92.395 171.725 ;
        RECT 89.925 170.535 90.095 170.705 ;
        RECT 92.685 170.535 92.855 170.705 ;
        RECT 102.805 171.555 102.975 171.725 ;
        RECT 102.345 170.535 102.515 170.705 ;
        RECT 106.025 171.555 106.195 171.725 ;
        RECT 112.005 172.235 112.175 172.405 ;
        RECT 112.925 171.555 113.095 171.725 ;
        RECT 113.845 171.555 114.015 171.725 ;
        RECT 114.765 171.555 114.935 171.725 ;
        RECT 115.685 172.235 115.855 172.405 ;
        RECT 118.905 172.235 119.075 172.405 ;
        RECT 116.145 171.555 116.315 171.725 ;
        RECT 117.065 171.555 117.235 171.725 ;
        RECT 117.985 171.895 118.155 172.065 ;
        RECT 114.765 170.535 114.935 170.705 ;
        RECT 123.045 171.215 123.215 171.385 ;
        RECT 123.530 170.875 123.700 171.045 ;
        RECT 123.925 171.215 124.095 171.385 ;
        RECT 124.380 171.555 124.550 171.725 ;
        RECT 125.115 171.215 125.285 171.385 ;
        RECT 125.630 170.875 125.800 171.045 ;
        RECT 127.200 170.875 127.370 171.045 ;
        RECT 127.635 171.215 127.805 171.385 ;
        RECT 129.945 172.235 130.115 172.405 ;
        RECT 11.265 170.025 11.435 170.195 ;
        RECT 11.725 170.025 11.895 170.195 ;
        RECT 12.185 170.025 12.355 170.195 ;
        RECT 12.645 170.025 12.815 170.195 ;
        RECT 13.105 170.025 13.275 170.195 ;
        RECT 13.565 170.025 13.735 170.195 ;
        RECT 14.025 170.025 14.195 170.195 ;
        RECT 14.485 170.025 14.655 170.195 ;
        RECT 14.945 170.025 15.115 170.195 ;
        RECT 15.405 170.025 15.575 170.195 ;
        RECT 15.865 170.025 16.035 170.195 ;
        RECT 16.325 170.025 16.495 170.195 ;
        RECT 16.785 170.025 16.955 170.195 ;
        RECT 17.245 170.025 17.415 170.195 ;
        RECT 17.705 170.025 17.875 170.195 ;
        RECT 18.165 170.025 18.335 170.195 ;
        RECT 18.625 170.025 18.795 170.195 ;
        RECT 19.085 170.025 19.255 170.195 ;
        RECT 19.545 170.025 19.715 170.195 ;
        RECT 20.005 170.025 20.175 170.195 ;
        RECT 20.465 170.025 20.635 170.195 ;
        RECT 20.925 170.025 21.095 170.195 ;
        RECT 21.385 170.025 21.555 170.195 ;
        RECT 21.845 170.025 22.015 170.195 ;
        RECT 22.305 170.025 22.475 170.195 ;
        RECT 22.765 170.025 22.935 170.195 ;
        RECT 23.225 170.025 23.395 170.195 ;
        RECT 23.685 170.025 23.855 170.195 ;
        RECT 24.145 170.025 24.315 170.195 ;
        RECT 24.605 170.025 24.775 170.195 ;
        RECT 25.065 170.025 25.235 170.195 ;
        RECT 25.525 170.025 25.695 170.195 ;
        RECT 25.985 170.025 26.155 170.195 ;
        RECT 26.445 170.025 26.615 170.195 ;
        RECT 26.905 170.025 27.075 170.195 ;
        RECT 27.365 170.025 27.535 170.195 ;
        RECT 27.825 170.025 27.995 170.195 ;
        RECT 28.285 170.025 28.455 170.195 ;
        RECT 28.745 170.025 28.915 170.195 ;
        RECT 29.205 170.025 29.375 170.195 ;
        RECT 29.665 170.025 29.835 170.195 ;
        RECT 30.125 170.025 30.295 170.195 ;
        RECT 30.585 170.025 30.755 170.195 ;
        RECT 31.045 170.025 31.215 170.195 ;
        RECT 31.505 170.025 31.675 170.195 ;
        RECT 31.965 170.025 32.135 170.195 ;
        RECT 32.425 170.025 32.595 170.195 ;
        RECT 32.885 170.025 33.055 170.195 ;
        RECT 33.345 170.025 33.515 170.195 ;
        RECT 33.805 170.025 33.975 170.195 ;
        RECT 34.265 170.025 34.435 170.195 ;
        RECT 34.725 170.025 34.895 170.195 ;
        RECT 35.185 170.025 35.355 170.195 ;
        RECT 35.645 170.025 35.815 170.195 ;
        RECT 36.105 170.025 36.275 170.195 ;
        RECT 36.565 170.025 36.735 170.195 ;
        RECT 37.025 170.025 37.195 170.195 ;
        RECT 37.485 170.025 37.655 170.195 ;
        RECT 37.945 170.025 38.115 170.195 ;
        RECT 38.405 170.025 38.575 170.195 ;
        RECT 38.865 170.025 39.035 170.195 ;
        RECT 39.325 170.025 39.495 170.195 ;
        RECT 39.785 170.025 39.955 170.195 ;
        RECT 40.245 170.025 40.415 170.195 ;
        RECT 40.705 170.025 40.875 170.195 ;
        RECT 41.165 170.025 41.335 170.195 ;
        RECT 41.625 170.025 41.795 170.195 ;
        RECT 42.085 170.025 42.255 170.195 ;
        RECT 42.545 170.025 42.715 170.195 ;
        RECT 43.005 170.025 43.175 170.195 ;
        RECT 43.465 170.025 43.635 170.195 ;
        RECT 43.925 170.025 44.095 170.195 ;
        RECT 44.385 170.025 44.555 170.195 ;
        RECT 44.845 170.025 45.015 170.195 ;
        RECT 45.305 170.025 45.475 170.195 ;
        RECT 45.765 170.025 45.935 170.195 ;
        RECT 46.225 170.025 46.395 170.195 ;
        RECT 46.685 170.025 46.855 170.195 ;
        RECT 47.145 170.025 47.315 170.195 ;
        RECT 47.605 170.025 47.775 170.195 ;
        RECT 48.065 170.025 48.235 170.195 ;
        RECT 48.525 170.025 48.695 170.195 ;
        RECT 48.985 170.025 49.155 170.195 ;
        RECT 49.445 170.025 49.615 170.195 ;
        RECT 49.905 170.025 50.075 170.195 ;
        RECT 50.365 170.025 50.535 170.195 ;
        RECT 50.825 170.025 50.995 170.195 ;
        RECT 51.285 170.025 51.455 170.195 ;
        RECT 51.745 170.025 51.915 170.195 ;
        RECT 52.205 170.025 52.375 170.195 ;
        RECT 52.665 170.025 52.835 170.195 ;
        RECT 53.125 170.025 53.295 170.195 ;
        RECT 53.585 170.025 53.755 170.195 ;
        RECT 54.045 170.025 54.215 170.195 ;
        RECT 54.505 170.025 54.675 170.195 ;
        RECT 54.965 170.025 55.135 170.195 ;
        RECT 55.425 170.025 55.595 170.195 ;
        RECT 55.885 170.025 56.055 170.195 ;
        RECT 56.345 170.025 56.515 170.195 ;
        RECT 56.805 170.025 56.975 170.195 ;
        RECT 57.265 170.025 57.435 170.195 ;
        RECT 57.725 170.025 57.895 170.195 ;
        RECT 58.185 170.025 58.355 170.195 ;
        RECT 58.645 170.025 58.815 170.195 ;
        RECT 59.105 170.025 59.275 170.195 ;
        RECT 59.565 170.025 59.735 170.195 ;
        RECT 60.025 170.025 60.195 170.195 ;
        RECT 60.485 170.025 60.655 170.195 ;
        RECT 60.945 170.025 61.115 170.195 ;
        RECT 61.405 170.025 61.575 170.195 ;
        RECT 61.865 170.025 62.035 170.195 ;
        RECT 62.325 170.025 62.495 170.195 ;
        RECT 62.785 170.025 62.955 170.195 ;
        RECT 63.245 170.025 63.415 170.195 ;
        RECT 63.705 170.025 63.875 170.195 ;
        RECT 64.165 170.025 64.335 170.195 ;
        RECT 64.625 170.025 64.795 170.195 ;
        RECT 65.085 170.025 65.255 170.195 ;
        RECT 65.545 170.025 65.715 170.195 ;
        RECT 66.005 170.025 66.175 170.195 ;
        RECT 66.465 170.025 66.635 170.195 ;
        RECT 66.925 170.025 67.095 170.195 ;
        RECT 67.385 170.025 67.555 170.195 ;
        RECT 67.845 170.025 68.015 170.195 ;
        RECT 68.305 170.025 68.475 170.195 ;
        RECT 68.765 170.025 68.935 170.195 ;
        RECT 69.225 170.025 69.395 170.195 ;
        RECT 69.685 170.025 69.855 170.195 ;
        RECT 70.145 170.025 70.315 170.195 ;
        RECT 70.605 170.025 70.775 170.195 ;
        RECT 71.065 170.025 71.235 170.195 ;
        RECT 71.525 170.025 71.695 170.195 ;
        RECT 71.985 170.025 72.155 170.195 ;
        RECT 72.445 170.025 72.615 170.195 ;
        RECT 72.905 170.025 73.075 170.195 ;
        RECT 73.365 170.025 73.535 170.195 ;
        RECT 73.825 170.025 73.995 170.195 ;
        RECT 74.285 170.025 74.455 170.195 ;
        RECT 74.745 170.025 74.915 170.195 ;
        RECT 75.205 170.025 75.375 170.195 ;
        RECT 75.665 170.025 75.835 170.195 ;
        RECT 76.125 170.025 76.295 170.195 ;
        RECT 76.585 170.025 76.755 170.195 ;
        RECT 77.045 170.025 77.215 170.195 ;
        RECT 77.505 170.025 77.675 170.195 ;
        RECT 77.965 170.025 78.135 170.195 ;
        RECT 78.425 170.025 78.595 170.195 ;
        RECT 78.885 170.025 79.055 170.195 ;
        RECT 79.345 170.025 79.515 170.195 ;
        RECT 79.805 170.025 79.975 170.195 ;
        RECT 80.265 170.025 80.435 170.195 ;
        RECT 80.725 170.025 80.895 170.195 ;
        RECT 81.185 170.025 81.355 170.195 ;
        RECT 81.645 170.025 81.815 170.195 ;
        RECT 82.105 170.025 82.275 170.195 ;
        RECT 82.565 170.025 82.735 170.195 ;
        RECT 83.025 170.025 83.195 170.195 ;
        RECT 83.485 170.025 83.655 170.195 ;
        RECT 83.945 170.025 84.115 170.195 ;
        RECT 84.405 170.025 84.575 170.195 ;
        RECT 84.865 170.025 85.035 170.195 ;
        RECT 85.325 170.025 85.495 170.195 ;
        RECT 85.785 170.025 85.955 170.195 ;
        RECT 86.245 170.025 86.415 170.195 ;
        RECT 86.705 170.025 86.875 170.195 ;
        RECT 87.165 170.025 87.335 170.195 ;
        RECT 87.625 170.025 87.795 170.195 ;
        RECT 88.085 170.025 88.255 170.195 ;
        RECT 88.545 170.025 88.715 170.195 ;
        RECT 89.005 170.025 89.175 170.195 ;
        RECT 89.465 170.025 89.635 170.195 ;
        RECT 89.925 170.025 90.095 170.195 ;
        RECT 90.385 170.025 90.555 170.195 ;
        RECT 90.845 170.025 91.015 170.195 ;
        RECT 91.305 170.025 91.475 170.195 ;
        RECT 91.765 170.025 91.935 170.195 ;
        RECT 92.225 170.025 92.395 170.195 ;
        RECT 92.685 170.025 92.855 170.195 ;
        RECT 93.145 170.025 93.315 170.195 ;
        RECT 93.605 170.025 93.775 170.195 ;
        RECT 94.065 170.025 94.235 170.195 ;
        RECT 94.525 170.025 94.695 170.195 ;
        RECT 94.985 170.025 95.155 170.195 ;
        RECT 95.445 170.025 95.615 170.195 ;
        RECT 95.905 170.025 96.075 170.195 ;
        RECT 96.365 170.025 96.535 170.195 ;
        RECT 96.825 170.025 96.995 170.195 ;
        RECT 97.285 170.025 97.455 170.195 ;
        RECT 97.745 170.025 97.915 170.195 ;
        RECT 98.205 170.025 98.375 170.195 ;
        RECT 98.665 170.025 98.835 170.195 ;
        RECT 99.125 170.025 99.295 170.195 ;
        RECT 99.585 170.025 99.755 170.195 ;
        RECT 100.045 170.025 100.215 170.195 ;
        RECT 100.505 170.025 100.675 170.195 ;
        RECT 100.965 170.025 101.135 170.195 ;
        RECT 101.425 170.025 101.595 170.195 ;
        RECT 101.885 170.025 102.055 170.195 ;
        RECT 102.345 170.025 102.515 170.195 ;
        RECT 102.805 170.025 102.975 170.195 ;
        RECT 103.265 170.025 103.435 170.195 ;
        RECT 103.725 170.025 103.895 170.195 ;
        RECT 104.185 170.025 104.355 170.195 ;
        RECT 104.645 170.025 104.815 170.195 ;
        RECT 105.105 170.025 105.275 170.195 ;
        RECT 105.565 170.025 105.735 170.195 ;
        RECT 106.025 170.025 106.195 170.195 ;
        RECT 106.485 170.025 106.655 170.195 ;
        RECT 106.945 170.025 107.115 170.195 ;
        RECT 107.405 170.025 107.575 170.195 ;
        RECT 107.865 170.025 108.035 170.195 ;
        RECT 108.325 170.025 108.495 170.195 ;
        RECT 108.785 170.025 108.955 170.195 ;
        RECT 109.245 170.025 109.415 170.195 ;
        RECT 109.705 170.025 109.875 170.195 ;
        RECT 110.165 170.025 110.335 170.195 ;
        RECT 110.625 170.025 110.795 170.195 ;
        RECT 111.085 170.025 111.255 170.195 ;
        RECT 111.545 170.025 111.715 170.195 ;
        RECT 112.005 170.025 112.175 170.195 ;
        RECT 112.465 170.025 112.635 170.195 ;
        RECT 112.925 170.025 113.095 170.195 ;
        RECT 113.385 170.025 113.555 170.195 ;
        RECT 113.845 170.025 114.015 170.195 ;
        RECT 114.305 170.025 114.475 170.195 ;
        RECT 114.765 170.025 114.935 170.195 ;
        RECT 115.225 170.025 115.395 170.195 ;
        RECT 115.685 170.025 115.855 170.195 ;
        RECT 116.145 170.025 116.315 170.195 ;
        RECT 116.605 170.025 116.775 170.195 ;
        RECT 117.065 170.025 117.235 170.195 ;
        RECT 117.525 170.025 117.695 170.195 ;
        RECT 117.985 170.025 118.155 170.195 ;
        RECT 118.445 170.025 118.615 170.195 ;
        RECT 118.905 170.025 119.075 170.195 ;
        RECT 119.365 170.025 119.535 170.195 ;
        RECT 119.825 170.025 119.995 170.195 ;
        RECT 120.285 170.025 120.455 170.195 ;
        RECT 120.745 170.025 120.915 170.195 ;
        RECT 121.205 170.025 121.375 170.195 ;
        RECT 121.665 170.025 121.835 170.195 ;
        RECT 122.125 170.025 122.295 170.195 ;
        RECT 122.585 170.025 122.755 170.195 ;
        RECT 123.045 170.025 123.215 170.195 ;
        RECT 123.505 170.025 123.675 170.195 ;
        RECT 123.965 170.025 124.135 170.195 ;
        RECT 124.425 170.025 124.595 170.195 ;
        RECT 124.885 170.025 125.055 170.195 ;
        RECT 125.345 170.025 125.515 170.195 ;
        RECT 125.805 170.025 125.975 170.195 ;
        RECT 126.265 170.025 126.435 170.195 ;
        RECT 126.725 170.025 126.895 170.195 ;
        RECT 127.185 170.025 127.355 170.195 ;
        RECT 127.645 170.025 127.815 170.195 ;
        RECT 128.105 170.025 128.275 170.195 ;
        RECT 128.565 170.025 128.735 170.195 ;
        RECT 129.025 170.025 129.195 170.195 ;
        RECT 129.485 170.025 129.655 170.195 ;
        RECT 129.945 170.025 130.115 170.195 ;
        RECT 130.405 170.025 130.575 170.195 ;
        RECT 130.865 170.025 131.035 170.195 ;
        RECT 131.325 170.025 131.495 170.195 ;
        RECT 131.785 170.025 131.955 170.195 ;
        RECT 132.245 170.025 132.415 170.195 ;
        RECT 132.705 170.025 132.875 170.195 ;
        RECT 133.165 170.025 133.335 170.195 ;
        RECT 133.625 170.025 133.795 170.195 ;
        RECT 134.085 170.025 134.255 170.195 ;
        RECT 134.545 170.025 134.715 170.195 ;
        RECT 135.005 170.025 135.175 170.195 ;
        RECT 135.465 170.025 135.635 170.195 ;
        RECT 135.925 170.025 136.095 170.195 ;
        RECT 136.385 170.025 136.555 170.195 ;
        RECT 136.845 170.025 137.015 170.195 ;
        RECT 137.305 170.025 137.475 170.195 ;
        RECT 137.765 170.025 137.935 170.195 ;
        RECT 138.225 170.025 138.395 170.195 ;
        RECT 138.685 170.025 138.855 170.195 ;
        RECT 139.145 170.025 139.315 170.195 ;
        RECT 139.605 170.025 139.775 170.195 ;
        RECT 140.065 170.025 140.235 170.195 ;
        RECT 140.525 170.025 140.695 170.195 ;
        RECT 140.985 170.025 141.155 170.195 ;
        RECT 141.445 170.025 141.615 170.195 ;
        RECT 141.905 170.025 142.075 170.195 ;
        RECT 142.365 170.025 142.535 170.195 ;
        RECT 142.825 170.025 142.995 170.195 ;
        RECT 143.285 170.025 143.455 170.195 ;
        RECT 143.745 170.025 143.915 170.195 ;
        RECT 144.205 170.025 144.375 170.195 ;
        RECT 144.665 170.025 144.835 170.195 ;
        RECT 145.125 170.025 145.295 170.195 ;
        RECT 145.585 170.025 145.755 170.195 ;
        RECT 146.045 170.025 146.215 170.195 ;
        RECT 146.505 170.025 146.675 170.195 ;
        RECT 146.965 170.025 147.135 170.195 ;
        RECT 147.425 170.025 147.595 170.195 ;
        RECT 147.885 170.025 148.055 170.195 ;
        RECT 148.345 170.025 148.515 170.195 ;
        RECT 148.805 170.025 148.975 170.195 ;
        RECT 149.265 170.025 149.435 170.195 ;
        RECT 149.725 170.025 149.895 170.195 ;
        RECT 150.185 170.025 150.355 170.195 ;
        RECT 15.405 169.175 15.575 169.345 ;
        RECT 17.245 169.515 17.415 169.685 ;
        RECT 18.165 169.515 18.335 169.685 ;
        RECT 17.245 168.155 17.415 168.325 ;
        RECT 20.465 168.495 20.635 168.665 ;
        RECT 21.385 168.495 21.555 168.665 ;
        RECT 20.925 167.815 21.095 167.985 ;
        RECT 21.845 168.155 22.015 168.325 ;
        RECT 22.765 168.155 22.935 168.325 ;
        RECT 23.685 168.155 23.855 168.325 ;
        RECT 26.445 168.835 26.615 169.005 ;
        RECT 25.525 168.495 25.695 168.665 ;
        RECT 26.905 168.835 27.075 169.005 ;
        RECT 29.690 169.175 29.860 169.345 ;
        RECT 24.605 168.155 24.775 168.325 ;
        RECT 27.825 168.495 27.995 168.665 ;
        RECT 28.285 168.495 28.455 168.665 ;
        RECT 29.205 168.495 29.375 168.665 ;
        RECT 30.085 168.835 30.255 169.005 ;
        RECT 30.540 168.155 30.710 168.325 ;
        RECT 31.790 169.175 31.960 169.345 ;
        RECT 31.275 168.835 31.445 169.005 ;
        RECT 33.360 169.175 33.530 169.345 ;
        RECT 33.795 168.835 33.965 169.005 ;
        RECT 36.105 169.515 36.275 169.685 ;
        RECT 38.865 169.515 39.035 169.685 ;
        RECT 37.945 167.815 38.115 167.985 ;
        RECT 38.785 167.815 38.955 167.985 ;
        RECT 39.785 168.155 39.955 168.325 ;
        RECT 43.005 169.515 43.175 169.685 ;
        RECT 41.625 168.495 41.795 168.665 ;
        RECT 42.085 168.155 42.255 168.325 ;
        RECT 43.005 168.495 43.175 168.665 ;
        RECT 51.745 168.835 51.915 169.005 ;
        RECT 52.205 168.495 52.375 168.665 ;
        RECT 50.365 167.815 50.535 167.985 ;
        RECT 55.885 168.835 56.055 169.005 ;
        RECT 55.425 168.495 55.595 168.665 ;
        RECT 53.585 167.815 53.755 167.985 ;
        RECT 56.805 169.175 56.975 169.345 ;
        RECT 58.645 169.175 58.815 169.345 ;
        RECT 57.725 168.495 57.895 168.665 ;
        RECT 59.105 168.495 59.275 168.665 ;
        RECT 60.025 168.495 60.195 168.665 ;
        RECT 60.485 168.495 60.655 168.665 ;
        RECT 67.410 169.175 67.580 169.345 ;
        RECT 66.925 168.495 67.095 168.665 ;
        RECT 67.805 168.835 67.975 169.005 ;
        RECT 68.260 168.155 68.430 168.325 ;
        RECT 69.510 169.175 69.680 169.345 ;
        RECT 68.995 168.835 69.165 169.005 ;
        RECT 71.080 169.175 71.250 169.345 ;
        RECT 71.515 168.835 71.685 169.005 ;
        RECT 73.825 169.175 73.995 169.345 ;
        RECT 78.425 169.175 78.595 169.345 ;
        RECT 88.545 169.515 88.715 169.685 ;
        RECT 84.865 168.155 85.035 168.325 ;
        RECT 87.165 168.835 87.335 169.005 ;
        RECT 86.705 168.495 86.875 168.665 ;
        RECT 98.205 168.495 98.375 168.665 ;
        RECT 98.665 168.495 98.835 168.665 ;
        RECT 99.585 168.495 99.755 168.665 ;
        RECT 100.045 168.495 100.215 168.665 ;
        RECT 102.370 169.175 102.540 169.345 ;
        RECT 101.885 168.495 102.055 168.665 ;
        RECT 100.965 167.815 101.135 167.985 ;
        RECT 102.765 168.835 102.935 169.005 ;
        RECT 103.220 168.155 103.390 168.325 ;
        RECT 104.470 169.175 104.640 169.345 ;
        RECT 103.955 168.835 104.125 169.005 ;
        RECT 106.040 169.175 106.210 169.345 ;
        RECT 106.475 168.835 106.645 169.005 ;
        RECT 108.785 169.515 108.955 169.685 ;
        RECT 111.085 169.515 111.255 169.685 ;
        RECT 111.545 168.835 111.715 169.005 ;
        RECT 112.005 169.175 112.175 169.345 ;
        RECT 113.385 168.495 113.555 168.665 ;
        RECT 117.525 169.515 117.695 169.685 ;
        RECT 109.705 167.815 109.875 167.985 ;
        RECT 112.925 167.815 113.095 167.985 ;
        RECT 117.445 168.155 117.615 168.325 ;
        RECT 116.605 167.815 116.775 167.985 ;
        RECT 118.905 168.495 119.075 168.665 ;
        RECT 118.445 168.155 118.615 168.325 ;
        RECT 119.825 168.495 119.995 168.665 ;
        RECT 121.205 168.495 121.375 168.665 ;
        RECT 122.125 168.495 122.295 168.665 ;
        RECT 123.045 168.495 123.215 168.665 ;
        RECT 124.425 169.515 124.595 169.685 ;
        RECT 125.345 168.495 125.515 168.665 ;
        RECT 11.265 167.305 11.435 167.475 ;
        RECT 11.725 167.305 11.895 167.475 ;
        RECT 12.185 167.305 12.355 167.475 ;
        RECT 12.645 167.305 12.815 167.475 ;
        RECT 13.105 167.305 13.275 167.475 ;
        RECT 13.565 167.305 13.735 167.475 ;
        RECT 14.025 167.305 14.195 167.475 ;
        RECT 14.485 167.305 14.655 167.475 ;
        RECT 14.945 167.305 15.115 167.475 ;
        RECT 15.405 167.305 15.575 167.475 ;
        RECT 15.865 167.305 16.035 167.475 ;
        RECT 16.325 167.305 16.495 167.475 ;
        RECT 16.785 167.305 16.955 167.475 ;
        RECT 17.245 167.305 17.415 167.475 ;
        RECT 17.705 167.305 17.875 167.475 ;
        RECT 18.165 167.305 18.335 167.475 ;
        RECT 18.625 167.305 18.795 167.475 ;
        RECT 19.085 167.305 19.255 167.475 ;
        RECT 19.545 167.305 19.715 167.475 ;
        RECT 20.005 167.305 20.175 167.475 ;
        RECT 20.465 167.305 20.635 167.475 ;
        RECT 20.925 167.305 21.095 167.475 ;
        RECT 21.385 167.305 21.555 167.475 ;
        RECT 21.845 167.305 22.015 167.475 ;
        RECT 22.305 167.305 22.475 167.475 ;
        RECT 22.765 167.305 22.935 167.475 ;
        RECT 23.225 167.305 23.395 167.475 ;
        RECT 23.685 167.305 23.855 167.475 ;
        RECT 24.145 167.305 24.315 167.475 ;
        RECT 24.605 167.305 24.775 167.475 ;
        RECT 25.065 167.305 25.235 167.475 ;
        RECT 25.525 167.305 25.695 167.475 ;
        RECT 25.985 167.305 26.155 167.475 ;
        RECT 26.445 167.305 26.615 167.475 ;
        RECT 26.905 167.305 27.075 167.475 ;
        RECT 27.365 167.305 27.535 167.475 ;
        RECT 27.825 167.305 27.995 167.475 ;
        RECT 28.285 167.305 28.455 167.475 ;
        RECT 28.745 167.305 28.915 167.475 ;
        RECT 29.205 167.305 29.375 167.475 ;
        RECT 29.665 167.305 29.835 167.475 ;
        RECT 30.125 167.305 30.295 167.475 ;
        RECT 30.585 167.305 30.755 167.475 ;
        RECT 31.045 167.305 31.215 167.475 ;
        RECT 31.505 167.305 31.675 167.475 ;
        RECT 31.965 167.305 32.135 167.475 ;
        RECT 32.425 167.305 32.595 167.475 ;
        RECT 32.885 167.305 33.055 167.475 ;
        RECT 33.345 167.305 33.515 167.475 ;
        RECT 33.805 167.305 33.975 167.475 ;
        RECT 34.265 167.305 34.435 167.475 ;
        RECT 34.725 167.305 34.895 167.475 ;
        RECT 35.185 167.305 35.355 167.475 ;
        RECT 35.645 167.305 35.815 167.475 ;
        RECT 36.105 167.305 36.275 167.475 ;
        RECT 36.565 167.305 36.735 167.475 ;
        RECT 37.025 167.305 37.195 167.475 ;
        RECT 37.485 167.305 37.655 167.475 ;
        RECT 37.945 167.305 38.115 167.475 ;
        RECT 38.405 167.305 38.575 167.475 ;
        RECT 38.865 167.305 39.035 167.475 ;
        RECT 39.325 167.305 39.495 167.475 ;
        RECT 39.785 167.305 39.955 167.475 ;
        RECT 40.245 167.305 40.415 167.475 ;
        RECT 40.705 167.305 40.875 167.475 ;
        RECT 41.165 167.305 41.335 167.475 ;
        RECT 41.625 167.305 41.795 167.475 ;
        RECT 42.085 167.305 42.255 167.475 ;
        RECT 42.545 167.305 42.715 167.475 ;
        RECT 43.005 167.305 43.175 167.475 ;
        RECT 43.465 167.305 43.635 167.475 ;
        RECT 43.925 167.305 44.095 167.475 ;
        RECT 44.385 167.305 44.555 167.475 ;
        RECT 44.845 167.305 45.015 167.475 ;
        RECT 45.305 167.305 45.475 167.475 ;
        RECT 45.765 167.305 45.935 167.475 ;
        RECT 46.225 167.305 46.395 167.475 ;
        RECT 46.685 167.305 46.855 167.475 ;
        RECT 47.145 167.305 47.315 167.475 ;
        RECT 47.605 167.305 47.775 167.475 ;
        RECT 48.065 167.305 48.235 167.475 ;
        RECT 48.525 167.305 48.695 167.475 ;
        RECT 48.985 167.305 49.155 167.475 ;
        RECT 49.445 167.305 49.615 167.475 ;
        RECT 49.905 167.305 50.075 167.475 ;
        RECT 50.365 167.305 50.535 167.475 ;
        RECT 50.825 167.305 50.995 167.475 ;
        RECT 51.285 167.305 51.455 167.475 ;
        RECT 51.745 167.305 51.915 167.475 ;
        RECT 52.205 167.305 52.375 167.475 ;
        RECT 52.665 167.305 52.835 167.475 ;
        RECT 53.125 167.305 53.295 167.475 ;
        RECT 53.585 167.305 53.755 167.475 ;
        RECT 54.045 167.305 54.215 167.475 ;
        RECT 54.505 167.305 54.675 167.475 ;
        RECT 54.965 167.305 55.135 167.475 ;
        RECT 55.425 167.305 55.595 167.475 ;
        RECT 55.885 167.305 56.055 167.475 ;
        RECT 56.345 167.305 56.515 167.475 ;
        RECT 56.805 167.305 56.975 167.475 ;
        RECT 57.265 167.305 57.435 167.475 ;
        RECT 57.725 167.305 57.895 167.475 ;
        RECT 58.185 167.305 58.355 167.475 ;
        RECT 58.645 167.305 58.815 167.475 ;
        RECT 59.105 167.305 59.275 167.475 ;
        RECT 59.565 167.305 59.735 167.475 ;
        RECT 60.025 167.305 60.195 167.475 ;
        RECT 60.485 167.305 60.655 167.475 ;
        RECT 60.945 167.305 61.115 167.475 ;
        RECT 61.405 167.305 61.575 167.475 ;
        RECT 61.865 167.305 62.035 167.475 ;
        RECT 62.325 167.305 62.495 167.475 ;
        RECT 62.785 167.305 62.955 167.475 ;
        RECT 63.245 167.305 63.415 167.475 ;
        RECT 63.705 167.305 63.875 167.475 ;
        RECT 64.165 167.305 64.335 167.475 ;
        RECT 64.625 167.305 64.795 167.475 ;
        RECT 65.085 167.305 65.255 167.475 ;
        RECT 65.545 167.305 65.715 167.475 ;
        RECT 66.005 167.305 66.175 167.475 ;
        RECT 66.465 167.305 66.635 167.475 ;
        RECT 66.925 167.305 67.095 167.475 ;
        RECT 67.385 167.305 67.555 167.475 ;
        RECT 67.845 167.305 68.015 167.475 ;
        RECT 68.305 167.305 68.475 167.475 ;
        RECT 68.765 167.305 68.935 167.475 ;
        RECT 69.225 167.305 69.395 167.475 ;
        RECT 69.685 167.305 69.855 167.475 ;
        RECT 70.145 167.305 70.315 167.475 ;
        RECT 70.605 167.305 70.775 167.475 ;
        RECT 71.065 167.305 71.235 167.475 ;
        RECT 71.525 167.305 71.695 167.475 ;
        RECT 71.985 167.305 72.155 167.475 ;
        RECT 72.445 167.305 72.615 167.475 ;
        RECT 72.905 167.305 73.075 167.475 ;
        RECT 73.365 167.305 73.535 167.475 ;
        RECT 73.825 167.305 73.995 167.475 ;
        RECT 74.285 167.305 74.455 167.475 ;
        RECT 74.745 167.305 74.915 167.475 ;
        RECT 75.205 167.305 75.375 167.475 ;
        RECT 75.665 167.305 75.835 167.475 ;
        RECT 76.125 167.305 76.295 167.475 ;
        RECT 76.585 167.305 76.755 167.475 ;
        RECT 77.045 167.305 77.215 167.475 ;
        RECT 77.505 167.305 77.675 167.475 ;
        RECT 77.965 167.305 78.135 167.475 ;
        RECT 78.425 167.305 78.595 167.475 ;
        RECT 78.885 167.305 79.055 167.475 ;
        RECT 79.345 167.305 79.515 167.475 ;
        RECT 79.805 167.305 79.975 167.475 ;
        RECT 80.265 167.305 80.435 167.475 ;
        RECT 80.725 167.305 80.895 167.475 ;
        RECT 81.185 167.305 81.355 167.475 ;
        RECT 81.645 167.305 81.815 167.475 ;
        RECT 82.105 167.305 82.275 167.475 ;
        RECT 82.565 167.305 82.735 167.475 ;
        RECT 83.025 167.305 83.195 167.475 ;
        RECT 83.485 167.305 83.655 167.475 ;
        RECT 83.945 167.305 84.115 167.475 ;
        RECT 84.405 167.305 84.575 167.475 ;
        RECT 84.865 167.305 85.035 167.475 ;
        RECT 85.325 167.305 85.495 167.475 ;
        RECT 85.785 167.305 85.955 167.475 ;
        RECT 86.245 167.305 86.415 167.475 ;
        RECT 86.705 167.305 86.875 167.475 ;
        RECT 87.165 167.305 87.335 167.475 ;
        RECT 87.625 167.305 87.795 167.475 ;
        RECT 88.085 167.305 88.255 167.475 ;
        RECT 88.545 167.305 88.715 167.475 ;
        RECT 89.005 167.305 89.175 167.475 ;
        RECT 89.465 167.305 89.635 167.475 ;
        RECT 89.925 167.305 90.095 167.475 ;
        RECT 90.385 167.305 90.555 167.475 ;
        RECT 90.845 167.305 91.015 167.475 ;
        RECT 91.305 167.305 91.475 167.475 ;
        RECT 91.765 167.305 91.935 167.475 ;
        RECT 92.225 167.305 92.395 167.475 ;
        RECT 92.685 167.305 92.855 167.475 ;
        RECT 93.145 167.305 93.315 167.475 ;
        RECT 93.605 167.305 93.775 167.475 ;
        RECT 94.065 167.305 94.235 167.475 ;
        RECT 94.525 167.305 94.695 167.475 ;
        RECT 94.985 167.305 95.155 167.475 ;
        RECT 95.445 167.305 95.615 167.475 ;
        RECT 95.905 167.305 96.075 167.475 ;
        RECT 96.365 167.305 96.535 167.475 ;
        RECT 96.825 167.305 96.995 167.475 ;
        RECT 97.285 167.305 97.455 167.475 ;
        RECT 97.745 167.305 97.915 167.475 ;
        RECT 98.205 167.305 98.375 167.475 ;
        RECT 98.665 167.305 98.835 167.475 ;
        RECT 99.125 167.305 99.295 167.475 ;
        RECT 99.585 167.305 99.755 167.475 ;
        RECT 100.045 167.305 100.215 167.475 ;
        RECT 100.505 167.305 100.675 167.475 ;
        RECT 100.965 167.305 101.135 167.475 ;
        RECT 101.425 167.305 101.595 167.475 ;
        RECT 101.885 167.305 102.055 167.475 ;
        RECT 102.345 167.305 102.515 167.475 ;
        RECT 102.805 167.305 102.975 167.475 ;
        RECT 103.265 167.305 103.435 167.475 ;
        RECT 103.725 167.305 103.895 167.475 ;
        RECT 104.185 167.305 104.355 167.475 ;
        RECT 104.645 167.305 104.815 167.475 ;
        RECT 105.105 167.305 105.275 167.475 ;
        RECT 105.565 167.305 105.735 167.475 ;
        RECT 106.025 167.305 106.195 167.475 ;
        RECT 106.485 167.305 106.655 167.475 ;
        RECT 106.945 167.305 107.115 167.475 ;
        RECT 107.405 167.305 107.575 167.475 ;
        RECT 107.865 167.305 108.035 167.475 ;
        RECT 108.325 167.305 108.495 167.475 ;
        RECT 108.785 167.305 108.955 167.475 ;
        RECT 109.245 167.305 109.415 167.475 ;
        RECT 109.705 167.305 109.875 167.475 ;
        RECT 110.165 167.305 110.335 167.475 ;
        RECT 110.625 167.305 110.795 167.475 ;
        RECT 111.085 167.305 111.255 167.475 ;
        RECT 111.545 167.305 111.715 167.475 ;
        RECT 112.005 167.305 112.175 167.475 ;
        RECT 112.465 167.305 112.635 167.475 ;
        RECT 112.925 167.305 113.095 167.475 ;
        RECT 113.385 167.305 113.555 167.475 ;
        RECT 113.845 167.305 114.015 167.475 ;
        RECT 114.305 167.305 114.475 167.475 ;
        RECT 114.765 167.305 114.935 167.475 ;
        RECT 115.225 167.305 115.395 167.475 ;
        RECT 115.685 167.305 115.855 167.475 ;
        RECT 116.145 167.305 116.315 167.475 ;
        RECT 116.605 167.305 116.775 167.475 ;
        RECT 117.065 167.305 117.235 167.475 ;
        RECT 117.525 167.305 117.695 167.475 ;
        RECT 117.985 167.305 118.155 167.475 ;
        RECT 118.445 167.305 118.615 167.475 ;
        RECT 118.905 167.305 119.075 167.475 ;
        RECT 119.365 167.305 119.535 167.475 ;
        RECT 119.825 167.305 119.995 167.475 ;
        RECT 120.285 167.305 120.455 167.475 ;
        RECT 120.745 167.305 120.915 167.475 ;
        RECT 121.205 167.305 121.375 167.475 ;
        RECT 121.665 167.305 121.835 167.475 ;
        RECT 122.125 167.305 122.295 167.475 ;
        RECT 122.585 167.305 122.755 167.475 ;
        RECT 123.045 167.305 123.215 167.475 ;
        RECT 123.505 167.305 123.675 167.475 ;
        RECT 123.965 167.305 124.135 167.475 ;
        RECT 124.425 167.305 124.595 167.475 ;
        RECT 124.885 167.305 125.055 167.475 ;
        RECT 125.345 167.305 125.515 167.475 ;
        RECT 125.805 167.305 125.975 167.475 ;
        RECT 126.265 167.305 126.435 167.475 ;
        RECT 126.725 167.305 126.895 167.475 ;
        RECT 127.185 167.305 127.355 167.475 ;
        RECT 127.645 167.305 127.815 167.475 ;
        RECT 128.105 167.305 128.275 167.475 ;
        RECT 128.565 167.305 128.735 167.475 ;
        RECT 129.025 167.305 129.195 167.475 ;
        RECT 129.485 167.305 129.655 167.475 ;
        RECT 129.945 167.305 130.115 167.475 ;
        RECT 130.405 167.305 130.575 167.475 ;
        RECT 130.865 167.305 131.035 167.475 ;
        RECT 131.325 167.305 131.495 167.475 ;
        RECT 131.785 167.305 131.955 167.475 ;
        RECT 132.245 167.305 132.415 167.475 ;
        RECT 132.705 167.305 132.875 167.475 ;
        RECT 133.165 167.305 133.335 167.475 ;
        RECT 133.625 167.305 133.795 167.475 ;
        RECT 134.085 167.305 134.255 167.475 ;
        RECT 134.545 167.305 134.715 167.475 ;
        RECT 135.005 167.305 135.175 167.475 ;
        RECT 135.465 167.305 135.635 167.475 ;
        RECT 135.925 167.305 136.095 167.475 ;
        RECT 136.385 167.305 136.555 167.475 ;
        RECT 136.845 167.305 137.015 167.475 ;
        RECT 137.305 167.305 137.475 167.475 ;
        RECT 137.765 167.305 137.935 167.475 ;
        RECT 138.225 167.305 138.395 167.475 ;
        RECT 138.685 167.305 138.855 167.475 ;
        RECT 139.145 167.305 139.315 167.475 ;
        RECT 139.605 167.305 139.775 167.475 ;
        RECT 140.065 167.305 140.235 167.475 ;
        RECT 140.525 167.305 140.695 167.475 ;
        RECT 140.985 167.305 141.155 167.475 ;
        RECT 141.445 167.305 141.615 167.475 ;
        RECT 141.905 167.305 142.075 167.475 ;
        RECT 142.365 167.305 142.535 167.475 ;
        RECT 142.825 167.305 142.995 167.475 ;
        RECT 143.285 167.305 143.455 167.475 ;
        RECT 143.745 167.305 143.915 167.475 ;
        RECT 144.205 167.305 144.375 167.475 ;
        RECT 144.665 167.305 144.835 167.475 ;
        RECT 145.125 167.305 145.295 167.475 ;
        RECT 145.585 167.305 145.755 167.475 ;
        RECT 146.045 167.305 146.215 167.475 ;
        RECT 146.505 167.305 146.675 167.475 ;
        RECT 146.965 167.305 147.135 167.475 ;
        RECT 147.425 167.305 147.595 167.475 ;
        RECT 147.885 167.305 148.055 167.475 ;
        RECT 148.345 167.305 148.515 167.475 ;
        RECT 148.805 167.305 148.975 167.475 ;
        RECT 149.265 167.305 149.435 167.475 ;
        RECT 149.725 167.305 149.895 167.475 ;
        RECT 150.185 167.305 150.355 167.475 ;
        RECT 26.445 166.115 26.615 166.285 ;
        RECT 29.205 166.795 29.375 166.965 ;
        RECT 32.885 166.795 33.055 166.965 ;
        RECT 30.585 166.115 30.755 166.285 ;
        RECT 33.805 166.115 33.975 166.285 ;
        RECT 31.045 165.095 31.215 165.265 ;
        RECT 42.085 166.115 42.255 166.285 ;
        RECT 42.545 165.775 42.715 165.945 ;
        RECT 43.465 165.095 43.635 165.265 ;
        RECT 52.665 166.455 52.835 166.625 ;
        RECT 52.205 166.115 52.375 166.285 ;
        RECT 53.585 166.455 53.755 166.625 ;
        RECT 53.585 165.095 53.755 165.265 ;
        RECT 63.245 166.115 63.415 166.285 ;
        RECT 67.385 166.795 67.555 166.965 ;
        RECT 68.305 166.795 68.475 166.965 ;
        RECT 66.465 166.115 66.635 166.285 ;
        RECT 66.925 166.115 67.095 166.285 ;
        RECT 67.845 166.115 68.015 166.285 ;
        RECT 69.225 166.115 69.395 166.285 ;
        RECT 74.285 166.455 74.455 166.625 ;
        RECT 76.585 166.115 76.755 166.285 ;
        RECT 79.805 166.795 79.975 166.965 ;
        RECT 77.505 166.115 77.675 166.285 ;
        RECT 77.965 166.115 78.135 166.285 ;
        RECT 78.425 166.115 78.595 166.285 ;
        RECT 74.745 165.095 74.915 165.265 ;
        RECT 92.685 166.115 92.855 166.285 ;
        RECT 93.145 165.775 93.315 165.945 ;
        RECT 94.985 166.115 95.155 166.285 ;
        RECT 94.525 165.775 94.695 165.945 ;
        RECT 101.915 166.795 102.085 166.965 ;
        RECT 95.905 166.115 96.075 166.285 ;
        RECT 96.365 166.115 96.535 166.285 ;
        RECT 101.425 166.455 101.595 166.625 ;
        RECT 102.345 166.795 102.515 166.965 ;
        RECT 102.805 166.115 102.975 166.285 ;
        RECT 94.985 165.095 95.155 165.265 ;
        RECT 107.865 165.095 108.035 165.265 ;
        RECT 110.165 166.455 110.335 166.625 ;
        RECT 110.625 165.775 110.795 165.945 ;
        RECT 112.005 165.775 112.175 165.945 ;
        RECT 112.925 166.115 113.095 166.285 ;
        RECT 113.385 166.115 113.555 166.285 ;
        RECT 118.445 166.115 118.615 166.285 ;
        RECT 119.365 165.095 119.535 165.265 ;
        RECT 126.265 166.455 126.435 166.625 ;
        RECT 127.645 166.115 127.815 166.285 ;
        RECT 11.265 164.585 11.435 164.755 ;
        RECT 11.725 164.585 11.895 164.755 ;
        RECT 12.185 164.585 12.355 164.755 ;
        RECT 12.645 164.585 12.815 164.755 ;
        RECT 13.105 164.585 13.275 164.755 ;
        RECT 13.565 164.585 13.735 164.755 ;
        RECT 14.025 164.585 14.195 164.755 ;
        RECT 14.485 164.585 14.655 164.755 ;
        RECT 14.945 164.585 15.115 164.755 ;
        RECT 15.405 164.585 15.575 164.755 ;
        RECT 15.865 164.585 16.035 164.755 ;
        RECT 16.325 164.585 16.495 164.755 ;
        RECT 16.785 164.585 16.955 164.755 ;
        RECT 17.245 164.585 17.415 164.755 ;
        RECT 17.705 164.585 17.875 164.755 ;
        RECT 18.165 164.585 18.335 164.755 ;
        RECT 18.625 164.585 18.795 164.755 ;
        RECT 19.085 164.585 19.255 164.755 ;
        RECT 19.545 164.585 19.715 164.755 ;
        RECT 20.005 164.585 20.175 164.755 ;
        RECT 20.465 164.585 20.635 164.755 ;
        RECT 20.925 164.585 21.095 164.755 ;
        RECT 21.385 164.585 21.555 164.755 ;
        RECT 21.845 164.585 22.015 164.755 ;
        RECT 22.305 164.585 22.475 164.755 ;
        RECT 22.765 164.585 22.935 164.755 ;
        RECT 23.225 164.585 23.395 164.755 ;
        RECT 23.685 164.585 23.855 164.755 ;
        RECT 24.145 164.585 24.315 164.755 ;
        RECT 24.605 164.585 24.775 164.755 ;
        RECT 25.065 164.585 25.235 164.755 ;
        RECT 25.525 164.585 25.695 164.755 ;
        RECT 25.985 164.585 26.155 164.755 ;
        RECT 26.445 164.585 26.615 164.755 ;
        RECT 26.905 164.585 27.075 164.755 ;
        RECT 27.365 164.585 27.535 164.755 ;
        RECT 27.825 164.585 27.995 164.755 ;
        RECT 28.285 164.585 28.455 164.755 ;
        RECT 28.745 164.585 28.915 164.755 ;
        RECT 29.205 164.585 29.375 164.755 ;
        RECT 29.665 164.585 29.835 164.755 ;
        RECT 30.125 164.585 30.295 164.755 ;
        RECT 30.585 164.585 30.755 164.755 ;
        RECT 31.045 164.585 31.215 164.755 ;
        RECT 31.505 164.585 31.675 164.755 ;
        RECT 31.965 164.585 32.135 164.755 ;
        RECT 32.425 164.585 32.595 164.755 ;
        RECT 32.885 164.585 33.055 164.755 ;
        RECT 33.345 164.585 33.515 164.755 ;
        RECT 33.805 164.585 33.975 164.755 ;
        RECT 34.265 164.585 34.435 164.755 ;
        RECT 34.725 164.585 34.895 164.755 ;
        RECT 35.185 164.585 35.355 164.755 ;
        RECT 35.645 164.585 35.815 164.755 ;
        RECT 36.105 164.585 36.275 164.755 ;
        RECT 36.565 164.585 36.735 164.755 ;
        RECT 37.025 164.585 37.195 164.755 ;
        RECT 37.485 164.585 37.655 164.755 ;
        RECT 37.945 164.585 38.115 164.755 ;
        RECT 38.405 164.585 38.575 164.755 ;
        RECT 38.865 164.585 39.035 164.755 ;
        RECT 39.325 164.585 39.495 164.755 ;
        RECT 39.785 164.585 39.955 164.755 ;
        RECT 40.245 164.585 40.415 164.755 ;
        RECT 40.705 164.585 40.875 164.755 ;
        RECT 41.165 164.585 41.335 164.755 ;
        RECT 41.625 164.585 41.795 164.755 ;
        RECT 42.085 164.585 42.255 164.755 ;
        RECT 42.545 164.585 42.715 164.755 ;
        RECT 43.005 164.585 43.175 164.755 ;
        RECT 43.465 164.585 43.635 164.755 ;
        RECT 43.925 164.585 44.095 164.755 ;
        RECT 44.385 164.585 44.555 164.755 ;
        RECT 44.845 164.585 45.015 164.755 ;
        RECT 45.305 164.585 45.475 164.755 ;
        RECT 45.765 164.585 45.935 164.755 ;
        RECT 46.225 164.585 46.395 164.755 ;
        RECT 46.685 164.585 46.855 164.755 ;
        RECT 47.145 164.585 47.315 164.755 ;
        RECT 47.605 164.585 47.775 164.755 ;
        RECT 48.065 164.585 48.235 164.755 ;
        RECT 48.525 164.585 48.695 164.755 ;
        RECT 48.985 164.585 49.155 164.755 ;
        RECT 49.445 164.585 49.615 164.755 ;
        RECT 49.905 164.585 50.075 164.755 ;
        RECT 50.365 164.585 50.535 164.755 ;
        RECT 50.825 164.585 50.995 164.755 ;
        RECT 51.285 164.585 51.455 164.755 ;
        RECT 51.745 164.585 51.915 164.755 ;
        RECT 52.205 164.585 52.375 164.755 ;
        RECT 52.665 164.585 52.835 164.755 ;
        RECT 53.125 164.585 53.295 164.755 ;
        RECT 53.585 164.585 53.755 164.755 ;
        RECT 54.045 164.585 54.215 164.755 ;
        RECT 54.505 164.585 54.675 164.755 ;
        RECT 54.965 164.585 55.135 164.755 ;
        RECT 55.425 164.585 55.595 164.755 ;
        RECT 55.885 164.585 56.055 164.755 ;
        RECT 56.345 164.585 56.515 164.755 ;
        RECT 56.805 164.585 56.975 164.755 ;
        RECT 57.265 164.585 57.435 164.755 ;
        RECT 57.725 164.585 57.895 164.755 ;
        RECT 58.185 164.585 58.355 164.755 ;
        RECT 58.645 164.585 58.815 164.755 ;
        RECT 59.105 164.585 59.275 164.755 ;
        RECT 59.565 164.585 59.735 164.755 ;
        RECT 60.025 164.585 60.195 164.755 ;
        RECT 60.485 164.585 60.655 164.755 ;
        RECT 60.945 164.585 61.115 164.755 ;
        RECT 61.405 164.585 61.575 164.755 ;
        RECT 61.865 164.585 62.035 164.755 ;
        RECT 62.325 164.585 62.495 164.755 ;
        RECT 62.785 164.585 62.955 164.755 ;
        RECT 63.245 164.585 63.415 164.755 ;
        RECT 63.705 164.585 63.875 164.755 ;
        RECT 64.165 164.585 64.335 164.755 ;
        RECT 64.625 164.585 64.795 164.755 ;
        RECT 65.085 164.585 65.255 164.755 ;
        RECT 65.545 164.585 65.715 164.755 ;
        RECT 66.005 164.585 66.175 164.755 ;
        RECT 66.465 164.585 66.635 164.755 ;
        RECT 66.925 164.585 67.095 164.755 ;
        RECT 67.385 164.585 67.555 164.755 ;
        RECT 67.845 164.585 68.015 164.755 ;
        RECT 68.305 164.585 68.475 164.755 ;
        RECT 68.765 164.585 68.935 164.755 ;
        RECT 69.225 164.585 69.395 164.755 ;
        RECT 69.685 164.585 69.855 164.755 ;
        RECT 70.145 164.585 70.315 164.755 ;
        RECT 70.605 164.585 70.775 164.755 ;
        RECT 71.065 164.585 71.235 164.755 ;
        RECT 71.525 164.585 71.695 164.755 ;
        RECT 71.985 164.585 72.155 164.755 ;
        RECT 72.445 164.585 72.615 164.755 ;
        RECT 72.905 164.585 73.075 164.755 ;
        RECT 73.365 164.585 73.535 164.755 ;
        RECT 73.825 164.585 73.995 164.755 ;
        RECT 74.285 164.585 74.455 164.755 ;
        RECT 74.745 164.585 74.915 164.755 ;
        RECT 75.205 164.585 75.375 164.755 ;
        RECT 75.665 164.585 75.835 164.755 ;
        RECT 76.125 164.585 76.295 164.755 ;
        RECT 76.585 164.585 76.755 164.755 ;
        RECT 77.045 164.585 77.215 164.755 ;
        RECT 77.505 164.585 77.675 164.755 ;
        RECT 77.965 164.585 78.135 164.755 ;
        RECT 78.425 164.585 78.595 164.755 ;
        RECT 78.885 164.585 79.055 164.755 ;
        RECT 79.345 164.585 79.515 164.755 ;
        RECT 79.805 164.585 79.975 164.755 ;
        RECT 80.265 164.585 80.435 164.755 ;
        RECT 80.725 164.585 80.895 164.755 ;
        RECT 81.185 164.585 81.355 164.755 ;
        RECT 81.645 164.585 81.815 164.755 ;
        RECT 82.105 164.585 82.275 164.755 ;
        RECT 82.565 164.585 82.735 164.755 ;
        RECT 83.025 164.585 83.195 164.755 ;
        RECT 83.485 164.585 83.655 164.755 ;
        RECT 83.945 164.585 84.115 164.755 ;
        RECT 84.405 164.585 84.575 164.755 ;
        RECT 84.865 164.585 85.035 164.755 ;
        RECT 85.325 164.585 85.495 164.755 ;
        RECT 85.785 164.585 85.955 164.755 ;
        RECT 86.245 164.585 86.415 164.755 ;
        RECT 86.705 164.585 86.875 164.755 ;
        RECT 87.165 164.585 87.335 164.755 ;
        RECT 87.625 164.585 87.795 164.755 ;
        RECT 88.085 164.585 88.255 164.755 ;
        RECT 88.545 164.585 88.715 164.755 ;
        RECT 89.005 164.585 89.175 164.755 ;
        RECT 89.465 164.585 89.635 164.755 ;
        RECT 89.925 164.585 90.095 164.755 ;
        RECT 90.385 164.585 90.555 164.755 ;
        RECT 90.845 164.585 91.015 164.755 ;
        RECT 91.305 164.585 91.475 164.755 ;
        RECT 91.765 164.585 91.935 164.755 ;
        RECT 92.225 164.585 92.395 164.755 ;
        RECT 92.685 164.585 92.855 164.755 ;
        RECT 93.145 164.585 93.315 164.755 ;
        RECT 93.605 164.585 93.775 164.755 ;
        RECT 94.065 164.585 94.235 164.755 ;
        RECT 94.525 164.585 94.695 164.755 ;
        RECT 94.985 164.585 95.155 164.755 ;
        RECT 95.445 164.585 95.615 164.755 ;
        RECT 95.905 164.585 96.075 164.755 ;
        RECT 96.365 164.585 96.535 164.755 ;
        RECT 96.825 164.585 96.995 164.755 ;
        RECT 97.285 164.585 97.455 164.755 ;
        RECT 97.745 164.585 97.915 164.755 ;
        RECT 98.205 164.585 98.375 164.755 ;
        RECT 98.665 164.585 98.835 164.755 ;
        RECT 99.125 164.585 99.295 164.755 ;
        RECT 99.585 164.585 99.755 164.755 ;
        RECT 100.045 164.585 100.215 164.755 ;
        RECT 100.505 164.585 100.675 164.755 ;
        RECT 100.965 164.585 101.135 164.755 ;
        RECT 101.425 164.585 101.595 164.755 ;
        RECT 101.885 164.585 102.055 164.755 ;
        RECT 102.345 164.585 102.515 164.755 ;
        RECT 102.805 164.585 102.975 164.755 ;
        RECT 103.265 164.585 103.435 164.755 ;
        RECT 103.725 164.585 103.895 164.755 ;
        RECT 104.185 164.585 104.355 164.755 ;
        RECT 104.645 164.585 104.815 164.755 ;
        RECT 105.105 164.585 105.275 164.755 ;
        RECT 105.565 164.585 105.735 164.755 ;
        RECT 106.025 164.585 106.195 164.755 ;
        RECT 106.485 164.585 106.655 164.755 ;
        RECT 106.945 164.585 107.115 164.755 ;
        RECT 107.405 164.585 107.575 164.755 ;
        RECT 107.865 164.585 108.035 164.755 ;
        RECT 108.325 164.585 108.495 164.755 ;
        RECT 108.785 164.585 108.955 164.755 ;
        RECT 109.245 164.585 109.415 164.755 ;
        RECT 109.705 164.585 109.875 164.755 ;
        RECT 110.165 164.585 110.335 164.755 ;
        RECT 110.625 164.585 110.795 164.755 ;
        RECT 111.085 164.585 111.255 164.755 ;
        RECT 111.545 164.585 111.715 164.755 ;
        RECT 112.005 164.585 112.175 164.755 ;
        RECT 112.465 164.585 112.635 164.755 ;
        RECT 112.925 164.585 113.095 164.755 ;
        RECT 113.385 164.585 113.555 164.755 ;
        RECT 113.845 164.585 114.015 164.755 ;
        RECT 114.305 164.585 114.475 164.755 ;
        RECT 114.765 164.585 114.935 164.755 ;
        RECT 115.225 164.585 115.395 164.755 ;
        RECT 115.685 164.585 115.855 164.755 ;
        RECT 116.145 164.585 116.315 164.755 ;
        RECT 116.605 164.585 116.775 164.755 ;
        RECT 117.065 164.585 117.235 164.755 ;
        RECT 117.525 164.585 117.695 164.755 ;
        RECT 117.985 164.585 118.155 164.755 ;
        RECT 118.445 164.585 118.615 164.755 ;
        RECT 118.905 164.585 119.075 164.755 ;
        RECT 119.365 164.585 119.535 164.755 ;
        RECT 119.825 164.585 119.995 164.755 ;
        RECT 120.285 164.585 120.455 164.755 ;
        RECT 120.745 164.585 120.915 164.755 ;
        RECT 121.205 164.585 121.375 164.755 ;
        RECT 121.665 164.585 121.835 164.755 ;
        RECT 122.125 164.585 122.295 164.755 ;
        RECT 122.585 164.585 122.755 164.755 ;
        RECT 123.045 164.585 123.215 164.755 ;
        RECT 123.505 164.585 123.675 164.755 ;
        RECT 123.965 164.585 124.135 164.755 ;
        RECT 124.425 164.585 124.595 164.755 ;
        RECT 124.885 164.585 125.055 164.755 ;
        RECT 125.345 164.585 125.515 164.755 ;
        RECT 125.805 164.585 125.975 164.755 ;
        RECT 126.265 164.585 126.435 164.755 ;
        RECT 126.725 164.585 126.895 164.755 ;
        RECT 127.185 164.585 127.355 164.755 ;
        RECT 127.645 164.585 127.815 164.755 ;
        RECT 128.105 164.585 128.275 164.755 ;
        RECT 128.565 164.585 128.735 164.755 ;
        RECT 129.025 164.585 129.195 164.755 ;
        RECT 129.485 164.585 129.655 164.755 ;
        RECT 129.945 164.585 130.115 164.755 ;
        RECT 130.405 164.585 130.575 164.755 ;
        RECT 130.865 164.585 131.035 164.755 ;
        RECT 131.325 164.585 131.495 164.755 ;
        RECT 131.785 164.585 131.955 164.755 ;
        RECT 132.245 164.585 132.415 164.755 ;
        RECT 132.705 164.585 132.875 164.755 ;
        RECT 133.165 164.585 133.335 164.755 ;
        RECT 133.625 164.585 133.795 164.755 ;
        RECT 134.085 164.585 134.255 164.755 ;
        RECT 134.545 164.585 134.715 164.755 ;
        RECT 135.005 164.585 135.175 164.755 ;
        RECT 135.465 164.585 135.635 164.755 ;
        RECT 135.925 164.585 136.095 164.755 ;
        RECT 136.385 164.585 136.555 164.755 ;
        RECT 136.845 164.585 137.015 164.755 ;
        RECT 137.305 164.585 137.475 164.755 ;
        RECT 137.765 164.585 137.935 164.755 ;
        RECT 138.225 164.585 138.395 164.755 ;
        RECT 138.685 164.585 138.855 164.755 ;
        RECT 139.145 164.585 139.315 164.755 ;
        RECT 139.605 164.585 139.775 164.755 ;
        RECT 140.065 164.585 140.235 164.755 ;
        RECT 140.525 164.585 140.695 164.755 ;
        RECT 140.985 164.585 141.155 164.755 ;
        RECT 141.445 164.585 141.615 164.755 ;
        RECT 141.905 164.585 142.075 164.755 ;
        RECT 142.365 164.585 142.535 164.755 ;
        RECT 142.825 164.585 142.995 164.755 ;
        RECT 143.285 164.585 143.455 164.755 ;
        RECT 143.745 164.585 143.915 164.755 ;
        RECT 144.205 164.585 144.375 164.755 ;
        RECT 144.665 164.585 144.835 164.755 ;
        RECT 145.125 164.585 145.295 164.755 ;
        RECT 145.585 164.585 145.755 164.755 ;
        RECT 146.045 164.585 146.215 164.755 ;
        RECT 146.505 164.585 146.675 164.755 ;
        RECT 146.965 164.585 147.135 164.755 ;
        RECT 147.425 164.585 147.595 164.755 ;
        RECT 147.885 164.585 148.055 164.755 ;
        RECT 148.345 164.585 148.515 164.755 ;
        RECT 148.805 164.585 148.975 164.755 ;
        RECT 149.265 164.585 149.435 164.755 ;
        RECT 149.725 164.585 149.895 164.755 ;
        RECT 150.185 164.585 150.355 164.755 ;
        RECT 16.810 163.735 16.980 163.905 ;
        RECT 16.325 163.055 16.495 163.225 ;
        RECT 17.205 163.395 17.375 163.565 ;
        RECT 17.660 163.055 17.830 163.225 ;
        RECT 18.910 163.735 19.080 163.905 ;
        RECT 18.395 163.395 18.565 163.565 ;
        RECT 20.480 163.735 20.650 163.905 ;
        RECT 20.915 163.395 21.085 163.565 ;
        RECT 23.225 164.075 23.395 164.245 ;
        RECT 30.585 163.395 30.755 163.565 ;
        RECT 30.125 163.055 30.295 163.225 ;
        RECT 31.965 162.375 32.135 162.545 ;
        RECT 32.885 163.395 33.055 163.565 ;
        RECT 33.345 163.055 33.515 163.225 ;
        RECT 35.185 163.735 35.355 163.905 ;
        RECT 37.945 163.395 38.115 163.565 ;
        RECT 38.865 162.375 39.035 162.545 ;
        RECT 39.325 162.715 39.495 162.885 ;
        RECT 39.785 163.055 39.955 163.225 ;
        RECT 41.625 163.055 41.795 163.225 ;
        RECT 40.705 162.715 40.875 162.885 ;
        RECT 43.005 163.055 43.175 163.225 ;
        RECT 44.050 163.395 44.220 163.565 ;
        RECT 44.845 163.735 45.015 163.905 ;
        RECT 48.065 163.395 48.235 163.565 ;
        RECT 47.605 163.055 47.775 163.225 ;
        RECT 49.445 162.375 49.615 162.545 ;
        RECT 52.205 163.395 52.375 163.565 ;
        RECT 52.665 163.055 52.835 163.225 ;
        RECT 53.125 163.395 53.295 163.565 ;
        RECT 53.585 163.055 53.755 163.225 ;
        RECT 54.965 163.055 55.135 163.225 ;
        RECT 54.505 162.375 54.675 162.545 ;
        RECT 55.885 162.715 56.055 162.885 ;
        RECT 56.345 163.055 56.515 163.225 ;
        RECT 56.805 163.055 56.975 163.225 ;
        RECT 66.925 163.055 67.095 163.225 ;
        RECT 68.765 164.075 68.935 164.245 ;
        RECT 69.685 164.075 69.855 164.245 ;
        RECT 57.725 162.375 57.895 162.545 ;
        RECT 68.765 162.375 68.935 162.545 ;
        RECT 74.395 164.075 74.565 164.245 ;
        RECT 75.205 164.075 75.375 164.245 ;
        RECT 71.065 162.715 71.235 162.885 ;
        RECT 71.985 162.715 72.155 162.885 ;
        RECT 73.365 162.715 73.535 162.885 ;
        RECT 70.145 162.375 70.315 162.545 ;
        RECT 74.365 162.715 74.535 162.885 ;
        RECT 82.565 164.075 82.735 164.245 ;
        RECT 76.125 163.055 76.295 163.225 ;
        RECT 85.325 162.375 85.495 162.545 ;
        RECT 87.635 163.395 87.805 163.565 ;
        RECT 88.070 163.735 88.240 163.905 ;
        RECT 89.640 163.735 89.810 163.905 ;
        RECT 90.155 163.395 90.325 163.565 ;
        RECT 90.890 162.715 91.060 162.885 ;
        RECT 91.345 163.395 91.515 163.565 ;
        RECT 91.740 163.735 91.910 163.905 ;
        RECT 92.685 163.735 92.855 163.905 ;
        RECT 92.225 163.395 92.395 163.565 ;
        RECT 95.445 164.075 95.615 164.245 ;
        RECT 93.605 163.055 93.775 163.225 ;
        RECT 94.525 163.055 94.695 163.225 ;
        RECT 94.985 163.055 95.155 163.225 ;
        RECT 95.905 163.055 96.075 163.225 ;
        RECT 106.025 163.055 106.195 163.225 ;
        RECT 106.945 163.055 107.115 163.225 ;
        RECT 106.485 162.375 106.655 162.545 ;
        RECT 11.265 161.865 11.435 162.035 ;
        RECT 11.725 161.865 11.895 162.035 ;
        RECT 12.185 161.865 12.355 162.035 ;
        RECT 12.645 161.865 12.815 162.035 ;
        RECT 13.105 161.865 13.275 162.035 ;
        RECT 13.565 161.865 13.735 162.035 ;
        RECT 14.025 161.865 14.195 162.035 ;
        RECT 14.485 161.865 14.655 162.035 ;
        RECT 14.945 161.865 15.115 162.035 ;
        RECT 15.405 161.865 15.575 162.035 ;
        RECT 15.865 161.865 16.035 162.035 ;
        RECT 16.325 161.865 16.495 162.035 ;
        RECT 16.785 161.865 16.955 162.035 ;
        RECT 17.245 161.865 17.415 162.035 ;
        RECT 17.705 161.865 17.875 162.035 ;
        RECT 18.165 161.865 18.335 162.035 ;
        RECT 18.625 161.865 18.795 162.035 ;
        RECT 19.085 161.865 19.255 162.035 ;
        RECT 19.545 161.865 19.715 162.035 ;
        RECT 20.005 161.865 20.175 162.035 ;
        RECT 20.465 161.865 20.635 162.035 ;
        RECT 20.925 161.865 21.095 162.035 ;
        RECT 21.385 161.865 21.555 162.035 ;
        RECT 21.845 161.865 22.015 162.035 ;
        RECT 22.305 161.865 22.475 162.035 ;
        RECT 22.765 161.865 22.935 162.035 ;
        RECT 23.225 161.865 23.395 162.035 ;
        RECT 23.685 161.865 23.855 162.035 ;
        RECT 24.145 161.865 24.315 162.035 ;
        RECT 24.605 161.865 24.775 162.035 ;
        RECT 25.065 161.865 25.235 162.035 ;
        RECT 25.525 161.865 25.695 162.035 ;
        RECT 25.985 161.865 26.155 162.035 ;
        RECT 26.445 161.865 26.615 162.035 ;
        RECT 26.905 161.865 27.075 162.035 ;
        RECT 27.365 161.865 27.535 162.035 ;
        RECT 27.825 161.865 27.995 162.035 ;
        RECT 28.285 161.865 28.455 162.035 ;
        RECT 28.745 161.865 28.915 162.035 ;
        RECT 29.205 161.865 29.375 162.035 ;
        RECT 29.665 161.865 29.835 162.035 ;
        RECT 30.125 161.865 30.295 162.035 ;
        RECT 30.585 161.865 30.755 162.035 ;
        RECT 31.045 161.865 31.215 162.035 ;
        RECT 31.505 161.865 31.675 162.035 ;
        RECT 31.965 161.865 32.135 162.035 ;
        RECT 32.425 161.865 32.595 162.035 ;
        RECT 32.885 161.865 33.055 162.035 ;
        RECT 33.345 161.865 33.515 162.035 ;
        RECT 33.805 161.865 33.975 162.035 ;
        RECT 34.265 161.865 34.435 162.035 ;
        RECT 34.725 161.865 34.895 162.035 ;
        RECT 35.185 161.865 35.355 162.035 ;
        RECT 35.645 161.865 35.815 162.035 ;
        RECT 36.105 161.865 36.275 162.035 ;
        RECT 36.565 161.865 36.735 162.035 ;
        RECT 37.025 161.865 37.195 162.035 ;
        RECT 37.485 161.865 37.655 162.035 ;
        RECT 37.945 161.865 38.115 162.035 ;
        RECT 38.405 161.865 38.575 162.035 ;
        RECT 38.865 161.865 39.035 162.035 ;
        RECT 39.325 161.865 39.495 162.035 ;
        RECT 39.785 161.865 39.955 162.035 ;
        RECT 40.245 161.865 40.415 162.035 ;
        RECT 40.705 161.865 40.875 162.035 ;
        RECT 41.165 161.865 41.335 162.035 ;
        RECT 41.625 161.865 41.795 162.035 ;
        RECT 42.085 161.865 42.255 162.035 ;
        RECT 42.545 161.865 42.715 162.035 ;
        RECT 43.005 161.865 43.175 162.035 ;
        RECT 43.465 161.865 43.635 162.035 ;
        RECT 43.925 161.865 44.095 162.035 ;
        RECT 44.385 161.865 44.555 162.035 ;
        RECT 44.845 161.865 45.015 162.035 ;
        RECT 45.305 161.865 45.475 162.035 ;
        RECT 45.765 161.865 45.935 162.035 ;
        RECT 46.225 161.865 46.395 162.035 ;
        RECT 46.685 161.865 46.855 162.035 ;
        RECT 47.145 161.865 47.315 162.035 ;
        RECT 47.605 161.865 47.775 162.035 ;
        RECT 48.065 161.865 48.235 162.035 ;
        RECT 48.525 161.865 48.695 162.035 ;
        RECT 48.985 161.865 49.155 162.035 ;
        RECT 49.445 161.865 49.615 162.035 ;
        RECT 49.905 161.865 50.075 162.035 ;
        RECT 50.365 161.865 50.535 162.035 ;
        RECT 50.825 161.865 50.995 162.035 ;
        RECT 51.285 161.865 51.455 162.035 ;
        RECT 51.745 161.865 51.915 162.035 ;
        RECT 52.205 161.865 52.375 162.035 ;
        RECT 52.665 161.865 52.835 162.035 ;
        RECT 53.125 161.865 53.295 162.035 ;
        RECT 53.585 161.865 53.755 162.035 ;
        RECT 54.045 161.865 54.215 162.035 ;
        RECT 54.505 161.865 54.675 162.035 ;
        RECT 54.965 161.865 55.135 162.035 ;
        RECT 55.425 161.865 55.595 162.035 ;
        RECT 55.885 161.865 56.055 162.035 ;
        RECT 56.345 161.865 56.515 162.035 ;
        RECT 56.805 161.865 56.975 162.035 ;
        RECT 57.265 161.865 57.435 162.035 ;
        RECT 57.725 161.865 57.895 162.035 ;
        RECT 58.185 161.865 58.355 162.035 ;
        RECT 58.645 161.865 58.815 162.035 ;
        RECT 59.105 161.865 59.275 162.035 ;
        RECT 59.565 161.865 59.735 162.035 ;
        RECT 60.025 161.865 60.195 162.035 ;
        RECT 60.485 161.865 60.655 162.035 ;
        RECT 60.945 161.865 61.115 162.035 ;
        RECT 61.405 161.865 61.575 162.035 ;
        RECT 61.865 161.865 62.035 162.035 ;
        RECT 62.325 161.865 62.495 162.035 ;
        RECT 62.785 161.865 62.955 162.035 ;
        RECT 63.245 161.865 63.415 162.035 ;
        RECT 63.705 161.865 63.875 162.035 ;
        RECT 64.165 161.865 64.335 162.035 ;
        RECT 64.625 161.865 64.795 162.035 ;
        RECT 65.085 161.865 65.255 162.035 ;
        RECT 65.545 161.865 65.715 162.035 ;
        RECT 66.005 161.865 66.175 162.035 ;
        RECT 66.465 161.865 66.635 162.035 ;
        RECT 66.925 161.865 67.095 162.035 ;
        RECT 67.385 161.865 67.555 162.035 ;
        RECT 67.845 161.865 68.015 162.035 ;
        RECT 68.305 161.865 68.475 162.035 ;
        RECT 68.765 161.865 68.935 162.035 ;
        RECT 69.225 161.865 69.395 162.035 ;
        RECT 69.685 161.865 69.855 162.035 ;
        RECT 70.145 161.865 70.315 162.035 ;
        RECT 70.605 161.865 70.775 162.035 ;
        RECT 71.065 161.865 71.235 162.035 ;
        RECT 71.525 161.865 71.695 162.035 ;
        RECT 71.985 161.865 72.155 162.035 ;
        RECT 72.445 161.865 72.615 162.035 ;
        RECT 72.905 161.865 73.075 162.035 ;
        RECT 73.365 161.865 73.535 162.035 ;
        RECT 73.825 161.865 73.995 162.035 ;
        RECT 74.285 161.865 74.455 162.035 ;
        RECT 74.745 161.865 74.915 162.035 ;
        RECT 75.205 161.865 75.375 162.035 ;
        RECT 75.665 161.865 75.835 162.035 ;
        RECT 76.125 161.865 76.295 162.035 ;
        RECT 76.585 161.865 76.755 162.035 ;
        RECT 77.045 161.865 77.215 162.035 ;
        RECT 77.505 161.865 77.675 162.035 ;
        RECT 77.965 161.865 78.135 162.035 ;
        RECT 78.425 161.865 78.595 162.035 ;
        RECT 78.885 161.865 79.055 162.035 ;
        RECT 79.345 161.865 79.515 162.035 ;
        RECT 79.805 161.865 79.975 162.035 ;
        RECT 80.265 161.865 80.435 162.035 ;
        RECT 80.725 161.865 80.895 162.035 ;
        RECT 81.185 161.865 81.355 162.035 ;
        RECT 81.645 161.865 81.815 162.035 ;
        RECT 82.105 161.865 82.275 162.035 ;
        RECT 82.565 161.865 82.735 162.035 ;
        RECT 83.025 161.865 83.195 162.035 ;
        RECT 83.485 161.865 83.655 162.035 ;
        RECT 83.945 161.865 84.115 162.035 ;
        RECT 84.405 161.865 84.575 162.035 ;
        RECT 84.865 161.865 85.035 162.035 ;
        RECT 85.325 161.865 85.495 162.035 ;
        RECT 85.785 161.865 85.955 162.035 ;
        RECT 86.245 161.865 86.415 162.035 ;
        RECT 86.705 161.865 86.875 162.035 ;
        RECT 87.165 161.865 87.335 162.035 ;
        RECT 87.625 161.865 87.795 162.035 ;
        RECT 88.085 161.865 88.255 162.035 ;
        RECT 88.545 161.865 88.715 162.035 ;
        RECT 89.005 161.865 89.175 162.035 ;
        RECT 89.465 161.865 89.635 162.035 ;
        RECT 89.925 161.865 90.095 162.035 ;
        RECT 90.385 161.865 90.555 162.035 ;
        RECT 90.845 161.865 91.015 162.035 ;
        RECT 91.305 161.865 91.475 162.035 ;
        RECT 91.765 161.865 91.935 162.035 ;
        RECT 92.225 161.865 92.395 162.035 ;
        RECT 92.685 161.865 92.855 162.035 ;
        RECT 93.145 161.865 93.315 162.035 ;
        RECT 93.605 161.865 93.775 162.035 ;
        RECT 94.065 161.865 94.235 162.035 ;
        RECT 94.525 161.865 94.695 162.035 ;
        RECT 94.985 161.865 95.155 162.035 ;
        RECT 95.445 161.865 95.615 162.035 ;
        RECT 95.905 161.865 96.075 162.035 ;
        RECT 96.365 161.865 96.535 162.035 ;
        RECT 96.825 161.865 96.995 162.035 ;
        RECT 97.285 161.865 97.455 162.035 ;
        RECT 97.745 161.865 97.915 162.035 ;
        RECT 98.205 161.865 98.375 162.035 ;
        RECT 98.665 161.865 98.835 162.035 ;
        RECT 99.125 161.865 99.295 162.035 ;
        RECT 99.585 161.865 99.755 162.035 ;
        RECT 100.045 161.865 100.215 162.035 ;
        RECT 100.505 161.865 100.675 162.035 ;
        RECT 100.965 161.865 101.135 162.035 ;
        RECT 101.425 161.865 101.595 162.035 ;
        RECT 101.885 161.865 102.055 162.035 ;
        RECT 102.345 161.865 102.515 162.035 ;
        RECT 102.805 161.865 102.975 162.035 ;
        RECT 103.265 161.865 103.435 162.035 ;
        RECT 103.725 161.865 103.895 162.035 ;
        RECT 104.185 161.865 104.355 162.035 ;
        RECT 104.645 161.865 104.815 162.035 ;
        RECT 105.105 161.865 105.275 162.035 ;
        RECT 105.565 161.865 105.735 162.035 ;
        RECT 106.025 161.865 106.195 162.035 ;
        RECT 106.485 161.865 106.655 162.035 ;
        RECT 106.945 161.865 107.115 162.035 ;
        RECT 107.405 161.865 107.575 162.035 ;
        RECT 107.865 161.865 108.035 162.035 ;
        RECT 108.325 161.865 108.495 162.035 ;
        RECT 108.785 161.865 108.955 162.035 ;
        RECT 109.245 161.865 109.415 162.035 ;
        RECT 109.705 161.865 109.875 162.035 ;
        RECT 110.165 161.865 110.335 162.035 ;
        RECT 110.625 161.865 110.795 162.035 ;
        RECT 111.085 161.865 111.255 162.035 ;
        RECT 111.545 161.865 111.715 162.035 ;
        RECT 112.005 161.865 112.175 162.035 ;
        RECT 112.465 161.865 112.635 162.035 ;
        RECT 112.925 161.865 113.095 162.035 ;
        RECT 113.385 161.865 113.555 162.035 ;
        RECT 113.845 161.865 114.015 162.035 ;
        RECT 114.305 161.865 114.475 162.035 ;
        RECT 114.765 161.865 114.935 162.035 ;
        RECT 115.225 161.865 115.395 162.035 ;
        RECT 115.685 161.865 115.855 162.035 ;
        RECT 116.145 161.865 116.315 162.035 ;
        RECT 116.605 161.865 116.775 162.035 ;
        RECT 117.065 161.865 117.235 162.035 ;
        RECT 117.525 161.865 117.695 162.035 ;
        RECT 117.985 161.865 118.155 162.035 ;
        RECT 118.445 161.865 118.615 162.035 ;
        RECT 118.905 161.865 119.075 162.035 ;
        RECT 119.365 161.865 119.535 162.035 ;
        RECT 119.825 161.865 119.995 162.035 ;
        RECT 120.285 161.865 120.455 162.035 ;
        RECT 120.745 161.865 120.915 162.035 ;
        RECT 121.205 161.865 121.375 162.035 ;
        RECT 121.665 161.865 121.835 162.035 ;
        RECT 122.125 161.865 122.295 162.035 ;
        RECT 122.585 161.865 122.755 162.035 ;
        RECT 123.045 161.865 123.215 162.035 ;
        RECT 123.505 161.865 123.675 162.035 ;
        RECT 123.965 161.865 124.135 162.035 ;
        RECT 124.425 161.865 124.595 162.035 ;
        RECT 124.885 161.865 125.055 162.035 ;
        RECT 125.345 161.865 125.515 162.035 ;
        RECT 125.805 161.865 125.975 162.035 ;
        RECT 126.265 161.865 126.435 162.035 ;
        RECT 126.725 161.865 126.895 162.035 ;
        RECT 127.185 161.865 127.355 162.035 ;
        RECT 127.645 161.865 127.815 162.035 ;
        RECT 128.105 161.865 128.275 162.035 ;
        RECT 128.565 161.865 128.735 162.035 ;
        RECT 129.025 161.865 129.195 162.035 ;
        RECT 129.485 161.865 129.655 162.035 ;
        RECT 129.945 161.865 130.115 162.035 ;
        RECT 130.405 161.865 130.575 162.035 ;
        RECT 130.865 161.865 131.035 162.035 ;
        RECT 131.325 161.865 131.495 162.035 ;
        RECT 131.785 161.865 131.955 162.035 ;
        RECT 132.245 161.865 132.415 162.035 ;
        RECT 132.705 161.865 132.875 162.035 ;
        RECT 133.165 161.865 133.335 162.035 ;
        RECT 133.625 161.865 133.795 162.035 ;
        RECT 134.085 161.865 134.255 162.035 ;
        RECT 134.545 161.865 134.715 162.035 ;
        RECT 135.005 161.865 135.175 162.035 ;
        RECT 135.465 161.865 135.635 162.035 ;
        RECT 135.925 161.865 136.095 162.035 ;
        RECT 136.385 161.865 136.555 162.035 ;
        RECT 136.845 161.865 137.015 162.035 ;
        RECT 137.305 161.865 137.475 162.035 ;
        RECT 137.765 161.865 137.935 162.035 ;
        RECT 138.225 161.865 138.395 162.035 ;
        RECT 138.685 161.865 138.855 162.035 ;
        RECT 139.145 161.865 139.315 162.035 ;
        RECT 139.605 161.865 139.775 162.035 ;
        RECT 140.065 161.865 140.235 162.035 ;
        RECT 140.525 161.865 140.695 162.035 ;
        RECT 140.985 161.865 141.155 162.035 ;
        RECT 141.445 161.865 141.615 162.035 ;
        RECT 141.905 161.865 142.075 162.035 ;
        RECT 142.365 161.865 142.535 162.035 ;
        RECT 142.825 161.865 142.995 162.035 ;
        RECT 143.285 161.865 143.455 162.035 ;
        RECT 143.745 161.865 143.915 162.035 ;
        RECT 144.205 161.865 144.375 162.035 ;
        RECT 144.665 161.865 144.835 162.035 ;
        RECT 145.125 161.865 145.295 162.035 ;
        RECT 145.585 161.865 145.755 162.035 ;
        RECT 146.045 161.865 146.215 162.035 ;
        RECT 146.505 161.865 146.675 162.035 ;
        RECT 146.965 161.865 147.135 162.035 ;
        RECT 147.425 161.865 147.595 162.035 ;
        RECT 147.885 161.865 148.055 162.035 ;
        RECT 148.345 161.865 148.515 162.035 ;
        RECT 148.805 161.865 148.975 162.035 ;
        RECT 149.265 161.865 149.435 162.035 ;
        RECT 149.725 161.865 149.895 162.035 ;
        RECT 150.185 161.865 150.355 162.035 ;
        RECT 23.225 160.335 23.395 160.505 ;
        RECT 23.710 159.995 23.880 160.165 ;
        RECT 24.105 160.335 24.275 160.505 ;
        RECT 24.560 160.675 24.730 160.845 ;
        RECT 25.295 160.335 25.465 160.505 ;
        RECT 25.810 159.995 25.980 160.165 ;
        RECT 27.380 159.995 27.550 160.165 ;
        RECT 27.815 160.335 27.985 160.505 ;
        RECT 30.125 159.655 30.295 159.825 ;
        RECT 37.945 160.675 38.115 160.845 ;
        RECT 38.405 160.675 38.575 160.845 ;
        RECT 40.245 160.675 40.415 160.845 ;
        RECT 44.385 161.355 44.555 161.525 ;
        RECT 44.845 160.675 45.015 160.845 ;
        RECT 41.165 159.995 41.335 160.165 ;
        RECT 49.905 160.675 50.075 160.845 ;
        RECT 53.125 161.355 53.295 161.525 ;
        RECT 52.205 160.675 52.375 160.845 ;
        RECT 51.285 160.335 51.455 160.505 ;
        RECT 52.205 159.655 52.375 159.825 ;
        RECT 55.425 159.995 55.595 160.165 ;
        RECT 57.735 160.335 57.905 160.505 ;
        RECT 58.170 159.995 58.340 160.165 ;
        RECT 60.255 160.335 60.425 160.505 ;
        RECT 59.740 159.995 59.910 160.165 ;
        RECT 61.100 161.015 61.270 161.185 ;
        RECT 61.445 160.335 61.615 160.505 ;
        RECT 63.245 161.355 63.415 161.525 ;
        RECT 62.325 160.335 62.495 160.505 ;
        RECT 61.840 159.995 62.010 160.165 ;
        RECT 64.165 160.675 64.335 160.845 ;
        RECT 66.925 160.675 67.095 160.845 ;
        RECT 68.305 160.675 68.475 160.845 ;
        RECT 69.225 160.675 69.395 160.845 ;
        RECT 70.145 160.675 70.315 160.845 ;
        RECT 66.005 159.655 66.175 159.825 ;
        RECT 73.365 160.335 73.535 160.505 ;
        RECT 73.825 159.995 73.995 160.165 ;
        RECT 74.745 160.335 74.915 160.505 ;
        RECT 75.205 160.675 75.375 160.845 ;
        RECT 75.665 160.675 75.835 160.845 ;
        RECT 76.125 160.335 76.295 160.505 ;
        RECT 77.045 160.675 77.215 160.845 ;
        RECT 78.885 161.355 79.055 161.525 ;
        RECT 79.805 159.995 79.975 160.165 ;
        RECT 78.885 159.655 79.055 159.825 ;
        RECT 80.265 161.355 80.435 161.525 ;
        RECT 81.185 160.335 81.355 160.505 ;
        RECT 81.645 160.335 81.815 160.505 ;
        RECT 82.105 160.675 82.275 160.845 ;
        RECT 82.565 160.675 82.735 160.845 ;
        RECT 83.485 160.675 83.655 160.845 ;
        RECT 89.005 160.675 89.175 160.845 ;
        RECT 84.405 159.995 84.575 160.165 ;
        RECT 91.765 160.675 91.935 160.845 ;
        RECT 96.825 160.675 96.995 160.845 ;
        RECT 97.310 159.995 97.480 160.165 ;
        RECT 97.705 160.335 97.875 160.505 ;
        RECT 98.105 160.675 98.275 160.845 ;
        RECT 98.895 160.335 99.065 160.505 ;
        RECT 99.410 159.995 99.580 160.165 ;
        RECT 100.980 159.995 101.150 160.165 ;
        RECT 101.415 160.335 101.585 160.505 ;
        RECT 103.725 161.355 103.895 161.525 ;
        RECT 106.485 160.675 106.655 160.845 ;
        RECT 106.970 159.995 107.140 160.165 ;
        RECT 107.365 160.335 107.535 160.505 ;
        RECT 107.710 161.015 107.880 161.185 ;
        RECT 108.555 160.335 108.725 160.505 ;
        RECT 109.070 159.995 109.240 160.165 ;
        RECT 110.640 159.995 110.810 160.165 ;
        RECT 111.075 160.335 111.245 160.505 ;
        RECT 113.385 161.355 113.555 161.525 ;
        RECT 11.265 159.145 11.435 159.315 ;
        RECT 11.725 159.145 11.895 159.315 ;
        RECT 12.185 159.145 12.355 159.315 ;
        RECT 12.645 159.145 12.815 159.315 ;
        RECT 13.105 159.145 13.275 159.315 ;
        RECT 13.565 159.145 13.735 159.315 ;
        RECT 14.025 159.145 14.195 159.315 ;
        RECT 14.485 159.145 14.655 159.315 ;
        RECT 14.945 159.145 15.115 159.315 ;
        RECT 15.405 159.145 15.575 159.315 ;
        RECT 15.865 159.145 16.035 159.315 ;
        RECT 16.325 159.145 16.495 159.315 ;
        RECT 16.785 159.145 16.955 159.315 ;
        RECT 17.245 159.145 17.415 159.315 ;
        RECT 17.705 159.145 17.875 159.315 ;
        RECT 18.165 159.145 18.335 159.315 ;
        RECT 18.625 159.145 18.795 159.315 ;
        RECT 19.085 159.145 19.255 159.315 ;
        RECT 19.545 159.145 19.715 159.315 ;
        RECT 20.005 159.145 20.175 159.315 ;
        RECT 20.465 159.145 20.635 159.315 ;
        RECT 20.925 159.145 21.095 159.315 ;
        RECT 21.385 159.145 21.555 159.315 ;
        RECT 21.845 159.145 22.015 159.315 ;
        RECT 22.305 159.145 22.475 159.315 ;
        RECT 22.765 159.145 22.935 159.315 ;
        RECT 23.225 159.145 23.395 159.315 ;
        RECT 23.685 159.145 23.855 159.315 ;
        RECT 24.145 159.145 24.315 159.315 ;
        RECT 24.605 159.145 24.775 159.315 ;
        RECT 25.065 159.145 25.235 159.315 ;
        RECT 25.525 159.145 25.695 159.315 ;
        RECT 25.985 159.145 26.155 159.315 ;
        RECT 26.445 159.145 26.615 159.315 ;
        RECT 26.905 159.145 27.075 159.315 ;
        RECT 27.365 159.145 27.535 159.315 ;
        RECT 27.825 159.145 27.995 159.315 ;
        RECT 28.285 159.145 28.455 159.315 ;
        RECT 28.745 159.145 28.915 159.315 ;
        RECT 29.205 159.145 29.375 159.315 ;
        RECT 29.665 159.145 29.835 159.315 ;
        RECT 30.125 159.145 30.295 159.315 ;
        RECT 30.585 159.145 30.755 159.315 ;
        RECT 31.045 159.145 31.215 159.315 ;
        RECT 31.505 159.145 31.675 159.315 ;
        RECT 31.965 159.145 32.135 159.315 ;
        RECT 32.425 159.145 32.595 159.315 ;
        RECT 32.885 159.145 33.055 159.315 ;
        RECT 33.345 159.145 33.515 159.315 ;
        RECT 33.805 159.145 33.975 159.315 ;
        RECT 34.265 159.145 34.435 159.315 ;
        RECT 34.725 159.145 34.895 159.315 ;
        RECT 35.185 159.145 35.355 159.315 ;
        RECT 35.645 159.145 35.815 159.315 ;
        RECT 36.105 159.145 36.275 159.315 ;
        RECT 36.565 159.145 36.735 159.315 ;
        RECT 37.025 159.145 37.195 159.315 ;
        RECT 37.485 159.145 37.655 159.315 ;
        RECT 37.945 159.145 38.115 159.315 ;
        RECT 38.405 159.145 38.575 159.315 ;
        RECT 38.865 159.145 39.035 159.315 ;
        RECT 39.325 159.145 39.495 159.315 ;
        RECT 39.785 159.145 39.955 159.315 ;
        RECT 40.245 159.145 40.415 159.315 ;
        RECT 40.705 159.145 40.875 159.315 ;
        RECT 41.165 159.145 41.335 159.315 ;
        RECT 41.625 159.145 41.795 159.315 ;
        RECT 42.085 159.145 42.255 159.315 ;
        RECT 42.545 159.145 42.715 159.315 ;
        RECT 43.005 159.145 43.175 159.315 ;
        RECT 43.465 159.145 43.635 159.315 ;
        RECT 43.925 159.145 44.095 159.315 ;
        RECT 44.385 159.145 44.555 159.315 ;
        RECT 44.845 159.145 45.015 159.315 ;
        RECT 45.305 159.145 45.475 159.315 ;
        RECT 45.765 159.145 45.935 159.315 ;
        RECT 46.225 159.145 46.395 159.315 ;
        RECT 46.685 159.145 46.855 159.315 ;
        RECT 47.145 159.145 47.315 159.315 ;
        RECT 47.605 159.145 47.775 159.315 ;
        RECT 48.065 159.145 48.235 159.315 ;
        RECT 48.525 159.145 48.695 159.315 ;
        RECT 48.985 159.145 49.155 159.315 ;
        RECT 49.445 159.145 49.615 159.315 ;
        RECT 49.905 159.145 50.075 159.315 ;
        RECT 50.365 159.145 50.535 159.315 ;
        RECT 50.825 159.145 50.995 159.315 ;
        RECT 51.285 159.145 51.455 159.315 ;
        RECT 51.745 159.145 51.915 159.315 ;
        RECT 52.205 159.145 52.375 159.315 ;
        RECT 52.665 159.145 52.835 159.315 ;
        RECT 53.125 159.145 53.295 159.315 ;
        RECT 53.585 159.145 53.755 159.315 ;
        RECT 54.045 159.145 54.215 159.315 ;
        RECT 54.505 159.145 54.675 159.315 ;
        RECT 54.965 159.145 55.135 159.315 ;
        RECT 55.425 159.145 55.595 159.315 ;
        RECT 55.885 159.145 56.055 159.315 ;
        RECT 56.345 159.145 56.515 159.315 ;
        RECT 56.805 159.145 56.975 159.315 ;
        RECT 57.265 159.145 57.435 159.315 ;
        RECT 57.725 159.145 57.895 159.315 ;
        RECT 58.185 159.145 58.355 159.315 ;
        RECT 58.645 159.145 58.815 159.315 ;
        RECT 59.105 159.145 59.275 159.315 ;
        RECT 59.565 159.145 59.735 159.315 ;
        RECT 60.025 159.145 60.195 159.315 ;
        RECT 60.485 159.145 60.655 159.315 ;
        RECT 60.945 159.145 61.115 159.315 ;
        RECT 61.405 159.145 61.575 159.315 ;
        RECT 61.865 159.145 62.035 159.315 ;
        RECT 62.325 159.145 62.495 159.315 ;
        RECT 62.785 159.145 62.955 159.315 ;
        RECT 63.245 159.145 63.415 159.315 ;
        RECT 63.705 159.145 63.875 159.315 ;
        RECT 64.165 159.145 64.335 159.315 ;
        RECT 64.625 159.145 64.795 159.315 ;
        RECT 65.085 159.145 65.255 159.315 ;
        RECT 65.545 159.145 65.715 159.315 ;
        RECT 66.005 159.145 66.175 159.315 ;
        RECT 66.465 159.145 66.635 159.315 ;
        RECT 66.925 159.145 67.095 159.315 ;
        RECT 67.385 159.145 67.555 159.315 ;
        RECT 67.845 159.145 68.015 159.315 ;
        RECT 68.305 159.145 68.475 159.315 ;
        RECT 68.765 159.145 68.935 159.315 ;
        RECT 69.225 159.145 69.395 159.315 ;
        RECT 69.685 159.145 69.855 159.315 ;
        RECT 70.145 159.145 70.315 159.315 ;
        RECT 70.605 159.145 70.775 159.315 ;
        RECT 71.065 159.145 71.235 159.315 ;
        RECT 71.525 159.145 71.695 159.315 ;
        RECT 71.985 159.145 72.155 159.315 ;
        RECT 72.445 159.145 72.615 159.315 ;
        RECT 72.905 159.145 73.075 159.315 ;
        RECT 73.365 159.145 73.535 159.315 ;
        RECT 73.825 159.145 73.995 159.315 ;
        RECT 74.285 159.145 74.455 159.315 ;
        RECT 74.745 159.145 74.915 159.315 ;
        RECT 75.205 159.145 75.375 159.315 ;
        RECT 75.665 159.145 75.835 159.315 ;
        RECT 76.125 159.145 76.295 159.315 ;
        RECT 76.585 159.145 76.755 159.315 ;
        RECT 77.045 159.145 77.215 159.315 ;
        RECT 77.505 159.145 77.675 159.315 ;
        RECT 77.965 159.145 78.135 159.315 ;
        RECT 78.425 159.145 78.595 159.315 ;
        RECT 78.885 159.145 79.055 159.315 ;
        RECT 79.345 159.145 79.515 159.315 ;
        RECT 79.805 159.145 79.975 159.315 ;
        RECT 80.265 159.145 80.435 159.315 ;
        RECT 80.725 159.145 80.895 159.315 ;
        RECT 81.185 159.145 81.355 159.315 ;
        RECT 81.645 159.145 81.815 159.315 ;
        RECT 82.105 159.145 82.275 159.315 ;
        RECT 82.565 159.145 82.735 159.315 ;
        RECT 83.025 159.145 83.195 159.315 ;
        RECT 83.485 159.145 83.655 159.315 ;
        RECT 83.945 159.145 84.115 159.315 ;
        RECT 84.405 159.145 84.575 159.315 ;
        RECT 84.865 159.145 85.035 159.315 ;
        RECT 85.325 159.145 85.495 159.315 ;
        RECT 85.785 159.145 85.955 159.315 ;
        RECT 86.245 159.145 86.415 159.315 ;
        RECT 86.705 159.145 86.875 159.315 ;
        RECT 87.165 159.145 87.335 159.315 ;
        RECT 87.625 159.145 87.795 159.315 ;
        RECT 88.085 159.145 88.255 159.315 ;
        RECT 88.545 159.145 88.715 159.315 ;
        RECT 89.005 159.145 89.175 159.315 ;
        RECT 89.465 159.145 89.635 159.315 ;
        RECT 89.925 159.145 90.095 159.315 ;
        RECT 90.385 159.145 90.555 159.315 ;
        RECT 90.845 159.145 91.015 159.315 ;
        RECT 91.305 159.145 91.475 159.315 ;
        RECT 91.765 159.145 91.935 159.315 ;
        RECT 92.225 159.145 92.395 159.315 ;
        RECT 92.685 159.145 92.855 159.315 ;
        RECT 93.145 159.145 93.315 159.315 ;
        RECT 93.605 159.145 93.775 159.315 ;
        RECT 94.065 159.145 94.235 159.315 ;
        RECT 94.525 159.145 94.695 159.315 ;
        RECT 94.985 159.145 95.155 159.315 ;
        RECT 95.445 159.145 95.615 159.315 ;
        RECT 95.905 159.145 96.075 159.315 ;
        RECT 96.365 159.145 96.535 159.315 ;
        RECT 96.825 159.145 96.995 159.315 ;
        RECT 97.285 159.145 97.455 159.315 ;
        RECT 97.745 159.145 97.915 159.315 ;
        RECT 98.205 159.145 98.375 159.315 ;
        RECT 98.665 159.145 98.835 159.315 ;
        RECT 99.125 159.145 99.295 159.315 ;
        RECT 99.585 159.145 99.755 159.315 ;
        RECT 100.045 159.145 100.215 159.315 ;
        RECT 100.505 159.145 100.675 159.315 ;
        RECT 100.965 159.145 101.135 159.315 ;
        RECT 101.425 159.145 101.595 159.315 ;
        RECT 101.885 159.145 102.055 159.315 ;
        RECT 102.345 159.145 102.515 159.315 ;
        RECT 102.805 159.145 102.975 159.315 ;
        RECT 103.265 159.145 103.435 159.315 ;
        RECT 103.725 159.145 103.895 159.315 ;
        RECT 104.185 159.145 104.355 159.315 ;
        RECT 104.645 159.145 104.815 159.315 ;
        RECT 105.105 159.145 105.275 159.315 ;
        RECT 105.565 159.145 105.735 159.315 ;
        RECT 106.025 159.145 106.195 159.315 ;
        RECT 106.485 159.145 106.655 159.315 ;
        RECT 106.945 159.145 107.115 159.315 ;
        RECT 107.405 159.145 107.575 159.315 ;
        RECT 107.865 159.145 108.035 159.315 ;
        RECT 108.325 159.145 108.495 159.315 ;
        RECT 108.785 159.145 108.955 159.315 ;
        RECT 109.245 159.145 109.415 159.315 ;
        RECT 109.705 159.145 109.875 159.315 ;
        RECT 110.165 159.145 110.335 159.315 ;
        RECT 110.625 159.145 110.795 159.315 ;
        RECT 111.085 159.145 111.255 159.315 ;
        RECT 111.545 159.145 111.715 159.315 ;
        RECT 112.005 159.145 112.175 159.315 ;
        RECT 112.465 159.145 112.635 159.315 ;
        RECT 112.925 159.145 113.095 159.315 ;
        RECT 113.385 159.145 113.555 159.315 ;
        RECT 113.845 159.145 114.015 159.315 ;
        RECT 114.305 159.145 114.475 159.315 ;
        RECT 114.765 159.145 114.935 159.315 ;
        RECT 115.225 159.145 115.395 159.315 ;
        RECT 115.685 159.145 115.855 159.315 ;
        RECT 116.145 159.145 116.315 159.315 ;
        RECT 116.605 159.145 116.775 159.315 ;
        RECT 117.065 159.145 117.235 159.315 ;
        RECT 117.525 159.145 117.695 159.315 ;
        RECT 117.985 159.145 118.155 159.315 ;
        RECT 118.445 159.145 118.615 159.315 ;
        RECT 118.905 159.145 119.075 159.315 ;
        RECT 119.365 159.145 119.535 159.315 ;
        RECT 119.825 159.145 119.995 159.315 ;
        RECT 120.285 159.145 120.455 159.315 ;
        RECT 120.745 159.145 120.915 159.315 ;
        RECT 121.205 159.145 121.375 159.315 ;
        RECT 121.665 159.145 121.835 159.315 ;
        RECT 122.125 159.145 122.295 159.315 ;
        RECT 122.585 159.145 122.755 159.315 ;
        RECT 123.045 159.145 123.215 159.315 ;
        RECT 123.505 159.145 123.675 159.315 ;
        RECT 123.965 159.145 124.135 159.315 ;
        RECT 124.425 159.145 124.595 159.315 ;
        RECT 124.885 159.145 125.055 159.315 ;
        RECT 125.345 159.145 125.515 159.315 ;
        RECT 125.805 159.145 125.975 159.315 ;
        RECT 126.265 159.145 126.435 159.315 ;
        RECT 126.725 159.145 126.895 159.315 ;
        RECT 127.185 159.145 127.355 159.315 ;
        RECT 127.645 159.145 127.815 159.315 ;
        RECT 128.105 159.145 128.275 159.315 ;
        RECT 128.565 159.145 128.735 159.315 ;
        RECT 129.025 159.145 129.195 159.315 ;
        RECT 129.485 159.145 129.655 159.315 ;
        RECT 129.945 159.145 130.115 159.315 ;
        RECT 130.405 159.145 130.575 159.315 ;
        RECT 130.865 159.145 131.035 159.315 ;
        RECT 131.325 159.145 131.495 159.315 ;
        RECT 131.785 159.145 131.955 159.315 ;
        RECT 132.245 159.145 132.415 159.315 ;
        RECT 132.705 159.145 132.875 159.315 ;
        RECT 133.165 159.145 133.335 159.315 ;
        RECT 133.625 159.145 133.795 159.315 ;
        RECT 134.085 159.145 134.255 159.315 ;
        RECT 134.545 159.145 134.715 159.315 ;
        RECT 135.005 159.145 135.175 159.315 ;
        RECT 135.465 159.145 135.635 159.315 ;
        RECT 135.925 159.145 136.095 159.315 ;
        RECT 136.385 159.145 136.555 159.315 ;
        RECT 136.845 159.145 137.015 159.315 ;
        RECT 137.305 159.145 137.475 159.315 ;
        RECT 137.765 159.145 137.935 159.315 ;
        RECT 138.225 159.145 138.395 159.315 ;
        RECT 138.685 159.145 138.855 159.315 ;
        RECT 139.145 159.145 139.315 159.315 ;
        RECT 139.605 159.145 139.775 159.315 ;
        RECT 140.065 159.145 140.235 159.315 ;
        RECT 140.525 159.145 140.695 159.315 ;
        RECT 140.985 159.145 141.155 159.315 ;
        RECT 141.445 159.145 141.615 159.315 ;
        RECT 141.905 159.145 142.075 159.315 ;
        RECT 142.365 159.145 142.535 159.315 ;
        RECT 142.825 159.145 142.995 159.315 ;
        RECT 143.285 159.145 143.455 159.315 ;
        RECT 143.745 159.145 143.915 159.315 ;
        RECT 144.205 159.145 144.375 159.315 ;
        RECT 144.665 159.145 144.835 159.315 ;
        RECT 145.125 159.145 145.295 159.315 ;
        RECT 145.585 159.145 145.755 159.315 ;
        RECT 146.045 159.145 146.215 159.315 ;
        RECT 146.505 159.145 146.675 159.315 ;
        RECT 146.965 159.145 147.135 159.315 ;
        RECT 147.425 159.145 147.595 159.315 ;
        RECT 147.885 159.145 148.055 159.315 ;
        RECT 148.345 159.145 148.515 159.315 ;
        RECT 148.805 159.145 148.975 159.315 ;
        RECT 149.265 159.145 149.435 159.315 ;
        RECT 149.725 159.145 149.895 159.315 ;
        RECT 150.185 159.145 150.355 159.315 ;
        RECT 25.065 157.615 25.235 157.785 ;
        RECT 25.525 157.615 25.695 157.785 ;
        RECT 26.445 157.615 26.615 157.785 ;
        RECT 26.905 158.635 27.075 158.805 ;
        RECT 27.825 157.615 27.995 157.785 ;
        RECT 53.125 158.635 53.295 158.805 ;
        RECT 50.365 157.275 50.535 157.445 ;
        RECT 51.285 156.935 51.455 157.105 ;
        RECT 51.745 156.935 51.915 157.105 ;
        RECT 52.205 156.935 52.375 157.105 ;
        RECT 57.725 158.635 57.895 158.805 ;
        RECT 58.645 158.635 58.815 158.805 ;
        RECT 56.805 157.275 56.975 157.445 ;
        RECT 57.805 156.935 57.975 157.105 ;
        RECT 71.065 158.635 71.235 158.805 ;
        RECT 74.285 158.635 74.455 158.805 ;
        RECT 75.205 158.635 75.375 158.805 ;
        RECT 72.905 157.955 73.075 158.125 ;
        RECT 71.985 157.615 72.155 157.785 ;
        RECT 73.365 157.275 73.535 157.445 ;
        RECT 74.415 156.935 74.585 157.105 ;
        RECT 78.885 157.955 79.055 158.125 ;
        RECT 78.425 157.615 78.595 157.785 ;
        RECT 80.265 157.955 80.435 158.125 ;
        RECT 84.865 157.955 85.035 158.125 ;
        RECT 89.005 158.635 89.175 158.805 ;
        RECT 84.405 157.615 84.575 157.785 ;
        RECT 85.325 157.615 85.495 157.785 ;
        RECT 85.785 157.615 85.955 157.785 ;
        RECT 86.250 157.615 86.420 157.785 ;
        RECT 87.165 157.615 87.335 157.785 ;
        RECT 88.110 157.615 88.280 157.785 ;
        RECT 87.625 157.275 87.795 157.445 ;
        RECT 91.305 157.955 91.475 158.125 ;
        RECT 90.385 157.275 90.555 157.445 ;
        RECT 93.605 158.635 93.775 158.805 ;
        RECT 94.985 157.615 95.155 157.785 ;
        RECT 95.445 157.615 95.615 157.785 ;
        RECT 95.905 157.615 96.075 157.785 ;
        RECT 97.285 157.955 97.455 158.125 ;
        RECT 96.825 157.615 96.995 157.785 ;
        RECT 98.205 157.615 98.375 157.785 ;
        RECT 98.665 157.615 98.835 157.785 ;
        RECT 99.125 157.955 99.295 158.125 ;
        RECT 99.585 157.955 99.755 158.125 ;
        RECT 103.265 157.955 103.435 158.125 ;
        RECT 103.725 157.615 103.895 157.785 ;
        RECT 101.885 156.935 102.055 157.105 ;
        RECT 110.165 157.615 110.335 157.785 ;
        RECT 110.625 156.935 110.795 157.105 ;
        RECT 11.265 156.425 11.435 156.595 ;
        RECT 11.725 156.425 11.895 156.595 ;
        RECT 12.185 156.425 12.355 156.595 ;
        RECT 12.645 156.425 12.815 156.595 ;
        RECT 13.105 156.425 13.275 156.595 ;
        RECT 13.565 156.425 13.735 156.595 ;
        RECT 14.025 156.425 14.195 156.595 ;
        RECT 14.485 156.425 14.655 156.595 ;
        RECT 14.945 156.425 15.115 156.595 ;
        RECT 15.405 156.425 15.575 156.595 ;
        RECT 15.865 156.425 16.035 156.595 ;
        RECT 16.325 156.425 16.495 156.595 ;
        RECT 16.785 156.425 16.955 156.595 ;
        RECT 17.245 156.425 17.415 156.595 ;
        RECT 17.705 156.425 17.875 156.595 ;
        RECT 18.165 156.425 18.335 156.595 ;
        RECT 18.625 156.425 18.795 156.595 ;
        RECT 19.085 156.425 19.255 156.595 ;
        RECT 19.545 156.425 19.715 156.595 ;
        RECT 20.005 156.425 20.175 156.595 ;
        RECT 20.465 156.425 20.635 156.595 ;
        RECT 20.925 156.425 21.095 156.595 ;
        RECT 21.385 156.425 21.555 156.595 ;
        RECT 21.845 156.425 22.015 156.595 ;
        RECT 22.305 156.425 22.475 156.595 ;
        RECT 22.765 156.425 22.935 156.595 ;
        RECT 23.225 156.425 23.395 156.595 ;
        RECT 23.685 156.425 23.855 156.595 ;
        RECT 24.145 156.425 24.315 156.595 ;
        RECT 24.605 156.425 24.775 156.595 ;
        RECT 25.065 156.425 25.235 156.595 ;
        RECT 25.525 156.425 25.695 156.595 ;
        RECT 25.985 156.425 26.155 156.595 ;
        RECT 26.445 156.425 26.615 156.595 ;
        RECT 26.905 156.425 27.075 156.595 ;
        RECT 27.365 156.425 27.535 156.595 ;
        RECT 27.825 156.425 27.995 156.595 ;
        RECT 28.285 156.425 28.455 156.595 ;
        RECT 28.745 156.425 28.915 156.595 ;
        RECT 29.205 156.425 29.375 156.595 ;
        RECT 29.665 156.425 29.835 156.595 ;
        RECT 30.125 156.425 30.295 156.595 ;
        RECT 30.585 156.425 30.755 156.595 ;
        RECT 31.045 156.425 31.215 156.595 ;
        RECT 31.505 156.425 31.675 156.595 ;
        RECT 31.965 156.425 32.135 156.595 ;
        RECT 32.425 156.425 32.595 156.595 ;
        RECT 32.885 156.425 33.055 156.595 ;
        RECT 33.345 156.425 33.515 156.595 ;
        RECT 33.805 156.425 33.975 156.595 ;
        RECT 34.265 156.425 34.435 156.595 ;
        RECT 34.725 156.425 34.895 156.595 ;
        RECT 35.185 156.425 35.355 156.595 ;
        RECT 35.645 156.425 35.815 156.595 ;
        RECT 36.105 156.425 36.275 156.595 ;
        RECT 36.565 156.425 36.735 156.595 ;
        RECT 37.025 156.425 37.195 156.595 ;
        RECT 37.485 156.425 37.655 156.595 ;
        RECT 37.945 156.425 38.115 156.595 ;
        RECT 38.405 156.425 38.575 156.595 ;
        RECT 38.865 156.425 39.035 156.595 ;
        RECT 39.325 156.425 39.495 156.595 ;
        RECT 39.785 156.425 39.955 156.595 ;
        RECT 40.245 156.425 40.415 156.595 ;
        RECT 40.705 156.425 40.875 156.595 ;
        RECT 41.165 156.425 41.335 156.595 ;
        RECT 41.625 156.425 41.795 156.595 ;
        RECT 42.085 156.425 42.255 156.595 ;
        RECT 42.545 156.425 42.715 156.595 ;
        RECT 43.005 156.425 43.175 156.595 ;
        RECT 43.465 156.425 43.635 156.595 ;
        RECT 43.925 156.425 44.095 156.595 ;
        RECT 44.385 156.425 44.555 156.595 ;
        RECT 44.845 156.425 45.015 156.595 ;
        RECT 45.305 156.425 45.475 156.595 ;
        RECT 45.765 156.425 45.935 156.595 ;
        RECT 46.225 156.425 46.395 156.595 ;
        RECT 46.685 156.425 46.855 156.595 ;
        RECT 47.145 156.425 47.315 156.595 ;
        RECT 47.605 156.425 47.775 156.595 ;
        RECT 48.065 156.425 48.235 156.595 ;
        RECT 48.525 156.425 48.695 156.595 ;
        RECT 48.985 156.425 49.155 156.595 ;
        RECT 49.445 156.425 49.615 156.595 ;
        RECT 49.905 156.425 50.075 156.595 ;
        RECT 50.365 156.425 50.535 156.595 ;
        RECT 50.825 156.425 50.995 156.595 ;
        RECT 51.285 156.425 51.455 156.595 ;
        RECT 51.745 156.425 51.915 156.595 ;
        RECT 52.205 156.425 52.375 156.595 ;
        RECT 52.665 156.425 52.835 156.595 ;
        RECT 53.125 156.425 53.295 156.595 ;
        RECT 53.585 156.425 53.755 156.595 ;
        RECT 54.045 156.425 54.215 156.595 ;
        RECT 54.505 156.425 54.675 156.595 ;
        RECT 54.965 156.425 55.135 156.595 ;
        RECT 55.425 156.425 55.595 156.595 ;
        RECT 55.885 156.425 56.055 156.595 ;
        RECT 56.345 156.425 56.515 156.595 ;
        RECT 56.805 156.425 56.975 156.595 ;
        RECT 57.265 156.425 57.435 156.595 ;
        RECT 57.725 156.425 57.895 156.595 ;
        RECT 58.185 156.425 58.355 156.595 ;
        RECT 58.645 156.425 58.815 156.595 ;
        RECT 59.105 156.425 59.275 156.595 ;
        RECT 59.565 156.425 59.735 156.595 ;
        RECT 60.025 156.425 60.195 156.595 ;
        RECT 60.485 156.425 60.655 156.595 ;
        RECT 60.945 156.425 61.115 156.595 ;
        RECT 61.405 156.425 61.575 156.595 ;
        RECT 61.865 156.425 62.035 156.595 ;
        RECT 62.325 156.425 62.495 156.595 ;
        RECT 62.785 156.425 62.955 156.595 ;
        RECT 63.245 156.425 63.415 156.595 ;
        RECT 63.705 156.425 63.875 156.595 ;
        RECT 64.165 156.425 64.335 156.595 ;
        RECT 64.625 156.425 64.795 156.595 ;
        RECT 65.085 156.425 65.255 156.595 ;
        RECT 65.545 156.425 65.715 156.595 ;
        RECT 66.005 156.425 66.175 156.595 ;
        RECT 66.465 156.425 66.635 156.595 ;
        RECT 66.925 156.425 67.095 156.595 ;
        RECT 67.385 156.425 67.555 156.595 ;
        RECT 67.845 156.425 68.015 156.595 ;
        RECT 68.305 156.425 68.475 156.595 ;
        RECT 68.765 156.425 68.935 156.595 ;
        RECT 69.225 156.425 69.395 156.595 ;
        RECT 69.685 156.425 69.855 156.595 ;
        RECT 70.145 156.425 70.315 156.595 ;
        RECT 70.605 156.425 70.775 156.595 ;
        RECT 71.065 156.425 71.235 156.595 ;
        RECT 71.525 156.425 71.695 156.595 ;
        RECT 71.985 156.425 72.155 156.595 ;
        RECT 72.445 156.425 72.615 156.595 ;
        RECT 72.905 156.425 73.075 156.595 ;
        RECT 73.365 156.425 73.535 156.595 ;
        RECT 73.825 156.425 73.995 156.595 ;
        RECT 74.285 156.425 74.455 156.595 ;
        RECT 74.745 156.425 74.915 156.595 ;
        RECT 75.205 156.425 75.375 156.595 ;
        RECT 75.665 156.425 75.835 156.595 ;
        RECT 76.125 156.425 76.295 156.595 ;
        RECT 76.585 156.425 76.755 156.595 ;
        RECT 77.045 156.425 77.215 156.595 ;
        RECT 77.505 156.425 77.675 156.595 ;
        RECT 77.965 156.425 78.135 156.595 ;
        RECT 78.425 156.425 78.595 156.595 ;
        RECT 78.885 156.425 79.055 156.595 ;
        RECT 79.345 156.425 79.515 156.595 ;
        RECT 79.805 156.425 79.975 156.595 ;
        RECT 80.265 156.425 80.435 156.595 ;
        RECT 80.725 156.425 80.895 156.595 ;
        RECT 81.185 156.425 81.355 156.595 ;
        RECT 81.645 156.425 81.815 156.595 ;
        RECT 82.105 156.425 82.275 156.595 ;
        RECT 82.565 156.425 82.735 156.595 ;
        RECT 83.025 156.425 83.195 156.595 ;
        RECT 83.485 156.425 83.655 156.595 ;
        RECT 83.945 156.425 84.115 156.595 ;
        RECT 84.405 156.425 84.575 156.595 ;
        RECT 84.865 156.425 85.035 156.595 ;
        RECT 85.325 156.425 85.495 156.595 ;
        RECT 85.785 156.425 85.955 156.595 ;
        RECT 86.245 156.425 86.415 156.595 ;
        RECT 86.705 156.425 86.875 156.595 ;
        RECT 87.165 156.425 87.335 156.595 ;
        RECT 87.625 156.425 87.795 156.595 ;
        RECT 88.085 156.425 88.255 156.595 ;
        RECT 88.545 156.425 88.715 156.595 ;
        RECT 89.005 156.425 89.175 156.595 ;
        RECT 89.465 156.425 89.635 156.595 ;
        RECT 89.925 156.425 90.095 156.595 ;
        RECT 90.385 156.425 90.555 156.595 ;
        RECT 90.845 156.425 91.015 156.595 ;
        RECT 91.305 156.425 91.475 156.595 ;
        RECT 91.765 156.425 91.935 156.595 ;
        RECT 92.225 156.425 92.395 156.595 ;
        RECT 92.685 156.425 92.855 156.595 ;
        RECT 93.145 156.425 93.315 156.595 ;
        RECT 93.605 156.425 93.775 156.595 ;
        RECT 94.065 156.425 94.235 156.595 ;
        RECT 94.525 156.425 94.695 156.595 ;
        RECT 94.985 156.425 95.155 156.595 ;
        RECT 95.445 156.425 95.615 156.595 ;
        RECT 95.905 156.425 96.075 156.595 ;
        RECT 96.365 156.425 96.535 156.595 ;
        RECT 96.825 156.425 96.995 156.595 ;
        RECT 97.285 156.425 97.455 156.595 ;
        RECT 97.745 156.425 97.915 156.595 ;
        RECT 98.205 156.425 98.375 156.595 ;
        RECT 98.665 156.425 98.835 156.595 ;
        RECT 99.125 156.425 99.295 156.595 ;
        RECT 99.585 156.425 99.755 156.595 ;
        RECT 100.045 156.425 100.215 156.595 ;
        RECT 100.505 156.425 100.675 156.595 ;
        RECT 100.965 156.425 101.135 156.595 ;
        RECT 101.425 156.425 101.595 156.595 ;
        RECT 101.885 156.425 102.055 156.595 ;
        RECT 102.345 156.425 102.515 156.595 ;
        RECT 102.805 156.425 102.975 156.595 ;
        RECT 103.265 156.425 103.435 156.595 ;
        RECT 103.725 156.425 103.895 156.595 ;
        RECT 104.185 156.425 104.355 156.595 ;
        RECT 104.645 156.425 104.815 156.595 ;
        RECT 105.105 156.425 105.275 156.595 ;
        RECT 105.565 156.425 105.735 156.595 ;
        RECT 106.025 156.425 106.195 156.595 ;
        RECT 106.485 156.425 106.655 156.595 ;
        RECT 106.945 156.425 107.115 156.595 ;
        RECT 107.405 156.425 107.575 156.595 ;
        RECT 107.865 156.425 108.035 156.595 ;
        RECT 108.325 156.425 108.495 156.595 ;
        RECT 108.785 156.425 108.955 156.595 ;
        RECT 109.245 156.425 109.415 156.595 ;
        RECT 109.705 156.425 109.875 156.595 ;
        RECT 110.165 156.425 110.335 156.595 ;
        RECT 110.625 156.425 110.795 156.595 ;
        RECT 111.085 156.425 111.255 156.595 ;
        RECT 111.545 156.425 111.715 156.595 ;
        RECT 112.005 156.425 112.175 156.595 ;
        RECT 112.465 156.425 112.635 156.595 ;
        RECT 112.925 156.425 113.095 156.595 ;
        RECT 113.385 156.425 113.555 156.595 ;
        RECT 113.845 156.425 114.015 156.595 ;
        RECT 114.305 156.425 114.475 156.595 ;
        RECT 114.765 156.425 114.935 156.595 ;
        RECT 115.225 156.425 115.395 156.595 ;
        RECT 115.685 156.425 115.855 156.595 ;
        RECT 116.145 156.425 116.315 156.595 ;
        RECT 116.605 156.425 116.775 156.595 ;
        RECT 117.065 156.425 117.235 156.595 ;
        RECT 117.525 156.425 117.695 156.595 ;
        RECT 117.985 156.425 118.155 156.595 ;
        RECT 118.445 156.425 118.615 156.595 ;
        RECT 118.905 156.425 119.075 156.595 ;
        RECT 119.365 156.425 119.535 156.595 ;
        RECT 119.825 156.425 119.995 156.595 ;
        RECT 120.285 156.425 120.455 156.595 ;
        RECT 120.745 156.425 120.915 156.595 ;
        RECT 121.205 156.425 121.375 156.595 ;
        RECT 121.665 156.425 121.835 156.595 ;
        RECT 122.125 156.425 122.295 156.595 ;
        RECT 122.585 156.425 122.755 156.595 ;
        RECT 123.045 156.425 123.215 156.595 ;
        RECT 123.505 156.425 123.675 156.595 ;
        RECT 123.965 156.425 124.135 156.595 ;
        RECT 124.425 156.425 124.595 156.595 ;
        RECT 124.885 156.425 125.055 156.595 ;
        RECT 125.345 156.425 125.515 156.595 ;
        RECT 125.805 156.425 125.975 156.595 ;
        RECT 126.265 156.425 126.435 156.595 ;
        RECT 126.725 156.425 126.895 156.595 ;
        RECT 127.185 156.425 127.355 156.595 ;
        RECT 127.645 156.425 127.815 156.595 ;
        RECT 128.105 156.425 128.275 156.595 ;
        RECT 128.565 156.425 128.735 156.595 ;
        RECT 129.025 156.425 129.195 156.595 ;
        RECT 129.485 156.425 129.655 156.595 ;
        RECT 129.945 156.425 130.115 156.595 ;
        RECT 130.405 156.425 130.575 156.595 ;
        RECT 130.865 156.425 131.035 156.595 ;
        RECT 131.325 156.425 131.495 156.595 ;
        RECT 131.785 156.425 131.955 156.595 ;
        RECT 132.245 156.425 132.415 156.595 ;
        RECT 132.705 156.425 132.875 156.595 ;
        RECT 133.165 156.425 133.335 156.595 ;
        RECT 133.625 156.425 133.795 156.595 ;
        RECT 134.085 156.425 134.255 156.595 ;
        RECT 134.545 156.425 134.715 156.595 ;
        RECT 135.005 156.425 135.175 156.595 ;
        RECT 135.465 156.425 135.635 156.595 ;
        RECT 135.925 156.425 136.095 156.595 ;
        RECT 136.385 156.425 136.555 156.595 ;
        RECT 136.845 156.425 137.015 156.595 ;
        RECT 137.305 156.425 137.475 156.595 ;
        RECT 137.765 156.425 137.935 156.595 ;
        RECT 138.225 156.425 138.395 156.595 ;
        RECT 138.685 156.425 138.855 156.595 ;
        RECT 139.145 156.425 139.315 156.595 ;
        RECT 139.605 156.425 139.775 156.595 ;
        RECT 140.065 156.425 140.235 156.595 ;
        RECT 140.525 156.425 140.695 156.595 ;
        RECT 140.985 156.425 141.155 156.595 ;
        RECT 141.445 156.425 141.615 156.595 ;
        RECT 141.905 156.425 142.075 156.595 ;
        RECT 142.365 156.425 142.535 156.595 ;
        RECT 142.825 156.425 142.995 156.595 ;
        RECT 143.285 156.425 143.455 156.595 ;
        RECT 143.745 156.425 143.915 156.595 ;
        RECT 144.205 156.425 144.375 156.595 ;
        RECT 144.665 156.425 144.835 156.595 ;
        RECT 145.125 156.425 145.295 156.595 ;
        RECT 145.585 156.425 145.755 156.595 ;
        RECT 146.045 156.425 146.215 156.595 ;
        RECT 146.505 156.425 146.675 156.595 ;
        RECT 146.965 156.425 147.135 156.595 ;
        RECT 147.425 156.425 147.595 156.595 ;
        RECT 147.885 156.425 148.055 156.595 ;
        RECT 148.345 156.425 148.515 156.595 ;
        RECT 148.805 156.425 148.975 156.595 ;
        RECT 149.265 156.425 149.435 156.595 ;
        RECT 149.725 156.425 149.895 156.595 ;
        RECT 150.185 156.425 150.355 156.595 ;
        RECT 19.085 155.235 19.255 155.405 ;
        RECT 29.205 155.915 29.375 156.085 ;
        RECT 18.165 154.215 18.335 154.385 ;
        RECT 30.585 155.575 30.755 155.745 ;
        RECT 30.125 155.235 30.295 155.405 ;
        RECT 31.045 155.235 31.215 155.405 ;
        RECT 31.965 155.235 32.135 155.405 ;
        RECT 34.725 155.235 34.895 155.405 ;
        RECT 35.185 154.895 35.355 155.065 ;
        RECT 36.565 154.555 36.735 154.725 ;
        RECT 39.785 155.575 39.955 155.745 ;
        RECT 38.865 155.235 39.035 155.405 ;
        RECT 40.245 155.575 40.415 155.745 ;
        RECT 40.805 155.345 40.975 155.515 ;
        RECT 41.625 155.235 41.795 155.405 ;
        RECT 42.085 155.235 42.255 155.405 ;
        RECT 43.005 155.235 43.175 155.405 ;
        RECT 38.865 154.555 39.035 154.725 ;
        RECT 43.925 155.235 44.095 155.405 ;
        RECT 44.385 155.235 44.555 155.405 ;
        RECT 48.065 155.915 48.235 156.085 ;
        RECT 45.305 155.235 45.475 155.405 ;
        RECT 47.145 155.235 47.315 155.405 ;
        RECT 45.765 154.895 45.935 155.065 ;
        RECT 48.525 154.895 48.695 155.065 ;
        RECT 50.365 155.235 50.535 155.405 ;
        RECT 53.125 155.235 53.295 155.405 ;
        RECT 53.585 155.235 53.755 155.405 ;
        RECT 57.265 155.915 57.435 156.085 ;
        RECT 56.345 155.235 56.515 155.405 ;
        RECT 57.265 155.235 57.435 155.405 ;
        RECT 53.125 154.215 53.295 154.385 ;
        RECT 54.045 154.215 54.215 154.385 ;
        RECT 59.105 155.235 59.275 155.405 ;
        RECT 64.165 155.235 64.335 155.405 ;
        RECT 60.025 154.215 60.195 154.385 ;
        RECT 64.650 154.555 64.820 154.725 ;
        RECT 65.045 154.895 65.215 155.065 ;
        RECT 65.500 155.575 65.670 155.745 ;
        RECT 66.235 154.895 66.405 155.065 ;
        RECT 66.750 154.555 66.920 154.725 ;
        RECT 68.320 154.555 68.490 154.725 ;
        RECT 68.755 154.895 68.925 155.065 ;
        RECT 71.065 155.915 71.235 156.085 ;
        RECT 72.905 154.555 73.075 154.725 ;
        RECT 73.825 154.895 73.995 155.065 ;
        RECT 73.365 154.215 73.535 154.385 ;
        RECT 83.485 155.575 83.655 155.745 ;
        RECT 85.325 155.915 85.495 156.085 ;
        RECT 84.565 155.575 84.735 155.745 ;
        RECT 87.165 155.235 87.335 155.405 ;
        RECT 88.085 155.235 88.255 155.405 ;
        RECT 84.405 154.215 84.575 154.385 ;
        RECT 88.085 154.215 88.255 154.385 ;
        RECT 92.685 155.235 92.855 155.405 ;
        RECT 95.905 155.915 96.075 156.085 ;
        RECT 94.065 154.895 94.235 155.065 ;
        RECT 95.110 155.235 95.280 155.405 ;
        RECT 96.365 155.915 96.535 156.085 ;
        RECT 97.285 155.575 97.455 155.745 ;
        RECT 97.285 154.215 97.455 154.385 ;
        RECT 99.125 155.235 99.295 155.405 ;
        RECT 101.345 155.575 101.515 155.745 ;
        RECT 102.345 155.575 102.515 155.745 ;
        RECT 100.505 154.215 100.675 154.385 ;
        RECT 101.425 154.215 101.595 154.385 ;
        RECT 108.325 155.235 108.495 155.405 ;
        RECT 109.245 155.235 109.415 155.405 ;
        RECT 108.785 154.215 108.955 154.385 ;
        RECT 11.265 153.705 11.435 153.875 ;
        RECT 11.725 153.705 11.895 153.875 ;
        RECT 12.185 153.705 12.355 153.875 ;
        RECT 12.645 153.705 12.815 153.875 ;
        RECT 13.105 153.705 13.275 153.875 ;
        RECT 13.565 153.705 13.735 153.875 ;
        RECT 14.025 153.705 14.195 153.875 ;
        RECT 14.485 153.705 14.655 153.875 ;
        RECT 14.945 153.705 15.115 153.875 ;
        RECT 15.405 153.705 15.575 153.875 ;
        RECT 15.865 153.705 16.035 153.875 ;
        RECT 16.325 153.705 16.495 153.875 ;
        RECT 16.785 153.705 16.955 153.875 ;
        RECT 17.245 153.705 17.415 153.875 ;
        RECT 17.705 153.705 17.875 153.875 ;
        RECT 18.165 153.705 18.335 153.875 ;
        RECT 18.625 153.705 18.795 153.875 ;
        RECT 19.085 153.705 19.255 153.875 ;
        RECT 19.545 153.705 19.715 153.875 ;
        RECT 20.005 153.705 20.175 153.875 ;
        RECT 20.465 153.705 20.635 153.875 ;
        RECT 20.925 153.705 21.095 153.875 ;
        RECT 21.385 153.705 21.555 153.875 ;
        RECT 21.845 153.705 22.015 153.875 ;
        RECT 22.305 153.705 22.475 153.875 ;
        RECT 22.765 153.705 22.935 153.875 ;
        RECT 23.225 153.705 23.395 153.875 ;
        RECT 23.685 153.705 23.855 153.875 ;
        RECT 24.145 153.705 24.315 153.875 ;
        RECT 24.605 153.705 24.775 153.875 ;
        RECT 25.065 153.705 25.235 153.875 ;
        RECT 25.525 153.705 25.695 153.875 ;
        RECT 25.985 153.705 26.155 153.875 ;
        RECT 26.445 153.705 26.615 153.875 ;
        RECT 26.905 153.705 27.075 153.875 ;
        RECT 27.365 153.705 27.535 153.875 ;
        RECT 27.825 153.705 27.995 153.875 ;
        RECT 28.285 153.705 28.455 153.875 ;
        RECT 28.745 153.705 28.915 153.875 ;
        RECT 29.205 153.705 29.375 153.875 ;
        RECT 29.665 153.705 29.835 153.875 ;
        RECT 30.125 153.705 30.295 153.875 ;
        RECT 30.585 153.705 30.755 153.875 ;
        RECT 31.045 153.705 31.215 153.875 ;
        RECT 31.505 153.705 31.675 153.875 ;
        RECT 31.965 153.705 32.135 153.875 ;
        RECT 32.425 153.705 32.595 153.875 ;
        RECT 32.885 153.705 33.055 153.875 ;
        RECT 33.345 153.705 33.515 153.875 ;
        RECT 33.805 153.705 33.975 153.875 ;
        RECT 34.265 153.705 34.435 153.875 ;
        RECT 34.725 153.705 34.895 153.875 ;
        RECT 35.185 153.705 35.355 153.875 ;
        RECT 35.645 153.705 35.815 153.875 ;
        RECT 36.105 153.705 36.275 153.875 ;
        RECT 36.565 153.705 36.735 153.875 ;
        RECT 37.025 153.705 37.195 153.875 ;
        RECT 37.485 153.705 37.655 153.875 ;
        RECT 37.945 153.705 38.115 153.875 ;
        RECT 38.405 153.705 38.575 153.875 ;
        RECT 38.865 153.705 39.035 153.875 ;
        RECT 39.325 153.705 39.495 153.875 ;
        RECT 39.785 153.705 39.955 153.875 ;
        RECT 40.245 153.705 40.415 153.875 ;
        RECT 40.705 153.705 40.875 153.875 ;
        RECT 41.165 153.705 41.335 153.875 ;
        RECT 41.625 153.705 41.795 153.875 ;
        RECT 42.085 153.705 42.255 153.875 ;
        RECT 42.545 153.705 42.715 153.875 ;
        RECT 43.005 153.705 43.175 153.875 ;
        RECT 43.465 153.705 43.635 153.875 ;
        RECT 43.925 153.705 44.095 153.875 ;
        RECT 44.385 153.705 44.555 153.875 ;
        RECT 44.845 153.705 45.015 153.875 ;
        RECT 45.305 153.705 45.475 153.875 ;
        RECT 45.765 153.705 45.935 153.875 ;
        RECT 46.225 153.705 46.395 153.875 ;
        RECT 46.685 153.705 46.855 153.875 ;
        RECT 47.145 153.705 47.315 153.875 ;
        RECT 47.605 153.705 47.775 153.875 ;
        RECT 48.065 153.705 48.235 153.875 ;
        RECT 48.525 153.705 48.695 153.875 ;
        RECT 48.985 153.705 49.155 153.875 ;
        RECT 49.445 153.705 49.615 153.875 ;
        RECT 49.905 153.705 50.075 153.875 ;
        RECT 50.365 153.705 50.535 153.875 ;
        RECT 50.825 153.705 50.995 153.875 ;
        RECT 51.285 153.705 51.455 153.875 ;
        RECT 51.745 153.705 51.915 153.875 ;
        RECT 52.205 153.705 52.375 153.875 ;
        RECT 52.665 153.705 52.835 153.875 ;
        RECT 53.125 153.705 53.295 153.875 ;
        RECT 53.585 153.705 53.755 153.875 ;
        RECT 54.045 153.705 54.215 153.875 ;
        RECT 54.505 153.705 54.675 153.875 ;
        RECT 54.965 153.705 55.135 153.875 ;
        RECT 55.425 153.705 55.595 153.875 ;
        RECT 55.885 153.705 56.055 153.875 ;
        RECT 56.345 153.705 56.515 153.875 ;
        RECT 56.805 153.705 56.975 153.875 ;
        RECT 57.265 153.705 57.435 153.875 ;
        RECT 57.725 153.705 57.895 153.875 ;
        RECT 58.185 153.705 58.355 153.875 ;
        RECT 58.645 153.705 58.815 153.875 ;
        RECT 59.105 153.705 59.275 153.875 ;
        RECT 59.565 153.705 59.735 153.875 ;
        RECT 60.025 153.705 60.195 153.875 ;
        RECT 60.485 153.705 60.655 153.875 ;
        RECT 60.945 153.705 61.115 153.875 ;
        RECT 61.405 153.705 61.575 153.875 ;
        RECT 61.865 153.705 62.035 153.875 ;
        RECT 62.325 153.705 62.495 153.875 ;
        RECT 62.785 153.705 62.955 153.875 ;
        RECT 63.245 153.705 63.415 153.875 ;
        RECT 63.705 153.705 63.875 153.875 ;
        RECT 64.165 153.705 64.335 153.875 ;
        RECT 64.625 153.705 64.795 153.875 ;
        RECT 65.085 153.705 65.255 153.875 ;
        RECT 65.545 153.705 65.715 153.875 ;
        RECT 66.005 153.705 66.175 153.875 ;
        RECT 66.465 153.705 66.635 153.875 ;
        RECT 66.925 153.705 67.095 153.875 ;
        RECT 67.385 153.705 67.555 153.875 ;
        RECT 67.845 153.705 68.015 153.875 ;
        RECT 68.305 153.705 68.475 153.875 ;
        RECT 68.765 153.705 68.935 153.875 ;
        RECT 69.225 153.705 69.395 153.875 ;
        RECT 69.685 153.705 69.855 153.875 ;
        RECT 70.145 153.705 70.315 153.875 ;
        RECT 70.605 153.705 70.775 153.875 ;
        RECT 71.065 153.705 71.235 153.875 ;
        RECT 71.525 153.705 71.695 153.875 ;
        RECT 71.985 153.705 72.155 153.875 ;
        RECT 72.445 153.705 72.615 153.875 ;
        RECT 72.905 153.705 73.075 153.875 ;
        RECT 73.365 153.705 73.535 153.875 ;
        RECT 73.825 153.705 73.995 153.875 ;
        RECT 74.285 153.705 74.455 153.875 ;
        RECT 74.745 153.705 74.915 153.875 ;
        RECT 75.205 153.705 75.375 153.875 ;
        RECT 75.665 153.705 75.835 153.875 ;
        RECT 76.125 153.705 76.295 153.875 ;
        RECT 76.585 153.705 76.755 153.875 ;
        RECT 77.045 153.705 77.215 153.875 ;
        RECT 77.505 153.705 77.675 153.875 ;
        RECT 77.965 153.705 78.135 153.875 ;
        RECT 78.425 153.705 78.595 153.875 ;
        RECT 78.885 153.705 79.055 153.875 ;
        RECT 79.345 153.705 79.515 153.875 ;
        RECT 79.805 153.705 79.975 153.875 ;
        RECT 80.265 153.705 80.435 153.875 ;
        RECT 80.725 153.705 80.895 153.875 ;
        RECT 81.185 153.705 81.355 153.875 ;
        RECT 81.645 153.705 81.815 153.875 ;
        RECT 82.105 153.705 82.275 153.875 ;
        RECT 82.565 153.705 82.735 153.875 ;
        RECT 83.025 153.705 83.195 153.875 ;
        RECT 83.485 153.705 83.655 153.875 ;
        RECT 83.945 153.705 84.115 153.875 ;
        RECT 84.405 153.705 84.575 153.875 ;
        RECT 84.865 153.705 85.035 153.875 ;
        RECT 85.325 153.705 85.495 153.875 ;
        RECT 85.785 153.705 85.955 153.875 ;
        RECT 86.245 153.705 86.415 153.875 ;
        RECT 86.705 153.705 86.875 153.875 ;
        RECT 87.165 153.705 87.335 153.875 ;
        RECT 87.625 153.705 87.795 153.875 ;
        RECT 88.085 153.705 88.255 153.875 ;
        RECT 88.545 153.705 88.715 153.875 ;
        RECT 89.005 153.705 89.175 153.875 ;
        RECT 89.465 153.705 89.635 153.875 ;
        RECT 89.925 153.705 90.095 153.875 ;
        RECT 90.385 153.705 90.555 153.875 ;
        RECT 90.845 153.705 91.015 153.875 ;
        RECT 91.305 153.705 91.475 153.875 ;
        RECT 91.765 153.705 91.935 153.875 ;
        RECT 92.225 153.705 92.395 153.875 ;
        RECT 92.685 153.705 92.855 153.875 ;
        RECT 93.145 153.705 93.315 153.875 ;
        RECT 93.605 153.705 93.775 153.875 ;
        RECT 94.065 153.705 94.235 153.875 ;
        RECT 94.525 153.705 94.695 153.875 ;
        RECT 94.985 153.705 95.155 153.875 ;
        RECT 95.445 153.705 95.615 153.875 ;
        RECT 95.905 153.705 96.075 153.875 ;
        RECT 96.365 153.705 96.535 153.875 ;
        RECT 96.825 153.705 96.995 153.875 ;
        RECT 97.285 153.705 97.455 153.875 ;
        RECT 97.745 153.705 97.915 153.875 ;
        RECT 98.205 153.705 98.375 153.875 ;
        RECT 98.665 153.705 98.835 153.875 ;
        RECT 99.125 153.705 99.295 153.875 ;
        RECT 99.585 153.705 99.755 153.875 ;
        RECT 100.045 153.705 100.215 153.875 ;
        RECT 100.505 153.705 100.675 153.875 ;
        RECT 100.965 153.705 101.135 153.875 ;
        RECT 101.425 153.705 101.595 153.875 ;
        RECT 101.885 153.705 102.055 153.875 ;
        RECT 102.345 153.705 102.515 153.875 ;
        RECT 102.805 153.705 102.975 153.875 ;
        RECT 103.265 153.705 103.435 153.875 ;
        RECT 103.725 153.705 103.895 153.875 ;
        RECT 104.185 153.705 104.355 153.875 ;
        RECT 104.645 153.705 104.815 153.875 ;
        RECT 105.105 153.705 105.275 153.875 ;
        RECT 105.565 153.705 105.735 153.875 ;
        RECT 106.025 153.705 106.195 153.875 ;
        RECT 106.485 153.705 106.655 153.875 ;
        RECT 106.945 153.705 107.115 153.875 ;
        RECT 107.405 153.705 107.575 153.875 ;
        RECT 107.865 153.705 108.035 153.875 ;
        RECT 108.325 153.705 108.495 153.875 ;
        RECT 108.785 153.705 108.955 153.875 ;
        RECT 109.245 153.705 109.415 153.875 ;
        RECT 109.705 153.705 109.875 153.875 ;
        RECT 110.165 153.705 110.335 153.875 ;
        RECT 110.625 153.705 110.795 153.875 ;
        RECT 111.085 153.705 111.255 153.875 ;
        RECT 111.545 153.705 111.715 153.875 ;
        RECT 112.005 153.705 112.175 153.875 ;
        RECT 112.465 153.705 112.635 153.875 ;
        RECT 112.925 153.705 113.095 153.875 ;
        RECT 113.385 153.705 113.555 153.875 ;
        RECT 113.845 153.705 114.015 153.875 ;
        RECT 114.305 153.705 114.475 153.875 ;
        RECT 114.765 153.705 114.935 153.875 ;
        RECT 115.225 153.705 115.395 153.875 ;
        RECT 115.685 153.705 115.855 153.875 ;
        RECT 116.145 153.705 116.315 153.875 ;
        RECT 116.605 153.705 116.775 153.875 ;
        RECT 117.065 153.705 117.235 153.875 ;
        RECT 117.525 153.705 117.695 153.875 ;
        RECT 117.985 153.705 118.155 153.875 ;
        RECT 118.445 153.705 118.615 153.875 ;
        RECT 118.905 153.705 119.075 153.875 ;
        RECT 119.365 153.705 119.535 153.875 ;
        RECT 119.825 153.705 119.995 153.875 ;
        RECT 120.285 153.705 120.455 153.875 ;
        RECT 120.745 153.705 120.915 153.875 ;
        RECT 121.205 153.705 121.375 153.875 ;
        RECT 121.665 153.705 121.835 153.875 ;
        RECT 122.125 153.705 122.295 153.875 ;
        RECT 122.585 153.705 122.755 153.875 ;
        RECT 123.045 153.705 123.215 153.875 ;
        RECT 123.505 153.705 123.675 153.875 ;
        RECT 123.965 153.705 124.135 153.875 ;
        RECT 124.425 153.705 124.595 153.875 ;
        RECT 124.885 153.705 125.055 153.875 ;
        RECT 125.345 153.705 125.515 153.875 ;
        RECT 125.805 153.705 125.975 153.875 ;
        RECT 126.265 153.705 126.435 153.875 ;
        RECT 126.725 153.705 126.895 153.875 ;
        RECT 127.185 153.705 127.355 153.875 ;
        RECT 127.645 153.705 127.815 153.875 ;
        RECT 128.105 153.705 128.275 153.875 ;
        RECT 128.565 153.705 128.735 153.875 ;
        RECT 129.025 153.705 129.195 153.875 ;
        RECT 129.485 153.705 129.655 153.875 ;
        RECT 129.945 153.705 130.115 153.875 ;
        RECT 130.405 153.705 130.575 153.875 ;
        RECT 130.865 153.705 131.035 153.875 ;
        RECT 131.325 153.705 131.495 153.875 ;
        RECT 131.785 153.705 131.955 153.875 ;
        RECT 132.245 153.705 132.415 153.875 ;
        RECT 132.705 153.705 132.875 153.875 ;
        RECT 133.165 153.705 133.335 153.875 ;
        RECT 133.625 153.705 133.795 153.875 ;
        RECT 134.085 153.705 134.255 153.875 ;
        RECT 134.545 153.705 134.715 153.875 ;
        RECT 135.005 153.705 135.175 153.875 ;
        RECT 135.465 153.705 135.635 153.875 ;
        RECT 135.925 153.705 136.095 153.875 ;
        RECT 136.385 153.705 136.555 153.875 ;
        RECT 136.845 153.705 137.015 153.875 ;
        RECT 137.305 153.705 137.475 153.875 ;
        RECT 137.765 153.705 137.935 153.875 ;
        RECT 138.225 153.705 138.395 153.875 ;
        RECT 138.685 153.705 138.855 153.875 ;
        RECT 139.145 153.705 139.315 153.875 ;
        RECT 139.605 153.705 139.775 153.875 ;
        RECT 140.065 153.705 140.235 153.875 ;
        RECT 140.525 153.705 140.695 153.875 ;
        RECT 140.985 153.705 141.155 153.875 ;
        RECT 141.445 153.705 141.615 153.875 ;
        RECT 141.905 153.705 142.075 153.875 ;
        RECT 142.365 153.705 142.535 153.875 ;
        RECT 142.825 153.705 142.995 153.875 ;
        RECT 143.285 153.705 143.455 153.875 ;
        RECT 143.745 153.705 143.915 153.875 ;
        RECT 144.205 153.705 144.375 153.875 ;
        RECT 144.665 153.705 144.835 153.875 ;
        RECT 145.125 153.705 145.295 153.875 ;
        RECT 145.585 153.705 145.755 153.875 ;
        RECT 146.045 153.705 146.215 153.875 ;
        RECT 146.505 153.705 146.675 153.875 ;
        RECT 146.965 153.705 147.135 153.875 ;
        RECT 147.425 153.705 147.595 153.875 ;
        RECT 147.885 153.705 148.055 153.875 ;
        RECT 148.345 153.705 148.515 153.875 ;
        RECT 148.805 153.705 148.975 153.875 ;
        RECT 149.265 153.705 149.435 153.875 ;
        RECT 149.725 153.705 149.895 153.875 ;
        RECT 150.185 153.705 150.355 153.875 ;
        RECT 16.350 152.855 16.520 153.025 ;
        RECT 15.865 152.175 16.035 152.345 ;
        RECT 16.745 152.515 16.915 152.685 ;
        RECT 17.200 152.175 17.370 152.345 ;
        RECT 18.450 152.855 18.620 153.025 ;
        RECT 17.935 152.515 18.105 152.685 ;
        RECT 20.020 152.855 20.190 153.025 ;
        RECT 20.455 152.515 20.625 152.685 ;
        RECT 22.765 152.855 22.935 153.025 ;
        RECT 26.905 153.195 27.075 153.365 ;
        RECT 25.065 152.515 25.235 152.685 ;
        RECT 25.525 152.175 25.695 152.345 ;
        RECT 30.585 152.175 30.755 152.345 ;
        RECT 31.045 152.175 31.215 152.345 ;
        RECT 32.425 152.175 32.595 152.345 ;
        RECT 31.505 151.835 31.675 152.005 ;
        RECT 29.665 151.495 29.835 151.665 ;
        RECT 42.545 153.195 42.715 153.365 ;
        RECT 44.845 153.195 45.015 153.365 ;
        RECT 41.625 152.175 41.795 152.345 ;
        RECT 42.085 151.835 42.255 152.005 ;
        RECT 44.385 152.175 44.555 152.345 ;
        RECT 43.005 151.835 43.175 152.005 ;
        RECT 45.305 152.175 45.475 152.345 ;
        RECT 55.425 153.195 55.595 153.365 ;
        RECT 52.665 152.175 52.835 152.345 ;
        RECT 53.125 152.175 53.295 152.345 ;
        RECT 54.045 152.175 54.215 152.345 ;
        RECT 54.505 152.175 54.675 152.345 ;
        RECT 57.725 151.495 57.895 151.665 ;
        RECT 60.035 152.515 60.205 152.685 ;
        RECT 60.470 152.855 60.640 153.025 ;
        RECT 62.040 152.855 62.210 153.025 ;
        RECT 62.555 152.515 62.725 152.685 ;
        RECT 63.290 152.175 63.460 152.345 ;
        RECT 63.745 152.515 63.915 152.685 ;
        RECT 64.140 152.855 64.310 153.025 ;
        RECT 64.625 152.175 64.795 152.345 ;
        RECT 67.385 152.515 67.555 152.685 ;
        RECT 66.465 152.175 66.635 152.345 ;
        RECT 65.545 151.495 65.715 151.665 ;
        RECT 72.905 152.175 73.075 152.345 ;
        RECT 73.825 152.175 73.995 152.345 ;
        RECT 71.985 151.495 72.155 151.665 ;
        RECT 74.285 152.175 74.455 152.345 ;
        RECT 77.045 152.175 77.215 152.345 ;
        RECT 76.585 151.495 76.755 151.665 ;
        RECT 78.885 152.515 79.055 152.685 ;
        RECT 78.425 152.175 78.595 152.345 ;
        RECT 80.265 152.855 80.435 153.025 ;
        RECT 84.865 153.195 85.035 153.365 ;
        RECT 87.165 152.855 87.335 153.025 ;
        RECT 83.945 152.175 84.115 152.345 ;
        RECT 84.405 152.175 84.575 152.345 ;
        RECT 85.785 152.175 85.955 152.345 ;
        RECT 85.325 151.835 85.495 152.005 ;
        RECT 86.245 151.495 86.415 151.665 ;
        RECT 87.165 152.175 87.335 152.345 ;
        RECT 92.225 153.195 92.395 153.365 ;
        RECT 95.905 153.195 96.075 153.365 ;
        RECT 98.205 153.195 98.375 153.365 ;
        RECT 93.605 152.175 93.775 152.345 ;
        RECT 94.065 152.175 94.235 152.345 ;
        RECT 94.525 152.175 94.695 152.345 ;
        RECT 95.325 152.175 95.495 152.345 ;
        RECT 96.735 152.175 96.905 152.345 ;
        RECT 97.745 152.175 97.915 152.345 ;
        RECT 99.125 151.835 99.295 152.005 ;
        RECT 108.325 153.195 108.495 153.365 ;
        RECT 111.085 152.855 111.255 153.025 ;
        RECT 101.885 152.175 102.055 152.345 ;
        RECT 113.395 152.515 113.565 152.685 ;
        RECT 113.830 152.855 114.000 153.025 ;
        RECT 115.400 152.855 115.570 153.025 ;
        RECT 115.915 152.515 116.085 152.685 ;
        RECT 116.650 151.835 116.820 152.005 ;
        RECT 117.105 152.515 117.275 152.685 ;
        RECT 117.500 152.855 117.670 153.025 ;
        RECT 117.985 152.515 118.155 152.685 ;
        RECT 11.265 150.985 11.435 151.155 ;
        RECT 11.725 150.985 11.895 151.155 ;
        RECT 12.185 150.985 12.355 151.155 ;
        RECT 12.645 150.985 12.815 151.155 ;
        RECT 13.105 150.985 13.275 151.155 ;
        RECT 13.565 150.985 13.735 151.155 ;
        RECT 14.025 150.985 14.195 151.155 ;
        RECT 14.485 150.985 14.655 151.155 ;
        RECT 14.945 150.985 15.115 151.155 ;
        RECT 15.405 150.985 15.575 151.155 ;
        RECT 15.865 150.985 16.035 151.155 ;
        RECT 16.325 150.985 16.495 151.155 ;
        RECT 16.785 150.985 16.955 151.155 ;
        RECT 17.245 150.985 17.415 151.155 ;
        RECT 17.705 150.985 17.875 151.155 ;
        RECT 18.165 150.985 18.335 151.155 ;
        RECT 18.625 150.985 18.795 151.155 ;
        RECT 19.085 150.985 19.255 151.155 ;
        RECT 19.545 150.985 19.715 151.155 ;
        RECT 20.005 150.985 20.175 151.155 ;
        RECT 20.465 150.985 20.635 151.155 ;
        RECT 20.925 150.985 21.095 151.155 ;
        RECT 21.385 150.985 21.555 151.155 ;
        RECT 21.845 150.985 22.015 151.155 ;
        RECT 22.305 150.985 22.475 151.155 ;
        RECT 22.765 150.985 22.935 151.155 ;
        RECT 23.225 150.985 23.395 151.155 ;
        RECT 23.685 150.985 23.855 151.155 ;
        RECT 24.145 150.985 24.315 151.155 ;
        RECT 24.605 150.985 24.775 151.155 ;
        RECT 25.065 150.985 25.235 151.155 ;
        RECT 25.525 150.985 25.695 151.155 ;
        RECT 25.985 150.985 26.155 151.155 ;
        RECT 26.445 150.985 26.615 151.155 ;
        RECT 26.905 150.985 27.075 151.155 ;
        RECT 27.365 150.985 27.535 151.155 ;
        RECT 27.825 150.985 27.995 151.155 ;
        RECT 28.285 150.985 28.455 151.155 ;
        RECT 28.745 150.985 28.915 151.155 ;
        RECT 29.205 150.985 29.375 151.155 ;
        RECT 29.665 150.985 29.835 151.155 ;
        RECT 30.125 150.985 30.295 151.155 ;
        RECT 30.585 150.985 30.755 151.155 ;
        RECT 31.045 150.985 31.215 151.155 ;
        RECT 31.505 150.985 31.675 151.155 ;
        RECT 31.965 150.985 32.135 151.155 ;
        RECT 32.425 150.985 32.595 151.155 ;
        RECT 32.885 150.985 33.055 151.155 ;
        RECT 33.345 150.985 33.515 151.155 ;
        RECT 33.805 150.985 33.975 151.155 ;
        RECT 34.265 150.985 34.435 151.155 ;
        RECT 34.725 150.985 34.895 151.155 ;
        RECT 35.185 150.985 35.355 151.155 ;
        RECT 35.645 150.985 35.815 151.155 ;
        RECT 36.105 150.985 36.275 151.155 ;
        RECT 36.565 150.985 36.735 151.155 ;
        RECT 37.025 150.985 37.195 151.155 ;
        RECT 37.485 150.985 37.655 151.155 ;
        RECT 37.945 150.985 38.115 151.155 ;
        RECT 38.405 150.985 38.575 151.155 ;
        RECT 38.865 150.985 39.035 151.155 ;
        RECT 39.325 150.985 39.495 151.155 ;
        RECT 39.785 150.985 39.955 151.155 ;
        RECT 40.245 150.985 40.415 151.155 ;
        RECT 40.705 150.985 40.875 151.155 ;
        RECT 41.165 150.985 41.335 151.155 ;
        RECT 41.625 150.985 41.795 151.155 ;
        RECT 42.085 150.985 42.255 151.155 ;
        RECT 42.545 150.985 42.715 151.155 ;
        RECT 43.005 150.985 43.175 151.155 ;
        RECT 43.465 150.985 43.635 151.155 ;
        RECT 43.925 150.985 44.095 151.155 ;
        RECT 44.385 150.985 44.555 151.155 ;
        RECT 44.845 150.985 45.015 151.155 ;
        RECT 45.305 150.985 45.475 151.155 ;
        RECT 45.765 150.985 45.935 151.155 ;
        RECT 46.225 150.985 46.395 151.155 ;
        RECT 46.685 150.985 46.855 151.155 ;
        RECT 47.145 150.985 47.315 151.155 ;
        RECT 47.605 150.985 47.775 151.155 ;
        RECT 48.065 150.985 48.235 151.155 ;
        RECT 48.525 150.985 48.695 151.155 ;
        RECT 48.985 150.985 49.155 151.155 ;
        RECT 49.445 150.985 49.615 151.155 ;
        RECT 49.905 150.985 50.075 151.155 ;
        RECT 50.365 150.985 50.535 151.155 ;
        RECT 50.825 150.985 50.995 151.155 ;
        RECT 51.285 150.985 51.455 151.155 ;
        RECT 51.745 150.985 51.915 151.155 ;
        RECT 52.205 150.985 52.375 151.155 ;
        RECT 52.665 150.985 52.835 151.155 ;
        RECT 53.125 150.985 53.295 151.155 ;
        RECT 53.585 150.985 53.755 151.155 ;
        RECT 54.045 150.985 54.215 151.155 ;
        RECT 54.505 150.985 54.675 151.155 ;
        RECT 54.965 150.985 55.135 151.155 ;
        RECT 55.425 150.985 55.595 151.155 ;
        RECT 55.885 150.985 56.055 151.155 ;
        RECT 56.345 150.985 56.515 151.155 ;
        RECT 56.805 150.985 56.975 151.155 ;
        RECT 57.265 150.985 57.435 151.155 ;
        RECT 57.725 150.985 57.895 151.155 ;
        RECT 58.185 150.985 58.355 151.155 ;
        RECT 58.645 150.985 58.815 151.155 ;
        RECT 59.105 150.985 59.275 151.155 ;
        RECT 59.565 150.985 59.735 151.155 ;
        RECT 60.025 150.985 60.195 151.155 ;
        RECT 60.485 150.985 60.655 151.155 ;
        RECT 60.945 150.985 61.115 151.155 ;
        RECT 61.405 150.985 61.575 151.155 ;
        RECT 61.865 150.985 62.035 151.155 ;
        RECT 62.325 150.985 62.495 151.155 ;
        RECT 62.785 150.985 62.955 151.155 ;
        RECT 63.245 150.985 63.415 151.155 ;
        RECT 63.705 150.985 63.875 151.155 ;
        RECT 64.165 150.985 64.335 151.155 ;
        RECT 64.625 150.985 64.795 151.155 ;
        RECT 65.085 150.985 65.255 151.155 ;
        RECT 65.545 150.985 65.715 151.155 ;
        RECT 66.005 150.985 66.175 151.155 ;
        RECT 66.465 150.985 66.635 151.155 ;
        RECT 66.925 150.985 67.095 151.155 ;
        RECT 67.385 150.985 67.555 151.155 ;
        RECT 67.845 150.985 68.015 151.155 ;
        RECT 68.305 150.985 68.475 151.155 ;
        RECT 68.765 150.985 68.935 151.155 ;
        RECT 69.225 150.985 69.395 151.155 ;
        RECT 69.685 150.985 69.855 151.155 ;
        RECT 70.145 150.985 70.315 151.155 ;
        RECT 70.605 150.985 70.775 151.155 ;
        RECT 71.065 150.985 71.235 151.155 ;
        RECT 71.525 150.985 71.695 151.155 ;
        RECT 71.985 150.985 72.155 151.155 ;
        RECT 72.445 150.985 72.615 151.155 ;
        RECT 72.905 150.985 73.075 151.155 ;
        RECT 73.365 150.985 73.535 151.155 ;
        RECT 73.825 150.985 73.995 151.155 ;
        RECT 74.285 150.985 74.455 151.155 ;
        RECT 74.745 150.985 74.915 151.155 ;
        RECT 75.205 150.985 75.375 151.155 ;
        RECT 75.665 150.985 75.835 151.155 ;
        RECT 76.125 150.985 76.295 151.155 ;
        RECT 76.585 150.985 76.755 151.155 ;
        RECT 77.045 150.985 77.215 151.155 ;
        RECT 77.505 150.985 77.675 151.155 ;
        RECT 77.965 150.985 78.135 151.155 ;
        RECT 78.425 150.985 78.595 151.155 ;
        RECT 78.885 150.985 79.055 151.155 ;
        RECT 79.345 150.985 79.515 151.155 ;
        RECT 79.805 150.985 79.975 151.155 ;
        RECT 80.265 150.985 80.435 151.155 ;
        RECT 80.725 150.985 80.895 151.155 ;
        RECT 81.185 150.985 81.355 151.155 ;
        RECT 81.645 150.985 81.815 151.155 ;
        RECT 82.105 150.985 82.275 151.155 ;
        RECT 82.565 150.985 82.735 151.155 ;
        RECT 83.025 150.985 83.195 151.155 ;
        RECT 83.485 150.985 83.655 151.155 ;
        RECT 83.945 150.985 84.115 151.155 ;
        RECT 84.405 150.985 84.575 151.155 ;
        RECT 84.865 150.985 85.035 151.155 ;
        RECT 85.325 150.985 85.495 151.155 ;
        RECT 85.785 150.985 85.955 151.155 ;
        RECT 86.245 150.985 86.415 151.155 ;
        RECT 86.705 150.985 86.875 151.155 ;
        RECT 87.165 150.985 87.335 151.155 ;
        RECT 87.625 150.985 87.795 151.155 ;
        RECT 88.085 150.985 88.255 151.155 ;
        RECT 88.545 150.985 88.715 151.155 ;
        RECT 89.005 150.985 89.175 151.155 ;
        RECT 89.465 150.985 89.635 151.155 ;
        RECT 89.925 150.985 90.095 151.155 ;
        RECT 90.385 150.985 90.555 151.155 ;
        RECT 90.845 150.985 91.015 151.155 ;
        RECT 91.305 150.985 91.475 151.155 ;
        RECT 91.765 150.985 91.935 151.155 ;
        RECT 92.225 150.985 92.395 151.155 ;
        RECT 92.685 150.985 92.855 151.155 ;
        RECT 93.145 150.985 93.315 151.155 ;
        RECT 93.605 150.985 93.775 151.155 ;
        RECT 94.065 150.985 94.235 151.155 ;
        RECT 94.525 150.985 94.695 151.155 ;
        RECT 94.985 150.985 95.155 151.155 ;
        RECT 95.445 150.985 95.615 151.155 ;
        RECT 95.905 150.985 96.075 151.155 ;
        RECT 96.365 150.985 96.535 151.155 ;
        RECT 96.825 150.985 96.995 151.155 ;
        RECT 97.285 150.985 97.455 151.155 ;
        RECT 97.745 150.985 97.915 151.155 ;
        RECT 98.205 150.985 98.375 151.155 ;
        RECT 98.665 150.985 98.835 151.155 ;
        RECT 99.125 150.985 99.295 151.155 ;
        RECT 99.585 150.985 99.755 151.155 ;
        RECT 100.045 150.985 100.215 151.155 ;
        RECT 100.505 150.985 100.675 151.155 ;
        RECT 100.965 150.985 101.135 151.155 ;
        RECT 101.425 150.985 101.595 151.155 ;
        RECT 101.885 150.985 102.055 151.155 ;
        RECT 102.345 150.985 102.515 151.155 ;
        RECT 102.805 150.985 102.975 151.155 ;
        RECT 103.265 150.985 103.435 151.155 ;
        RECT 103.725 150.985 103.895 151.155 ;
        RECT 104.185 150.985 104.355 151.155 ;
        RECT 104.645 150.985 104.815 151.155 ;
        RECT 105.105 150.985 105.275 151.155 ;
        RECT 105.565 150.985 105.735 151.155 ;
        RECT 106.025 150.985 106.195 151.155 ;
        RECT 106.485 150.985 106.655 151.155 ;
        RECT 106.945 150.985 107.115 151.155 ;
        RECT 107.405 150.985 107.575 151.155 ;
        RECT 107.865 150.985 108.035 151.155 ;
        RECT 108.325 150.985 108.495 151.155 ;
        RECT 108.785 150.985 108.955 151.155 ;
        RECT 109.245 150.985 109.415 151.155 ;
        RECT 109.705 150.985 109.875 151.155 ;
        RECT 110.165 150.985 110.335 151.155 ;
        RECT 110.625 150.985 110.795 151.155 ;
        RECT 111.085 150.985 111.255 151.155 ;
        RECT 111.545 150.985 111.715 151.155 ;
        RECT 112.005 150.985 112.175 151.155 ;
        RECT 112.465 150.985 112.635 151.155 ;
        RECT 112.925 150.985 113.095 151.155 ;
        RECT 113.385 150.985 113.555 151.155 ;
        RECT 113.845 150.985 114.015 151.155 ;
        RECT 114.305 150.985 114.475 151.155 ;
        RECT 114.765 150.985 114.935 151.155 ;
        RECT 115.225 150.985 115.395 151.155 ;
        RECT 115.685 150.985 115.855 151.155 ;
        RECT 116.145 150.985 116.315 151.155 ;
        RECT 116.605 150.985 116.775 151.155 ;
        RECT 117.065 150.985 117.235 151.155 ;
        RECT 117.525 150.985 117.695 151.155 ;
        RECT 117.985 150.985 118.155 151.155 ;
        RECT 118.445 150.985 118.615 151.155 ;
        RECT 118.905 150.985 119.075 151.155 ;
        RECT 119.365 150.985 119.535 151.155 ;
        RECT 119.825 150.985 119.995 151.155 ;
        RECT 120.285 150.985 120.455 151.155 ;
        RECT 120.745 150.985 120.915 151.155 ;
        RECT 121.205 150.985 121.375 151.155 ;
        RECT 121.665 150.985 121.835 151.155 ;
        RECT 122.125 150.985 122.295 151.155 ;
        RECT 122.585 150.985 122.755 151.155 ;
        RECT 123.045 150.985 123.215 151.155 ;
        RECT 123.505 150.985 123.675 151.155 ;
        RECT 123.965 150.985 124.135 151.155 ;
        RECT 124.425 150.985 124.595 151.155 ;
        RECT 124.885 150.985 125.055 151.155 ;
        RECT 125.345 150.985 125.515 151.155 ;
        RECT 125.805 150.985 125.975 151.155 ;
        RECT 126.265 150.985 126.435 151.155 ;
        RECT 126.725 150.985 126.895 151.155 ;
        RECT 127.185 150.985 127.355 151.155 ;
        RECT 127.645 150.985 127.815 151.155 ;
        RECT 128.105 150.985 128.275 151.155 ;
        RECT 128.565 150.985 128.735 151.155 ;
        RECT 129.025 150.985 129.195 151.155 ;
        RECT 129.485 150.985 129.655 151.155 ;
        RECT 129.945 150.985 130.115 151.155 ;
        RECT 130.405 150.985 130.575 151.155 ;
        RECT 130.865 150.985 131.035 151.155 ;
        RECT 131.325 150.985 131.495 151.155 ;
        RECT 131.785 150.985 131.955 151.155 ;
        RECT 132.245 150.985 132.415 151.155 ;
        RECT 132.705 150.985 132.875 151.155 ;
        RECT 133.165 150.985 133.335 151.155 ;
        RECT 133.625 150.985 133.795 151.155 ;
        RECT 134.085 150.985 134.255 151.155 ;
        RECT 134.545 150.985 134.715 151.155 ;
        RECT 135.005 150.985 135.175 151.155 ;
        RECT 135.465 150.985 135.635 151.155 ;
        RECT 135.925 150.985 136.095 151.155 ;
        RECT 136.385 150.985 136.555 151.155 ;
        RECT 136.845 150.985 137.015 151.155 ;
        RECT 137.305 150.985 137.475 151.155 ;
        RECT 137.765 150.985 137.935 151.155 ;
        RECT 138.225 150.985 138.395 151.155 ;
        RECT 138.685 150.985 138.855 151.155 ;
        RECT 139.145 150.985 139.315 151.155 ;
        RECT 139.605 150.985 139.775 151.155 ;
        RECT 140.065 150.985 140.235 151.155 ;
        RECT 140.525 150.985 140.695 151.155 ;
        RECT 140.985 150.985 141.155 151.155 ;
        RECT 141.445 150.985 141.615 151.155 ;
        RECT 141.905 150.985 142.075 151.155 ;
        RECT 142.365 150.985 142.535 151.155 ;
        RECT 142.825 150.985 142.995 151.155 ;
        RECT 143.285 150.985 143.455 151.155 ;
        RECT 143.745 150.985 143.915 151.155 ;
        RECT 144.205 150.985 144.375 151.155 ;
        RECT 144.665 150.985 144.835 151.155 ;
        RECT 145.125 150.985 145.295 151.155 ;
        RECT 145.585 150.985 145.755 151.155 ;
        RECT 146.045 150.985 146.215 151.155 ;
        RECT 146.505 150.985 146.675 151.155 ;
        RECT 146.965 150.985 147.135 151.155 ;
        RECT 147.425 150.985 147.595 151.155 ;
        RECT 147.885 150.985 148.055 151.155 ;
        RECT 148.345 150.985 148.515 151.155 ;
        RECT 148.805 150.985 148.975 151.155 ;
        RECT 149.265 150.985 149.435 151.155 ;
        RECT 149.725 150.985 149.895 151.155 ;
        RECT 150.185 150.985 150.355 151.155 ;
        RECT 19.085 150.475 19.255 150.645 ;
        RECT 20.005 149.795 20.175 149.965 ;
        RECT 20.925 149.455 21.095 149.625 ;
        RECT 31.965 149.115 32.135 149.285 ;
        RECT 33.805 149.795 33.975 149.965 ;
        RECT 34.265 149.455 34.435 149.625 ;
        RECT 39.325 150.135 39.495 150.305 ;
        RECT 41.625 150.475 41.795 150.645 ;
        RECT 38.815 149.795 38.985 149.965 ;
        RECT 39.785 149.795 39.955 149.965 ;
        RECT 41.165 149.795 41.335 149.965 ;
        RECT 42.085 149.795 42.255 149.965 ;
        RECT 51.285 149.455 51.455 149.625 ;
        RECT 53.125 149.455 53.295 149.625 ;
        RECT 53.585 149.795 53.755 149.965 ;
        RECT 74.745 150.475 74.915 150.645 ;
        RECT 54.505 148.775 54.675 148.945 ;
        RECT 74.745 149.455 74.915 149.625 ;
        RECT 75.665 149.795 75.835 149.965 ;
        RECT 76.125 149.795 76.295 149.965 ;
        RECT 93.145 149.795 93.315 149.965 ;
        RECT 94.525 149.795 94.695 149.965 ;
        RECT 94.985 149.795 95.155 149.965 ;
        RECT 96.825 149.455 96.995 149.625 ;
        RECT 98.205 149.795 98.375 149.965 ;
        RECT 97.285 149.115 97.455 149.285 ;
        RECT 97.745 148.775 97.915 148.945 ;
        RECT 101.885 149.455 102.055 149.625 ;
        RECT 103.725 149.795 103.895 149.965 ;
        RECT 103.265 149.455 103.435 149.625 ;
        RECT 106.025 149.795 106.195 149.965 ;
        RECT 109.245 150.475 109.415 150.645 ;
        RECT 106.945 149.795 107.115 149.965 ;
        RECT 107.405 149.795 107.575 149.965 ;
        RECT 107.865 149.795 108.035 149.965 ;
        RECT 109.705 149.795 109.875 149.965 ;
        RECT 111.545 149.795 111.715 149.965 ;
        RECT 112.925 149.795 113.095 149.965 ;
        RECT 114.765 149.795 114.935 149.965 ;
        RECT 110.165 148.775 110.335 148.945 ;
        RECT 113.385 149.455 113.555 149.625 ;
        RECT 115.685 149.115 115.855 149.285 ;
        RECT 116.605 148.775 116.775 148.945 ;
        RECT 118.915 149.455 119.085 149.625 ;
        RECT 119.350 149.115 119.520 149.285 ;
        RECT 121.435 149.455 121.605 149.625 ;
        RECT 120.920 149.115 121.090 149.285 ;
        RECT 122.170 149.795 122.340 149.965 ;
        RECT 122.625 149.455 122.795 149.625 ;
        RECT 123.505 149.795 123.675 149.965 ;
        RECT 123.020 149.115 123.190 149.285 ;
        RECT 11.265 148.265 11.435 148.435 ;
        RECT 11.725 148.265 11.895 148.435 ;
        RECT 12.185 148.265 12.355 148.435 ;
        RECT 12.645 148.265 12.815 148.435 ;
        RECT 13.105 148.265 13.275 148.435 ;
        RECT 13.565 148.265 13.735 148.435 ;
        RECT 14.025 148.265 14.195 148.435 ;
        RECT 14.485 148.265 14.655 148.435 ;
        RECT 14.945 148.265 15.115 148.435 ;
        RECT 15.405 148.265 15.575 148.435 ;
        RECT 15.865 148.265 16.035 148.435 ;
        RECT 16.325 148.265 16.495 148.435 ;
        RECT 16.785 148.265 16.955 148.435 ;
        RECT 17.245 148.265 17.415 148.435 ;
        RECT 17.705 148.265 17.875 148.435 ;
        RECT 18.165 148.265 18.335 148.435 ;
        RECT 18.625 148.265 18.795 148.435 ;
        RECT 19.085 148.265 19.255 148.435 ;
        RECT 19.545 148.265 19.715 148.435 ;
        RECT 20.005 148.265 20.175 148.435 ;
        RECT 20.465 148.265 20.635 148.435 ;
        RECT 20.925 148.265 21.095 148.435 ;
        RECT 21.385 148.265 21.555 148.435 ;
        RECT 21.845 148.265 22.015 148.435 ;
        RECT 22.305 148.265 22.475 148.435 ;
        RECT 22.765 148.265 22.935 148.435 ;
        RECT 23.225 148.265 23.395 148.435 ;
        RECT 23.685 148.265 23.855 148.435 ;
        RECT 24.145 148.265 24.315 148.435 ;
        RECT 24.605 148.265 24.775 148.435 ;
        RECT 25.065 148.265 25.235 148.435 ;
        RECT 25.525 148.265 25.695 148.435 ;
        RECT 25.985 148.265 26.155 148.435 ;
        RECT 26.445 148.265 26.615 148.435 ;
        RECT 26.905 148.265 27.075 148.435 ;
        RECT 27.365 148.265 27.535 148.435 ;
        RECT 27.825 148.265 27.995 148.435 ;
        RECT 28.285 148.265 28.455 148.435 ;
        RECT 28.745 148.265 28.915 148.435 ;
        RECT 29.205 148.265 29.375 148.435 ;
        RECT 29.665 148.265 29.835 148.435 ;
        RECT 30.125 148.265 30.295 148.435 ;
        RECT 30.585 148.265 30.755 148.435 ;
        RECT 31.045 148.265 31.215 148.435 ;
        RECT 31.505 148.265 31.675 148.435 ;
        RECT 31.965 148.265 32.135 148.435 ;
        RECT 32.425 148.265 32.595 148.435 ;
        RECT 32.885 148.265 33.055 148.435 ;
        RECT 33.345 148.265 33.515 148.435 ;
        RECT 33.805 148.265 33.975 148.435 ;
        RECT 34.265 148.265 34.435 148.435 ;
        RECT 34.725 148.265 34.895 148.435 ;
        RECT 35.185 148.265 35.355 148.435 ;
        RECT 35.645 148.265 35.815 148.435 ;
        RECT 36.105 148.265 36.275 148.435 ;
        RECT 36.565 148.265 36.735 148.435 ;
        RECT 37.025 148.265 37.195 148.435 ;
        RECT 37.485 148.265 37.655 148.435 ;
        RECT 37.945 148.265 38.115 148.435 ;
        RECT 38.405 148.265 38.575 148.435 ;
        RECT 38.865 148.265 39.035 148.435 ;
        RECT 39.325 148.265 39.495 148.435 ;
        RECT 39.785 148.265 39.955 148.435 ;
        RECT 40.245 148.265 40.415 148.435 ;
        RECT 40.705 148.265 40.875 148.435 ;
        RECT 41.165 148.265 41.335 148.435 ;
        RECT 41.625 148.265 41.795 148.435 ;
        RECT 42.085 148.265 42.255 148.435 ;
        RECT 42.545 148.265 42.715 148.435 ;
        RECT 43.005 148.265 43.175 148.435 ;
        RECT 43.465 148.265 43.635 148.435 ;
        RECT 43.925 148.265 44.095 148.435 ;
        RECT 44.385 148.265 44.555 148.435 ;
        RECT 44.845 148.265 45.015 148.435 ;
        RECT 45.305 148.265 45.475 148.435 ;
        RECT 45.765 148.265 45.935 148.435 ;
        RECT 46.225 148.265 46.395 148.435 ;
        RECT 46.685 148.265 46.855 148.435 ;
        RECT 47.145 148.265 47.315 148.435 ;
        RECT 47.605 148.265 47.775 148.435 ;
        RECT 48.065 148.265 48.235 148.435 ;
        RECT 48.525 148.265 48.695 148.435 ;
        RECT 48.985 148.265 49.155 148.435 ;
        RECT 49.445 148.265 49.615 148.435 ;
        RECT 49.905 148.265 50.075 148.435 ;
        RECT 50.365 148.265 50.535 148.435 ;
        RECT 50.825 148.265 50.995 148.435 ;
        RECT 51.285 148.265 51.455 148.435 ;
        RECT 51.745 148.265 51.915 148.435 ;
        RECT 52.205 148.265 52.375 148.435 ;
        RECT 52.665 148.265 52.835 148.435 ;
        RECT 53.125 148.265 53.295 148.435 ;
        RECT 53.585 148.265 53.755 148.435 ;
        RECT 54.045 148.265 54.215 148.435 ;
        RECT 54.505 148.265 54.675 148.435 ;
        RECT 54.965 148.265 55.135 148.435 ;
        RECT 55.425 148.265 55.595 148.435 ;
        RECT 55.885 148.265 56.055 148.435 ;
        RECT 56.345 148.265 56.515 148.435 ;
        RECT 56.805 148.265 56.975 148.435 ;
        RECT 57.265 148.265 57.435 148.435 ;
        RECT 57.725 148.265 57.895 148.435 ;
        RECT 58.185 148.265 58.355 148.435 ;
        RECT 58.645 148.265 58.815 148.435 ;
        RECT 59.105 148.265 59.275 148.435 ;
        RECT 59.565 148.265 59.735 148.435 ;
        RECT 60.025 148.265 60.195 148.435 ;
        RECT 60.485 148.265 60.655 148.435 ;
        RECT 60.945 148.265 61.115 148.435 ;
        RECT 61.405 148.265 61.575 148.435 ;
        RECT 61.865 148.265 62.035 148.435 ;
        RECT 62.325 148.265 62.495 148.435 ;
        RECT 62.785 148.265 62.955 148.435 ;
        RECT 63.245 148.265 63.415 148.435 ;
        RECT 63.705 148.265 63.875 148.435 ;
        RECT 64.165 148.265 64.335 148.435 ;
        RECT 64.625 148.265 64.795 148.435 ;
        RECT 65.085 148.265 65.255 148.435 ;
        RECT 65.545 148.265 65.715 148.435 ;
        RECT 66.005 148.265 66.175 148.435 ;
        RECT 66.465 148.265 66.635 148.435 ;
        RECT 66.925 148.265 67.095 148.435 ;
        RECT 67.385 148.265 67.555 148.435 ;
        RECT 67.845 148.265 68.015 148.435 ;
        RECT 68.305 148.265 68.475 148.435 ;
        RECT 68.765 148.265 68.935 148.435 ;
        RECT 69.225 148.265 69.395 148.435 ;
        RECT 69.685 148.265 69.855 148.435 ;
        RECT 70.145 148.265 70.315 148.435 ;
        RECT 70.605 148.265 70.775 148.435 ;
        RECT 71.065 148.265 71.235 148.435 ;
        RECT 71.525 148.265 71.695 148.435 ;
        RECT 71.985 148.265 72.155 148.435 ;
        RECT 72.445 148.265 72.615 148.435 ;
        RECT 72.905 148.265 73.075 148.435 ;
        RECT 73.365 148.265 73.535 148.435 ;
        RECT 73.825 148.265 73.995 148.435 ;
        RECT 74.285 148.265 74.455 148.435 ;
        RECT 74.745 148.265 74.915 148.435 ;
        RECT 75.205 148.265 75.375 148.435 ;
        RECT 75.665 148.265 75.835 148.435 ;
        RECT 76.125 148.265 76.295 148.435 ;
        RECT 76.585 148.265 76.755 148.435 ;
        RECT 77.045 148.265 77.215 148.435 ;
        RECT 77.505 148.265 77.675 148.435 ;
        RECT 77.965 148.265 78.135 148.435 ;
        RECT 78.425 148.265 78.595 148.435 ;
        RECT 78.885 148.265 79.055 148.435 ;
        RECT 79.345 148.265 79.515 148.435 ;
        RECT 79.805 148.265 79.975 148.435 ;
        RECT 80.265 148.265 80.435 148.435 ;
        RECT 80.725 148.265 80.895 148.435 ;
        RECT 81.185 148.265 81.355 148.435 ;
        RECT 81.645 148.265 81.815 148.435 ;
        RECT 82.105 148.265 82.275 148.435 ;
        RECT 82.565 148.265 82.735 148.435 ;
        RECT 83.025 148.265 83.195 148.435 ;
        RECT 83.485 148.265 83.655 148.435 ;
        RECT 83.945 148.265 84.115 148.435 ;
        RECT 84.405 148.265 84.575 148.435 ;
        RECT 84.865 148.265 85.035 148.435 ;
        RECT 85.325 148.265 85.495 148.435 ;
        RECT 85.785 148.265 85.955 148.435 ;
        RECT 86.245 148.265 86.415 148.435 ;
        RECT 86.705 148.265 86.875 148.435 ;
        RECT 87.165 148.265 87.335 148.435 ;
        RECT 87.625 148.265 87.795 148.435 ;
        RECT 88.085 148.265 88.255 148.435 ;
        RECT 88.545 148.265 88.715 148.435 ;
        RECT 89.005 148.265 89.175 148.435 ;
        RECT 89.465 148.265 89.635 148.435 ;
        RECT 89.925 148.265 90.095 148.435 ;
        RECT 90.385 148.265 90.555 148.435 ;
        RECT 90.845 148.265 91.015 148.435 ;
        RECT 91.305 148.265 91.475 148.435 ;
        RECT 91.765 148.265 91.935 148.435 ;
        RECT 92.225 148.265 92.395 148.435 ;
        RECT 92.685 148.265 92.855 148.435 ;
        RECT 93.145 148.265 93.315 148.435 ;
        RECT 93.605 148.265 93.775 148.435 ;
        RECT 94.065 148.265 94.235 148.435 ;
        RECT 94.525 148.265 94.695 148.435 ;
        RECT 94.985 148.265 95.155 148.435 ;
        RECT 95.445 148.265 95.615 148.435 ;
        RECT 95.905 148.265 96.075 148.435 ;
        RECT 96.365 148.265 96.535 148.435 ;
        RECT 96.825 148.265 96.995 148.435 ;
        RECT 97.285 148.265 97.455 148.435 ;
        RECT 97.745 148.265 97.915 148.435 ;
        RECT 98.205 148.265 98.375 148.435 ;
        RECT 98.665 148.265 98.835 148.435 ;
        RECT 99.125 148.265 99.295 148.435 ;
        RECT 99.585 148.265 99.755 148.435 ;
        RECT 100.045 148.265 100.215 148.435 ;
        RECT 100.505 148.265 100.675 148.435 ;
        RECT 100.965 148.265 101.135 148.435 ;
        RECT 101.425 148.265 101.595 148.435 ;
        RECT 101.885 148.265 102.055 148.435 ;
        RECT 102.345 148.265 102.515 148.435 ;
        RECT 102.805 148.265 102.975 148.435 ;
        RECT 103.265 148.265 103.435 148.435 ;
        RECT 103.725 148.265 103.895 148.435 ;
        RECT 104.185 148.265 104.355 148.435 ;
        RECT 104.645 148.265 104.815 148.435 ;
        RECT 105.105 148.265 105.275 148.435 ;
        RECT 105.565 148.265 105.735 148.435 ;
        RECT 106.025 148.265 106.195 148.435 ;
        RECT 106.485 148.265 106.655 148.435 ;
        RECT 106.945 148.265 107.115 148.435 ;
        RECT 107.405 148.265 107.575 148.435 ;
        RECT 107.865 148.265 108.035 148.435 ;
        RECT 108.325 148.265 108.495 148.435 ;
        RECT 108.785 148.265 108.955 148.435 ;
        RECT 109.245 148.265 109.415 148.435 ;
        RECT 109.705 148.265 109.875 148.435 ;
        RECT 110.165 148.265 110.335 148.435 ;
        RECT 110.625 148.265 110.795 148.435 ;
        RECT 111.085 148.265 111.255 148.435 ;
        RECT 111.545 148.265 111.715 148.435 ;
        RECT 112.005 148.265 112.175 148.435 ;
        RECT 112.465 148.265 112.635 148.435 ;
        RECT 112.925 148.265 113.095 148.435 ;
        RECT 113.385 148.265 113.555 148.435 ;
        RECT 113.845 148.265 114.015 148.435 ;
        RECT 114.305 148.265 114.475 148.435 ;
        RECT 114.765 148.265 114.935 148.435 ;
        RECT 115.225 148.265 115.395 148.435 ;
        RECT 115.685 148.265 115.855 148.435 ;
        RECT 116.145 148.265 116.315 148.435 ;
        RECT 116.605 148.265 116.775 148.435 ;
        RECT 117.065 148.265 117.235 148.435 ;
        RECT 117.525 148.265 117.695 148.435 ;
        RECT 117.985 148.265 118.155 148.435 ;
        RECT 118.445 148.265 118.615 148.435 ;
        RECT 118.905 148.265 119.075 148.435 ;
        RECT 119.365 148.265 119.535 148.435 ;
        RECT 119.825 148.265 119.995 148.435 ;
        RECT 120.285 148.265 120.455 148.435 ;
        RECT 120.745 148.265 120.915 148.435 ;
        RECT 121.205 148.265 121.375 148.435 ;
        RECT 121.665 148.265 121.835 148.435 ;
        RECT 122.125 148.265 122.295 148.435 ;
        RECT 122.585 148.265 122.755 148.435 ;
        RECT 123.045 148.265 123.215 148.435 ;
        RECT 123.505 148.265 123.675 148.435 ;
        RECT 123.965 148.265 124.135 148.435 ;
        RECT 124.425 148.265 124.595 148.435 ;
        RECT 124.885 148.265 125.055 148.435 ;
        RECT 125.345 148.265 125.515 148.435 ;
        RECT 125.805 148.265 125.975 148.435 ;
        RECT 126.265 148.265 126.435 148.435 ;
        RECT 126.725 148.265 126.895 148.435 ;
        RECT 127.185 148.265 127.355 148.435 ;
        RECT 127.645 148.265 127.815 148.435 ;
        RECT 128.105 148.265 128.275 148.435 ;
        RECT 128.565 148.265 128.735 148.435 ;
        RECT 129.025 148.265 129.195 148.435 ;
        RECT 129.485 148.265 129.655 148.435 ;
        RECT 129.945 148.265 130.115 148.435 ;
        RECT 130.405 148.265 130.575 148.435 ;
        RECT 130.865 148.265 131.035 148.435 ;
        RECT 131.325 148.265 131.495 148.435 ;
        RECT 131.785 148.265 131.955 148.435 ;
        RECT 132.245 148.265 132.415 148.435 ;
        RECT 132.705 148.265 132.875 148.435 ;
        RECT 133.165 148.265 133.335 148.435 ;
        RECT 133.625 148.265 133.795 148.435 ;
        RECT 134.085 148.265 134.255 148.435 ;
        RECT 134.545 148.265 134.715 148.435 ;
        RECT 135.005 148.265 135.175 148.435 ;
        RECT 135.465 148.265 135.635 148.435 ;
        RECT 135.925 148.265 136.095 148.435 ;
        RECT 136.385 148.265 136.555 148.435 ;
        RECT 136.845 148.265 137.015 148.435 ;
        RECT 137.305 148.265 137.475 148.435 ;
        RECT 137.765 148.265 137.935 148.435 ;
        RECT 138.225 148.265 138.395 148.435 ;
        RECT 138.685 148.265 138.855 148.435 ;
        RECT 139.145 148.265 139.315 148.435 ;
        RECT 139.605 148.265 139.775 148.435 ;
        RECT 140.065 148.265 140.235 148.435 ;
        RECT 140.525 148.265 140.695 148.435 ;
        RECT 140.985 148.265 141.155 148.435 ;
        RECT 141.445 148.265 141.615 148.435 ;
        RECT 141.905 148.265 142.075 148.435 ;
        RECT 142.365 148.265 142.535 148.435 ;
        RECT 142.825 148.265 142.995 148.435 ;
        RECT 143.285 148.265 143.455 148.435 ;
        RECT 143.745 148.265 143.915 148.435 ;
        RECT 144.205 148.265 144.375 148.435 ;
        RECT 144.665 148.265 144.835 148.435 ;
        RECT 145.125 148.265 145.295 148.435 ;
        RECT 145.585 148.265 145.755 148.435 ;
        RECT 146.045 148.265 146.215 148.435 ;
        RECT 146.505 148.265 146.675 148.435 ;
        RECT 146.965 148.265 147.135 148.435 ;
        RECT 147.425 148.265 147.595 148.435 ;
        RECT 147.885 148.265 148.055 148.435 ;
        RECT 148.345 148.265 148.515 148.435 ;
        RECT 148.805 148.265 148.975 148.435 ;
        RECT 149.265 148.265 149.435 148.435 ;
        RECT 149.725 148.265 149.895 148.435 ;
        RECT 150.185 148.265 150.355 148.435 ;
        RECT 18.625 147.075 18.795 147.245 ;
        RECT 20.465 147.415 20.635 147.585 ;
        RECT 21.385 146.735 21.555 146.905 ;
        RECT 23.225 147.415 23.395 147.585 ;
        RECT 23.685 147.415 23.855 147.585 ;
        RECT 24.605 146.735 24.775 146.905 ;
        RECT 25.525 146.735 25.695 146.905 ;
        RECT 25.065 146.395 25.235 146.565 ;
        RECT 26.445 147.075 26.615 147.245 ;
        RECT 26.905 146.735 27.075 146.905 ;
        RECT 27.365 146.735 27.535 146.905 ;
        RECT 27.825 146.735 27.995 146.905 ;
        RECT 28.745 146.055 28.915 146.225 ;
        RECT 29.205 147.075 29.375 147.245 ;
        RECT 30.125 146.735 30.295 146.905 ;
        RECT 38.430 147.415 38.600 147.585 ;
        RECT 31.505 146.735 31.675 146.905 ;
        RECT 32.425 146.735 32.595 146.905 ;
        RECT 37.945 146.735 38.115 146.905 ;
        RECT 38.825 147.075 38.995 147.245 ;
        RECT 39.280 146.395 39.450 146.565 ;
        RECT 40.530 147.415 40.700 147.585 ;
        RECT 40.015 147.075 40.185 147.245 ;
        RECT 42.100 147.415 42.270 147.585 ;
        RECT 42.535 147.075 42.705 147.245 ;
        RECT 44.845 147.415 45.015 147.585 ;
        RECT 45.765 147.755 45.935 147.925 ;
        RECT 46.685 146.395 46.855 146.565 ;
        RECT 47.605 146.735 47.775 146.905 ;
        RECT 48.065 146.735 48.235 146.905 ;
        RECT 51.745 147.755 51.915 147.925 ;
        RECT 52.665 147.755 52.835 147.925 ;
        RECT 50.825 146.735 50.995 146.905 ;
        RECT 48.985 146.055 49.155 146.225 ;
        RECT 51.745 146.735 51.915 146.905 ;
        RECT 54.505 147.415 54.675 147.585 ;
        RECT 52.205 146.735 52.375 146.905 ;
        RECT 53.585 146.735 53.755 146.905 ;
        RECT 57.265 147.075 57.435 147.245 ;
        RECT 56.805 146.735 56.975 146.905 ;
        RECT 58.645 147.075 58.815 147.245 ;
        RECT 60.945 147.415 61.115 147.585 ;
        RECT 59.565 146.735 59.735 146.905 ;
        RECT 60.025 146.055 60.195 146.225 ;
        RECT 60.945 146.395 61.115 146.565 ;
        RECT 62.325 147.075 62.495 147.245 ;
        RECT 62.785 146.735 62.955 146.905 ;
        RECT 61.405 146.055 61.575 146.225 ;
        RECT 64.165 146.735 64.335 146.905 ;
        RECT 64.625 147.075 64.795 147.245 ;
        RECT 68.765 147.755 68.935 147.925 ;
        RECT 66.010 146.735 66.180 146.905 ;
        RECT 66.465 147.075 66.635 147.245 ;
        RECT 66.925 146.735 67.095 146.905 ;
        RECT 67.385 147.075 67.555 147.245 ;
        RECT 65.085 146.055 65.255 146.225 ;
        RECT 69.645 146.785 69.815 146.955 ;
        RECT 70.145 146.735 70.315 146.905 ;
        RECT 71.065 146.735 71.235 146.905 ;
        RECT 71.525 146.735 71.695 146.905 ;
        RECT 77.505 146.395 77.675 146.565 ;
        RECT 79.805 147.075 79.975 147.245 ;
        RECT 81.185 146.735 81.355 146.905 ;
        RECT 81.645 146.735 81.815 146.905 ;
        RECT 82.105 146.735 82.275 146.905 ;
        RECT 77.965 146.055 78.135 146.225 ;
        RECT 83.025 146.735 83.195 146.905 ;
        RECT 86.245 147.075 86.415 147.245 ;
        RECT 86.705 146.735 86.875 146.905 ;
        RECT 88.545 147.415 88.715 147.585 ;
        RECT 99.585 146.735 99.755 146.905 ;
        RECT 104.205 147.755 104.375 147.925 ;
        RECT 105.125 147.755 105.295 147.925 ;
        RECT 100.045 146.055 100.215 146.225 ;
        RECT 102.805 147.075 102.975 147.245 ;
        RECT 103.265 146.735 103.435 146.905 ;
        RECT 107.405 147.075 107.575 147.245 ;
        RECT 108.325 147.755 108.495 147.925 ;
        RECT 107.865 146.735 108.035 146.905 ;
        RECT 108.785 146.735 108.955 146.905 ;
        RECT 111.085 147.075 111.255 147.245 ;
        RECT 110.625 146.735 110.795 146.905 ;
        RECT 116.145 147.415 116.315 147.585 ;
        RECT 113.385 146.735 113.555 146.905 ;
        RECT 114.305 146.735 114.475 146.905 ;
        RECT 112.465 146.055 112.635 146.225 ;
        RECT 115.225 146.735 115.395 146.905 ;
        RECT 114.765 146.395 114.935 146.565 ;
        RECT 116.605 147.755 116.775 147.925 ;
        RECT 117.525 146.735 117.695 146.905 ;
        RECT 117.985 146.735 118.155 146.905 ;
        RECT 11.265 145.545 11.435 145.715 ;
        RECT 11.725 145.545 11.895 145.715 ;
        RECT 12.185 145.545 12.355 145.715 ;
        RECT 12.645 145.545 12.815 145.715 ;
        RECT 13.105 145.545 13.275 145.715 ;
        RECT 13.565 145.545 13.735 145.715 ;
        RECT 14.025 145.545 14.195 145.715 ;
        RECT 14.485 145.545 14.655 145.715 ;
        RECT 14.945 145.545 15.115 145.715 ;
        RECT 15.405 145.545 15.575 145.715 ;
        RECT 15.865 145.545 16.035 145.715 ;
        RECT 16.325 145.545 16.495 145.715 ;
        RECT 16.785 145.545 16.955 145.715 ;
        RECT 17.245 145.545 17.415 145.715 ;
        RECT 17.705 145.545 17.875 145.715 ;
        RECT 18.165 145.545 18.335 145.715 ;
        RECT 18.625 145.545 18.795 145.715 ;
        RECT 19.085 145.545 19.255 145.715 ;
        RECT 19.545 145.545 19.715 145.715 ;
        RECT 20.005 145.545 20.175 145.715 ;
        RECT 20.465 145.545 20.635 145.715 ;
        RECT 20.925 145.545 21.095 145.715 ;
        RECT 21.385 145.545 21.555 145.715 ;
        RECT 21.845 145.545 22.015 145.715 ;
        RECT 22.305 145.545 22.475 145.715 ;
        RECT 22.765 145.545 22.935 145.715 ;
        RECT 23.225 145.545 23.395 145.715 ;
        RECT 23.685 145.545 23.855 145.715 ;
        RECT 24.145 145.545 24.315 145.715 ;
        RECT 24.605 145.545 24.775 145.715 ;
        RECT 25.065 145.545 25.235 145.715 ;
        RECT 25.525 145.545 25.695 145.715 ;
        RECT 25.985 145.545 26.155 145.715 ;
        RECT 26.445 145.545 26.615 145.715 ;
        RECT 26.905 145.545 27.075 145.715 ;
        RECT 27.365 145.545 27.535 145.715 ;
        RECT 27.825 145.545 27.995 145.715 ;
        RECT 28.285 145.545 28.455 145.715 ;
        RECT 28.745 145.545 28.915 145.715 ;
        RECT 29.205 145.545 29.375 145.715 ;
        RECT 29.665 145.545 29.835 145.715 ;
        RECT 30.125 145.545 30.295 145.715 ;
        RECT 30.585 145.545 30.755 145.715 ;
        RECT 31.045 145.545 31.215 145.715 ;
        RECT 31.505 145.545 31.675 145.715 ;
        RECT 31.965 145.545 32.135 145.715 ;
        RECT 32.425 145.545 32.595 145.715 ;
        RECT 32.885 145.545 33.055 145.715 ;
        RECT 33.345 145.545 33.515 145.715 ;
        RECT 33.805 145.545 33.975 145.715 ;
        RECT 34.265 145.545 34.435 145.715 ;
        RECT 34.725 145.545 34.895 145.715 ;
        RECT 35.185 145.545 35.355 145.715 ;
        RECT 35.645 145.545 35.815 145.715 ;
        RECT 36.105 145.545 36.275 145.715 ;
        RECT 36.565 145.545 36.735 145.715 ;
        RECT 37.025 145.545 37.195 145.715 ;
        RECT 37.485 145.545 37.655 145.715 ;
        RECT 37.945 145.545 38.115 145.715 ;
        RECT 38.405 145.545 38.575 145.715 ;
        RECT 38.865 145.545 39.035 145.715 ;
        RECT 39.325 145.545 39.495 145.715 ;
        RECT 39.785 145.545 39.955 145.715 ;
        RECT 40.245 145.545 40.415 145.715 ;
        RECT 40.705 145.545 40.875 145.715 ;
        RECT 41.165 145.545 41.335 145.715 ;
        RECT 41.625 145.545 41.795 145.715 ;
        RECT 42.085 145.545 42.255 145.715 ;
        RECT 42.545 145.545 42.715 145.715 ;
        RECT 43.005 145.545 43.175 145.715 ;
        RECT 43.465 145.545 43.635 145.715 ;
        RECT 43.925 145.545 44.095 145.715 ;
        RECT 44.385 145.545 44.555 145.715 ;
        RECT 44.845 145.545 45.015 145.715 ;
        RECT 45.305 145.545 45.475 145.715 ;
        RECT 45.765 145.545 45.935 145.715 ;
        RECT 46.225 145.545 46.395 145.715 ;
        RECT 46.685 145.545 46.855 145.715 ;
        RECT 47.145 145.545 47.315 145.715 ;
        RECT 47.605 145.545 47.775 145.715 ;
        RECT 48.065 145.545 48.235 145.715 ;
        RECT 48.525 145.545 48.695 145.715 ;
        RECT 48.985 145.545 49.155 145.715 ;
        RECT 49.445 145.545 49.615 145.715 ;
        RECT 49.905 145.545 50.075 145.715 ;
        RECT 50.365 145.545 50.535 145.715 ;
        RECT 50.825 145.545 50.995 145.715 ;
        RECT 51.285 145.545 51.455 145.715 ;
        RECT 51.745 145.545 51.915 145.715 ;
        RECT 52.205 145.545 52.375 145.715 ;
        RECT 52.665 145.545 52.835 145.715 ;
        RECT 53.125 145.545 53.295 145.715 ;
        RECT 53.585 145.545 53.755 145.715 ;
        RECT 54.045 145.545 54.215 145.715 ;
        RECT 54.505 145.545 54.675 145.715 ;
        RECT 54.965 145.545 55.135 145.715 ;
        RECT 55.425 145.545 55.595 145.715 ;
        RECT 55.885 145.545 56.055 145.715 ;
        RECT 56.345 145.545 56.515 145.715 ;
        RECT 56.805 145.545 56.975 145.715 ;
        RECT 57.265 145.545 57.435 145.715 ;
        RECT 57.725 145.545 57.895 145.715 ;
        RECT 58.185 145.545 58.355 145.715 ;
        RECT 58.645 145.545 58.815 145.715 ;
        RECT 59.105 145.545 59.275 145.715 ;
        RECT 59.565 145.545 59.735 145.715 ;
        RECT 60.025 145.545 60.195 145.715 ;
        RECT 60.485 145.545 60.655 145.715 ;
        RECT 60.945 145.545 61.115 145.715 ;
        RECT 61.405 145.545 61.575 145.715 ;
        RECT 61.865 145.545 62.035 145.715 ;
        RECT 62.325 145.545 62.495 145.715 ;
        RECT 62.785 145.545 62.955 145.715 ;
        RECT 63.245 145.545 63.415 145.715 ;
        RECT 63.705 145.545 63.875 145.715 ;
        RECT 64.165 145.545 64.335 145.715 ;
        RECT 64.625 145.545 64.795 145.715 ;
        RECT 65.085 145.545 65.255 145.715 ;
        RECT 65.545 145.545 65.715 145.715 ;
        RECT 66.005 145.545 66.175 145.715 ;
        RECT 66.465 145.545 66.635 145.715 ;
        RECT 66.925 145.545 67.095 145.715 ;
        RECT 67.385 145.545 67.555 145.715 ;
        RECT 67.845 145.545 68.015 145.715 ;
        RECT 68.305 145.545 68.475 145.715 ;
        RECT 68.765 145.545 68.935 145.715 ;
        RECT 69.225 145.545 69.395 145.715 ;
        RECT 69.685 145.545 69.855 145.715 ;
        RECT 70.145 145.545 70.315 145.715 ;
        RECT 70.605 145.545 70.775 145.715 ;
        RECT 71.065 145.545 71.235 145.715 ;
        RECT 71.525 145.545 71.695 145.715 ;
        RECT 71.985 145.545 72.155 145.715 ;
        RECT 72.445 145.545 72.615 145.715 ;
        RECT 72.905 145.545 73.075 145.715 ;
        RECT 73.365 145.545 73.535 145.715 ;
        RECT 73.825 145.545 73.995 145.715 ;
        RECT 74.285 145.545 74.455 145.715 ;
        RECT 74.745 145.545 74.915 145.715 ;
        RECT 75.205 145.545 75.375 145.715 ;
        RECT 75.665 145.545 75.835 145.715 ;
        RECT 76.125 145.545 76.295 145.715 ;
        RECT 76.585 145.545 76.755 145.715 ;
        RECT 77.045 145.545 77.215 145.715 ;
        RECT 77.505 145.545 77.675 145.715 ;
        RECT 77.965 145.545 78.135 145.715 ;
        RECT 78.425 145.545 78.595 145.715 ;
        RECT 78.885 145.545 79.055 145.715 ;
        RECT 79.345 145.545 79.515 145.715 ;
        RECT 79.805 145.545 79.975 145.715 ;
        RECT 80.265 145.545 80.435 145.715 ;
        RECT 80.725 145.545 80.895 145.715 ;
        RECT 81.185 145.545 81.355 145.715 ;
        RECT 81.645 145.545 81.815 145.715 ;
        RECT 82.105 145.545 82.275 145.715 ;
        RECT 82.565 145.545 82.735 145.715 ;
        RECT 83.025 145.545 83.195 145.715 ;
        RECT 83.485 145.545 83.655 145.715 ;
        RECT 83.945 145.545 84.115 145.715 ;
        RECT 84.405 145.545 84.575 145.715 ;
        RECT 84.865 145.545 85.035 145.715 ;
        RECT 85.325 145.545 85.495 145.715 ;
        RECT 85.785 145.545 85.955 145.715 ;
        RECT 86.245 145.545 86.415 145.715 ;
        RECT 86.705 145.545 86.875 145.715 ;
        RECT 87.165 145.545 87.335 145.715 ;
        RECT 87.625 145.545 87.795 145.715 ;
        RECT 88.085 145.545 88.255 145.715 ;
        RECT 88.545 145.545 88.715 145.715 ;
        RECT 89.005 145.545 89.175 145.715 ;
        RECT 89.465 145.545 89.635 145.715 ;
        RECT 89.925 145.545 90.095 145.715 ;
        RECT 90.385 145.545 90.555 145.715 ;
        RECT 90.845 145.545 91.015 145.715 ;
        RECT 91.305 145.545 91.475 145.715 ;
        RECT 91.765 145.545 91.935 145.715 ;
        RECT 92.225 145.545 92.395 145.715 ;
        RECT 92.685 145.545 92.855 145.715 ;
        RECT 93.145 145.545 93.315 145.715 ;
        RECT 93.605 145.545 93.775 145.715 ;
        RECT 94.065 145.545 94.235 145.715 ;
        RECT 94.525 145.545 94.695 145.715 ;
        RECT 94.985 145.545 95.155 145.715 ;
        RECT 95.445 145.545 95.615 145.715 ;
        RECT 95.905 145.545 96.075 145.715 ;
        RECT 96.365 145.545 96.535 145.715 ;
        RECT 96.825 145.545 96.995 145.715 ;
        RECT 97.285 145.545 97.455 145.715 ;
        RECT 97.745 145.545 97.915 145.715 ;
        RECT 98.205 145.545 98.375 145.715 ;
        RECT 98.665 145.545 98.835 145.715 ;
        RECT 99.125 145.545 99.295 145.715 ;
        RECT 99.585 145.545 99.755 145.715 ;
        RECT 100.045 145.545 100.215 145.715 ;
        RECT 100.505 145.545 100.675 145.715 ;
        RECT 100.965 145.545 101.135 145.715 ;
        RECT 101.425 145.545 101.595 145.715 ;
        RECT 101.885 145.545 102.055 145.715 ;
        RECT 102.345 145.545 102.515 145.715 ;
        RECT 102.805 145.545 102.975 145.715 ;
        RECT 103.265 145.545 103.435 145.715 ;
        RECT 103.725 145.545 103.895 145.715 ;
        RECT 104.185 145.545 104.355 145.715 ;
        RECT 104.645 145.545 104.815 145.715 ;
        RECT 105.105 145.545 105.275 145.715 ;
        RECT 105.565 145.545 105.735 145.715 ;
        RECT 106.025 145.545 106.195 145.715 ;
        RECT 106.485 145.545 106.655 145.715 ;
        RECT 106.945 145.545 107.115 145.715 ;
        RECT 107.405 145.545 107.575 145.715 ;
        RECT 107.865 145.545 108.035 145.715 ;
        RECT 108.325 145.545 108.495 145.715 ;
        RECT 108.785 145.545 108.955 145.715 ;
        RECT 109.245 145.545 109.415 145.715 ;
        RECT 109.705 145.545 109.875 145.715 ;
        RECT 110.165 145.545 110.335 145.715 ;
        RECT 110.625 145.545 110.795 145.715 ;
        RECT 111.085 145.545 111.255 145.715 ;
        RECT 111.545 145.545 111.715 145.715 ;
        RECT 112.005 145.545 112.175 145.715 ;
        RECT 112.465 145.545 112.635 145.715 ;
        RECT 112.925 145.545 113.095 145.715 ;
        RECT 113.385 145.545 113.555 145.715 ;
        RECT 113.845 145.545 114.015 145.715 ;
        RECT 114.305 145.545 114.475 145.715 ;
        RECT 114.765 145.545 114.935 145.715 ;
        RECT 115.225 145.545 115.395 145.715 ;
        RECT 115.685 145.545 115.855 145.715 ;
        RECT 116.145 145.545 116.315 145.715 ;
        RECT 116.605 145.545 116.775 145.715 ;
        RECT 117.065 145.545 117.235 145.715 ;
        RECT 117.525 145.545 117.695 145.715 ;
        RECT 117.985 145.545 118.155 145.715 ;
        RECT 118.445 145.545 118.615 145.715 ;
        RECT 118.905 145.545 119.075 145.715 ;
        RECT 119.365 145.545 119.535 145.715 ;
        RECT 119.825 145.545 119.995 145.715 ;
        RECT 120.285 145.545 120.455 145.715 ;
        RECT 120.745 145.545 120.915 145.715 ;
        RECT 121.205 145.545 121.375 145.715 ;
        RECT 121.665 145.545 121.835 145.715 ;
        RECT 122.125 145.545 122.295 145.715 ;
        RECT 122.585 145.545 122.755 145.715 ;
        RECT 123.045 145.545 123.215 145.715 ;
        RECT 123.505 145.545 123.675 145.715 ;
        RECT 123.965 145.545 124.135 145.715 ;
        RECT 124.425 145.545 124.595 145.715 ;
        RECT 124.885 145.545 125.055 145.715 ;
        RECT 125.345 145.545 125.515 145.715 ;
        RECT 125.805 145.545 125.975 145.715 ;
        RECT 126.265 145.545 126.435 145.715 ;
        RECT 126.725 145.545 126.895 145.715 ;
        RECT 127.185 145.545 127.355 145.715 ;
        RECT 127.645 145.545 127.815 145.715 ;
        RECT 128.105 145.545 128.275 145.715 ;
        RECT 128.565 145.545 128.735 145.715 ;
        RECT 129.025 145.545 129.195 145.715 ;
        RECT 129.485 145.545 129.655 145.715 ;
        RECT 129.945 145.545 130.115 145.715 ;
        RECT 130.405 145.545 130.575 145.715 ;
        RECT 130.865 145.545 131.035 145.715 ;
        RECT 131.325 145.545 131.495 145.715 ;
        RECT 131.785 145.545 131.955 145.715 ;
        RECT 132.245 145.545 132.415 145.715 ;
        RECT 132.705 145.545 132.875 145.715 ;
        RECT 133.165 145.545 133.335 145.715 ;
        RECT 133.625 145.545 133.795 145.715 ;
        RECT 134.085 145.545 134.255 145.715 ;
        RECT 134.545 145.545 134.715 145.715 ;
        RECT 135.005 145.545 135.175 145.715 ;
        RECT 135.465 145.545 135.635 145.715 ;
        RECT 135.925 145.545 136.095 145.715 ;
        RECT 136.385 145.545 136.555 145.715 ;
        RECT 136.845 145.545 137.015 145.715 ;
        RECT 137.305 145.545 137.475 145.715 ;
        RECT 137.765 145.545 137.935 145.715 ;
        RECT 138.225 145.545 138.395 145.715 ;
        RECT 138.685 145.545 138.855 145.715 ;
        RECT 139.145 145.545 139.315 145.715 ;
        RECT 139.605 145.545 139.775 145.715 ;
        RECT 140.065 145.545 140.235 145.715 ;
        RECT 140.525 145.545 140.695 145.715 ;
        RECT 140.985 145.545 141.155 145.715 ;
        RECT 141.445 145.545 141.615 145.715 ;
        RECT 141.905 145.545 142.075 145.715 ;
        RECT 142.365 145.545 142.535 145.715 ;
        RECT 142.825 145.545 142.995 145.715 ;
        RECT 143.285 145.545 143.455 145.715 ;
        RECT 143.745 145.545 143.915 145.715 ;
        RECT 144.205 145.545 144.375 145.715 ;
        RECT 144.665 145.545 144.835 145.715 ;
        RECT 145.125 145.545 145.295 145.715 ;
        RECT 145.585 145.545 145.755 145.715 ;
        RECT 146.045 145.545 146.215 145.715 ;
        RECT 146.505 145.545 146.675 145.715 ;
        RECT 146.965 145.545 147.135 145.715 ;
        RECT 147.425 145.545 147.595 145.715 ;
        RECT 147.885 145.545 148.055 145.715 ;
        RECT 148.345 145.545 148.515 145.715 ;
        RECT 148.805 145.545 148.975 145.715 ;
        RECT 149.265 145.545 149.435 145.715 ;
        RECT 149.725 145.545 149.895 145.715 ;
        RECT 150.185 145.545 150.355 145.715 ;
        RECT 24.145 144.355 24.315 144.525 ;
        RECT 25.065 144.355 25.235 144.525 ;
        RECT 25.525 144.355 25.695 144.525 ;
        RECT 24.145 143.675 24.315 143.845 ;
        RECT 27.365 144.355 27.535 144.525 ;
        RECT 26.905 144.015 27.075 144.185 ;
        RECT 29.205 144.015 29.375 144.185 ;
        RECT 38.405 144.355 38.575 144.525 ;
        RECT 39.325 144.355 39.495 144.525 ;
        RECT 37.485 144.015 37.655 144.185 ;
        RECT 39.785 145.035 39.955 145.205 ;
        RECT 40.705 144.355 40.875 144.525 ;
        RECT 50.825 144.355 50.995 144.525 ;
        RECT 51.745 144.355 51.915 144.525 ;
        RECT 51.745 143.675 51.915 143.845 ;
        RECT 53.125 144.015 53.295 144.185 ;
        RECT 61.420 144.355 61.590 144.525 ;
        RECT 60.485 144.015 60.655 144.185 ;
        RECT 62.325 143.335 62.495 143.505 ;
        RECT 63.705 144.015 63.875 144.185 ;
        RECT 64.190 143.675 64.360 143.845 ;
        RECT 64.585 144.015 64.755 144.185 ;
        RECT 65.040 144.355 65.210 144.525 ;
        RECT 65.775 144.015 65.945 144.185 ;
        RECT 66.290 143.675 66.460 143.845 ;
        RECT 67.860 143.675 68.030 143.845 ;
        RECT 68.295 144.015 68.465 144.185 ;
        RECT 70.605 145.035 70.775 145.205 ;
        RECT 71.065 144.015 71.235 144.185 ;
        RECT 71.550 143.675 71.720 143.845 ;
        RECT 71.945 144.015 72.115 144.185 ;
        RECT 72.400 144.695 72.570 144.865 ;
        RECT 73.135 144.015 73.305 144.185 ;
        RECT 73.650 143.675 73.820 143.845 ;
        RECT 75.220 143.675 75.390 143.845 ;
        RECT 75.655 144.015 75.825 144.185 ;
        RECT 77.965 145.035 78.135 145.205 ;
        RECT 79.805 145.035 79.975 145.205 ;
        RECT 78.425 144.015 78.595 144.185 ;
        RECT 79.805 144.355 79.975 144.525 ;
        RECT 79.345 143.675 79.515 143.845 ;
        RECT 82.105 144.355 82.275 144.525 ;
        RECT 83.025 144.355 83.195 144.525 ;
        RECT 83.945 144.695 84.115 144.865 ;
        RECT 86.245 145.035 86.415 145.205 ;
        RECT 87.005 144.695 87.175 144.865 ;
        RECT 88.085 144.695 88.255 144.865 ;
        RECT 89.005 145.035 89.175 145.205 ;
        RECT 87.165 143.335 87.335 143.505 ;
        RECT 89.925 144.355 90.095 144.525 ;
        RECT 90.845 144.355 91.015 144.525 ;
        RECT 94.985 145.035 95.155 145.205 ;
        RECT 93.145 144.355 93.315 144.525 ;
        RECT 92.685 144.015 92.855 144.185 ;
        RECT 102.805 144.695 102.975 144.865 ;
        RECT 104.185 143.675 104.355 143.845 ;
        RECT 105.105 143.335 105.275 143.505 ;
        RECT 115.685 144.355 115.855 144.525 ;
        RECT 116.605 143.335 116.775 143.505 ;
        RECT 11.265 142.825 11.435 142.995 ;
        RECT 11.725 142.825 11.895 142.995 ;
        RECT 12.185 142.825 12.355 142.995 ;
        RECT 12.645 142.825 12.815 142.995 ;
        RECT 13.105 142.825 13.275 142.995 ;
        RECT 13.565 142.825 13.735 142.995 ;
        RECT 14.025 142.825 14.195 142.995 ;
        RECT 14.485 142.825 14.655 142.995 ;
        RECT 14.945 142.825 15.115 142.995 ;
        RECT 15.405 142.825 15.575 142.995 ;
        RECT 15.865 142.825 16.035 142.995 ;
        RECT 16.325 142.825 16.495 142.995 ;
        RECT 16.785 142.825 16.955 142.995 ;
        RECT 17.245 142.825 17.415 142.995 ;
        RECT 17.705 142.825 17.875 142.995 ;
        RECT 18.165 142.825 18.335 142.995 ;
        RECT 18.625 142.825 18.795 142.995 ;
        RECT 19.085 142.825 19.255 142.995 ;
        RECT 19.545 142.825 19.715 142.995 ;
        RECT 20.005 142.825 20.175 142.995 ;
        RECT 20.465 142.825 20.635 142.995 ;
        RECT 20.925 142.825 21.095 142.995 ;
        RECT 21.385 142.825 21.555 142.995 ;
        RECT 21.845 142.825 22.015 142.995 ;
        RECT 22.305 142.825 22.475 142.995 ;
        RECT 22.765 142.825 22.935 142.995 ;
        RECT 23.225 142.825 23.395 142.995 ;
        RECT 23.685 142.825 23.855 142.995 ;
        RECT 24.145 142.825 24.315 142.995 ;
        RECT 24.605 142.825 24.775 142.995 ;
        RECT 25.065 142.825 25.235 142.995 ;
        RECT 25.525 142.825 25.695 142.995 ;
        RECT 25.985 142.825 26.155 142.995 ;
        RECT 26.445 142.825 26.615 142.995 ;
        RECT 26.905 142.825 27.075 142.995 ;
        RECT 27.365 142.825 27.535 142.995 ;
        RECT 27.825 142.825 27.995 142.995 ;
        RECT 28.285 142.825 28.455 142.995 ;
        RECT 28.745 142.825 28.915 142.995 ;
        RECT 29.205 142.825 29.375 142.995 ;
        RECT 29.665 142.825 29.835 142.995 ;
        RECT 30.125 142.825 30.295 142.995 ;
        RECT 30.585 142.825 30.755 142.995 ;
        RECT 31.045 142.825 31.215 142.995 ;
        RECT 31.505 142.825 31.675 142.995 ;
        RECT 31.965 142.825 32.135 142.995 ;
        RECT 32.425 142.825 32.595 142.995 ;
        RECT 32.885 142.825 33.055 142.995 ;
        RECT 33.345 142.825 33.515 142.995 ;
        RECT 33.805 142.825 33.975 142.995 ;
        RECT 34.265 142.825 34.435 142.995 ;
        RECT 34.725 142.825 34.895 142.995 ;
        RECT 35.185 142.825 35.355 142.995 ;
        RECT 35.645 142.825 35.815 142.995 ;
        RECT 36.105 142.825 36.275 142.995 ;
        RECT 36.565 142.825 36.735 142.995 ;
        RECT 37.025 142.825 37.195 142.995 ;
        RECT 37.485 142.825 37.655 142.995 ;
        RECT 37.945 142.825 38.115 142.995 ;
        RECT 38.405 142.825 38.575 142.995 ;
        RECT 38.865 142.825 39.035 142.995 ;
        RECT 39.325 142.825 39.495 142.995 ;
        RECT 39.785 142.825 39.955 142.995 ;
        RECT 40.245 142.825 40.415 142.995 ;
        RECT 40.705 142.825 40.875 142.995 ;
        RECT 41.165 142.825 41.335 142.995 ;
        RECT 41.625 142.825 41.795 142.995 ;
        RECT 42.085 142.825 42.255 142.995 ;
        RECT 42.545 142.825 42.715 142.995 ;
        RECT 43.005 142.825 43.175 142.995 ;
        RECT 43.465 142.825 43.635 142.995 ;
        RECT 43.925 142.825 44.095 142.995 ;
        RECT 44.385 142.825 44.555 142.995 ;
        RECT 44.845 142.825 45.015 142.995 ;
        RECT 45.305 142.825 45.475 142.995 ;
        RECT 45.765 142.825 45.935 142.995 ;
        RECT 46.225 142.825 46.395 142.995 ;
        RECT 46.685 142.825 46.855 142.995 ;
        RECT 47.145 142.825 47.315 142.995 ;
        RECT 47.605 142.825 47.775 142.995 ;
        RECT 48.065 142.825 48.235 142.995 ;
        RECT 48.525 142.825 48.695 142.995 ;
        RECT 48.985 142.825 49.155 142.995 ;
        RECT 49.445 142.825 49.615 142.995 ;
        RECT 49.905 142.825 50.075 142.995 ;
        RECT 50.365 142.825 50.535 142.995 ;
        RECT 50.825 142.825 50.995 142.995 ;
        RECT 51.285 142.825 51.455 142.995 ;
        RECT 51.745 142.825 51.915 142.995 ;
        RECT 52.205 142.825 52.375 142.995 ;
        RECT 52.665 142.825 52.835 142.995 ;
        RECT 53.125 142.825 53.295 142.995 ;
        RECT 53.585 142.825 53.755 142.995 ;
        RECT 54.045 142.825 54.215 142.995 ;
        RECT 54.505 142.825 54.675 142.995 ;
        RECT 54.965 142.825 55.135 142.995 ;
        RECT 55.425 142.825 55.595 142.995 ;
        RECT 55.885 142.825 56.055 142.995 ;
        RECT 56.345 142.825 56.515 142.995 ;
        RECT 56.805 142.825 56.975 142.995 ;
        RECT 57.265 142.825 57.435 142.995 ;
        RECT 57.725 142.825 57.895 142.995 ;
        RECT 58.185 142.825 58.355 142.995 ;
        RECT 58.645 142.825 58.815 142.995 ;
        RECT 59.105 142.825 59.275 142.995 ;
        RECT 59.565 142.825 59.735 142.995 ;
        RECT 60.025 142.825 60.195 142.995 ;
        RECT 60.485 142.825 60.655 142.995 ;
        RECT 60.945 142.825 61.115 142.995 ;
        RECT 61.405 142.825 61.575 142.995 ;
        RECT 61.865 142.825 62.035 142.995 ;
        RECT 62.325 142.825 62.495 142.995 ;
        RECT 62.785 142.825 62.955 142.995 ;
        RECT 63.245 142.825 63.415 142.995 ;
        RECT 63.705 142.825 63.875 142.995 ;
        RECT 64.165 142.825 64.335 142.995 ;
        RECT 64.625 142.825 64.795 142.995 ;
        RECT 65.085 142.825 65.255 142.995 ;
        RECT 65.545 142.825 65.715 142.995 ;
        RECT 66.005 142.825 66.175 142.995 ;
        RECT 66.465 142.825 66.635 142.995 ;
        RECT 66.925 142.825 67.095 142.995 ;
        RECT 67.385 142.825 67.555 142.995 ;
        RECT 67.845 142.825 68.015 142.995 ;
        RECT 68.305 142.825 68.475 142.995 ;
        RECT 68.765 142.825 68.935 142.995 ;
        RECT 69.225 142.825 69.395 142.995 ;
        RECT 69.685 142.825 69.855 142.995 ;
        RECT 70.145 142.825 70.315 142.995 ;
        RECT 70.605 142.825 70.775 142.995 ;
        RECT 71.065 142.825 71.235 142.995 ;
        RECT 71.525 142.825 71.695 142.995 ;
        RECT 71.985 142.825 72.155 142.995 ;
        RECT 72.445 142.825 72.615 142.995 ;
        RECT 72.905 142.825 73.075 142.995 ;
        RECT 73.365 142.825 73.535 142.995 ;
        RECT 73.825 142.825 73.995 142.995 ;
        RECT 74.285 142.825 74.455 142.995 ;
        RECT 74.745 142.825 74.915 142.995 ;
        RECT 75.205 142.825 75.375 142.995 ;
        RECT 75.665 142.825 75.835 142.995 ;
        RECT 76.125 142.825 76.295 142.995 ;
        RECT 76.585 142.825 76.755 142.995 ;
        RECT 77.045 142.825 77.215 142.995 ;
        RECT 77.505 142.825 77.675 142.995 ;
        RECT 77.965 142.825 78.135 142.995 ;
        RECT 78.425 142.825 78.595 142.995 ;
        RECT 78.885 142.825 79.055 142.995 ;
        RECT 79.345 142.825 79.515 142.995 ;
        RECT 79.805 142.825 79.975 142.995 ;
        RECT 80.265 142.825 80.435 142.995 ;
        RECT 80.725 142.825 80.895 142.995 ;
        RECT 81.185 142.825 81.355 142.995 ;
        RECT 81.645 142.825 81.815 142.995 ;
        RECT 82.105 142.825 82.275 142.995 ;
        RECT 82.565 142.825 82.735 142.995 ;
        RECT 83.025 142.825 83.195 142.995 ;
        RECT 83.485 142.825 83.655 142.995 ;
        RECT 83.945 142.825 84.115 142.995 ;
        RECT 84.405 142.825 84.575 142.995 ;
        RECT 84.865 142.825 85.035 142.995 ;
        RECT 85.325 142.825 85.495 142.995 ;
        RECT 85.785 142.825 85.955 142.995 ;
        RECT 86.245 142.825 86.415 142.995 ;
        RECT 86.705 142.825 86.875 142.995 ;
        RECT 87.165 142.825 87.335 142.995 ;
        RECT 87.625 142.825 87.795 142.995 ;
        RECT 88.085 142.825 88.255 142.995 ;
        RECT 88.545 142.825 88.715 142.995 ;
        RECT 89.005 142.825 89.175 142.995 ;
        RECT 89.465 142.825 89.635 142.995 ;
        RECT 89.925 142.825 90.095 142.995 ;
        RECT 90.385 142.825 90.555 142.995 ;
        RECT 90.845 142.825 91.015 142.995 ;
        RECT 91.305 142.825 91.475 142.995 ;
        RECT 91.765 142.825 91.935 142.995 ;
        RECT 92.225 142.825 92.395 142.995 ;
        RECT 92.685 142.825 92.855 142.995 ;
        RECT 93.145 142.825 93.315 142.995 ;
        RECT 93.605 142.825 93.775 142.995 ;
        RECT 94.065 142.825 94.235 142.995 ;
        RECT 94.525 142.825 94.695 142.995 ;
        RECT 94.985 142.825 95.155 142.995 ;
        RECT 95.445 142.825 95.615 142.995 ;
        RECT 95.905 142.825 96.075 142.995 ;
        RECT 96.365 142.825 96.535 142.995 ;
        RECT 96.825 142.825 96.995 142.995 ;
        RECT 97.285 142.825 97.455 142.995 ;
        RECT 97.745 142.825 97.915 142.995 ;
        RECT 98.205 142.825 98.375 142.995 ;
        RECT 98.665 142.825 98.835 142.995 ;
        RECT 99.125 142.825 99.295 142.995 ;
        RECT 99.585 142.825 99.755 142.995 ;
        RECT 100.045 142.825 100.215 142.995 ;
        RECT 100.505 142.825 100.675 142.995 ;
        RECT 100.965 142.825 101.135 142.995 ;
        RECT 101.425 142.825 101.595 142.995 ;
        RECT 101.885 142.825 102.055 142.995 ;
        RECT 102.345 142.825 102.515 142.995 ;
        RECT 102.805 142.825 102.975 142.995 ;
        RECT 103.265 142.825 103.435 142.995 ;
        RECT 103.725 142.825 103.895 142.995 ;
        RECT 104.185 142.825 104.355 142.995 ;
        RECT 104.645 142.825 104.815 142.995 ;
        RECT 105.105 142.825 105.275 142.995 ;
        RECT 105.565 142.825 105.735 142.995 ;
        RECT 106.025 142.825 106.195 142.995 ;
        RECT 106.485 142.825 106.655 142.995 ;
        RECT 106.945 142.825 107.115 142.995 ;
        RECT 107.405 142.825 107.575 142.995 ;
        RECT 107.865 142.825 108.035 142.995 ;
        RECT 108.325 142.825 108.495 142.995 ;
        RECT 108.785 142.825 108.955 142.995 ;
        RECT 109.245 142.825 109.415 142.995 ;
        RECT 109.705 142.825 109.875 142.995 ;
        RECT 110.165 142.825 110.335 142.995 ;
        RECT 110.625 142.825 110.795 142.995 ;
        RECT 111.085 142.825 111.255 142.995 ;
        RECT 111.545 142.825 111.715 142.995 ;
        RECT 112.005 142.825 112.175 142.995 ;
        RECT 112.465 142.825 112.635 142.995 ;
        RECT 112.925 142.825 113.095 142.995 ;
        RECT 113.385 142.825 113.555 142.995 ;
        RECT 113.845 142.825 114.015 142.995 ;
        RECT 114.305 142.825 114.475 142.995 ;
        RECT 114.765 142.825 114.935 142.995 ;
        RECT 115.225 142.825 115.395 142.995 ;
        RECT 115.685 142.825 115.855 142.995 ;
        RECT 116.145 142.825 116.315 142.995 ;
        RECT 116.605 142.825 116.775 142.995 ;
        RECT 117.065 142.825 117.235 142.995 ;
        RECT 117.525 142.825 117.695 142.995 ;
        RECT 117.985 142.825 118.155 142.995 ;
        RECT 118.445 142.825 118.615 142.995 ;
        RECT 118.905 142.825 119.075 142.995 ;
        RECT 119.365 142.825 119.535 142.995 ;
        RECT 119.825 142.825 119.995 142.995 ;
        RECT 120.285 142.825 120.455 142.995 ;
        RECT 120.745 142.825 120.915 142.995 ;
        RECT 121.205 142.825 121.375 142.995 ;
        RECT 121.665 142.825 121.835 142.995 ;
        RECT 122.125 142.825 122.295 142.995 ;
        RECT 122.585 142.825 122.755 142.995 ;
        RECT 123.045 142.825 123.215 142.995 ;
        RECT 123.505 142.825 123.675 142.995 ;
        RECT 123.965 142.825 124.135 142.995 ;
        RECT 124.425 142.825 124.595 142.995 ;
        RECT 124.885 142.825 125.055 142.995 ;
        RECT 125.345 142.825 125.515 142.995 ;
        RECT 125.805 142.825 125.975 142.995 ;
        RECT 126.265 142.825 126.435 142.995 ;
        RECT 126.725 142.825 126.895 142.995 ;
        RECT 127.185 142.825 127.355 142.995 ;
        RECT 127.645 142.825 127.815 142.995 ;
        RECT 128.105 142.825 128.275 142.995 ;
        RECT 128.565 142.825 128.735 142.995 ;
        RECT 129.025 142.825 129.195 142.995 ;
        RECT 129.485 142.825 129.655 142.995 ;
        RECT 129.945 142.825 130.115 142.995 ;
        RECT 130.405 142.825 130.575 142.995 ;
        RECT 130.865 142.825 131.035 142.995 ;
        RECT 131.325 142.825 131.495 142.995 ;
        RECT 131.785 142.825 131.955 142.995 ;
        RECT 132.245 142.825 132.415 142.995 ;
        RECT 132.705 142.825 132.875 142.995 ;
        RECT 133.165 142.825 133.335 142.995 ;
        RECT 133.625 142.825 133.795 142.995 ;
        RECT 134.085 142.825 134.255 142.995 ;
        RECT 134.545 142.825 134.715 142.995 ;
        RECT 135.005 142.825 135.175 142.995 ;
        RECT 135.465 142.825 135.635 142.995 ;
        RECT 135.925 142.825 136.095 142.995 ;
        RECT 136.385 142.825 136.555 142.995 ;
        RECT 136.845 142.825 137.015 142.995 ;
        RECT 137.305 142.825 137.475 142.995 ;
        RECT 137.765 142.825 137.935 142.995 ;
        RECT 138.225 142.825 138.395 142.995 ;
        RECT 138.685 142.825 138.855 142.995 ;
        RECT 139.145 142.825 139.315 142.995 ;
        RECT 139.605 142.825 139.775 142.995 ;
        RECT 140.065 142.825 140.235 142.995 ;
        RECT 140.525 142.825 140.695 142.995 ;
        RECT 140.985 142.825 141.155 142.995 ;
        RECT 141.445 142.825 141.615 142.995 ;
        RECT 141.905 142.825 142.075 142.995 ;
        RECT 142.365 142.825 142.535 142.995 ;
        RECT 142.825 142.825 142.995 142.995 ;
        RECT 143.285 142.825 143.455 142.995 ;
        RECT 143.745 142.825 143.915 142.995 ;
        RECT 144.205 142.825 144.375 142.995 ;
        RECT 144.665 142.825 144.835 142.995 ;
        RECT 145.125 142.825 145.295 142.995 ;
        RECT 145.585 142.825 145.755 142.995 ;
        RECT 146.045 142.825 146.215 142.995 ;
        RECT 146.505 142.825 146.675 142.995 ;
        RECT 146.965 142.825 147.135 142.995 ;
        RECT 147.425 142.825 147.595 142.995 ;
        RECT 147.885 142.825 148.055 142.995 ;
        RECT 148.345 142.825 148.515 142.995 ;
        RECT 148.805 142.825 148.975 142.995 ;
        RECT 149.265 142.825 149.435 142.995 ;
        RECT 149.725 142.825 149.895 142.995 ;
        RECT 150.185 142.825 150.355 142.995 ;
        RECT 18.625 141.295 18.795 141.465 ;
        RECT 17.705 140.615 17.875 140.785 ;
        RECT 28.285 141.295 28.455 141.465 ;
        RECT 29.205 141.295 29.375 141.465 ;
        RECT 38.405 142.315 38.575 142.485 ;
        RECT 35.645 141.295 35.815 141.465 ;
        RECT 29.205 140.615 29.375 140.785 ;
        RECT 36.565 140.955 36.735 141.125 ;
        RECT 37.025 141.295 37.195 141.465 ;
        RECT 37.485 141.295 37.655 141.465 ;
        RECT 42.545 141.635 42.715 141.805 ;
        RECT 43.925 141.975 44.095 142.145 ;
        RECT 44.845 140.615 45.015 140.785 ;
        RECT 45.765 141.975 45.935 142.145 ;
        RECT 45.305 140.615 45.475 140.785 ;
        RECT 47.605 141.295 47.775 141.465 ;
        RECT 53.125 142.315 53.295 142.485 ;
        RECT 52.665 141.295 52.835 141.465 ;
        RECT 65.545 142.315 65.715 142.485 ;
        RECT 66.465 141.295 66.635 141.465 ;
        RECT 76.585 141.295 76.755 141.465 ;
        RECT 77.505 141.295 77.675 141.465 ;
        RECT 77.045 140.615 77.215 140.785 ;
        RECT 104.185 141.635 104.355 141.805 ;
        RECT 102.805 141.295 102.975 141.465 ;
        RECT 103.725 141.295 103.895 141.465 ;
        RECT 105.105 141.295 105.275 141.465 ;
        RECT 101.885 140.615 102.055 140.785 ;
        RECT 106.025 141.295 106.195 141.465 ;
        RECT 105.565 140.615 105.735 140.785 ;
        RECT 107.405 141.635 107.575 141.805 ;
        RECT 107.865 141.295 108.035 141.465 ;
        RECT 109.705 141.635 109.875 141.805 ;
        RECT 111.085 141.295 111.255 141.465 ;
        RECT 112.005 141.295 112.175 141.465 ;
        RECT 112.465 141.295 112.635 141.465 ;
        RECT 112.925 141.295 113.095 141.465 ;
        RECT 114.305 141.975 114.475 142.145 ;
        RECT 113.845 140.615 114.015 140.785 ;
        RECT 116.615 141.635 116.785 141.805 ;
        RECT 117.050 141.975 117.220 142.145 ;
        RECT 118.620 141.975 118.790 142.145 ;
        RECT 119.135 141.635 119.305 141.805 ;
        RECT 119.870 140.955 120.040 141.125 ;
        RECT 120.325 141.635 120.495 141.805 ;
        RECT 120.720 141.975 120.890 142.145 ;
        RECT 121.205 141.295 121.375 141.465 ;
        RECT 11.265 140.105 11.435 140.275 ;
        RECT 11.725 140.105 11.895 140.275 ;
        RECT 12.185 140.105 12.355 140.275 ;
        RECT 12.645 140.105 12.815 140.275 ;
        RECT 13.105 140.105 13.275 140.275 ;
        RECT 13.565 140.105 13.735 140.275 ;
        RECT 14.025 140.105 14.195 140.275 ;
        RECT 14.485 140.105 14.655 140.275 ;
        RECT 14.945 140.105 15.115 140.275 ;
        RECT 15.405 140.105 15.575 140.275 ;
        RECT 15.865 140.105 16.035 140.275 ;
        RECT 16.325 140.105 16.495 140.275 ;
        RECT 16.785 140.105 16.955 140.275 ;
        RECT 17.245 140.105 17.415 140.275 ;
        RECT 17.705 140.105 17.875 140.275 ;
        RECT 18.165 140.105 18.335 140.275 ;
        RECT 18.625 140.105 18.795 140.275 ;
        RECT 19.085 140.105 19.255 140.275 ;
        RECT 19.545 140.105 19.715 140.275 ;
        RECT 20.005 140.105 20.175 140.275 ;
        RECT 20.465 140.105 20.635 140.275 ;
        RECT 20.925 140.105 21.095 140.275 ;
        RECT 21.385 140.105 21.555 140.275 ;
        RECT 21.845 140.105 22.015 140.275 ;
        RECT 22.305 140.105 22.475 140.275 ;
        RECT 22.765 140.105 22.935 140.275 ;
        RECT 23.225 140.105 23.395 140.275 ;
        RECT 23.685 140.105 23.855 140.275 ;
        RECT 24.145 140.105 24.315 140.275 ;
        RECT 24.605 140.105 24.775 140.275 ;
        RECT 25.065 140.105 25.235 140.275 ;
        RECT 25.525 140.105 25.695 140.275 ;
        RECT 25.985 140.105 26.155 140.275 ;
        RECT 26.445 140.105 26.615 140.275 ;
        RECT 26.905 140.105 27.075 140.275 ;
        RECT 27.365 140.105 27.535 140.275 ;
        RECT 27.825 140.105 27.995 140.275 ;
        RECT 28.285 140.105 28.455 140.275 ;
        RECT 28.745 140.105 28.915 140.275 ;
        RECT 29.205 140.105 29.375 140.275 ;
        RECT 29.665 140.105 29.835 140.275 ;
        RECT 30.125 140.105 30.295 140.275 ;
        RECT 30.585 140.105 30.755 140.275 ;
        RECT 31.045 140.105 31.215 140.275 ;
        RECT 31.505 140.105 31.675 140.275 ;
        RECT 31.965 140.105 32.135 140.275 ;
        RECT 32.425 140.105 32.595 140.275 ;
        RECT 32.885 140.105 33.055 140.275 ;
        RECT 33.345 140.105 33.515 140.275 ;
        RECT 33.805 140.105 33.975 140.275 ;
        RECT 34.265 140.105 34.435 140.275 ;
        RECT 34.725 140.105 34.895 140.275 ;
        RECT 35.185 140.105 35.355 140.275 ;
        RECT 35.645 140.105 35.815 140.275 ;
        RECT 36.105 140.105 36.275 140.275 ;
        RECT 36.565 140.105 36.735 140.275 ;
        RECT 37.025 140.105 37.195 140.275 ;
        RECT 37.485 140.105 37.655 140.275 ;
        RECT 37.945 140.105 38.115 140.275 ;
        RECT 38.405 140.105 38.575 140.275 ;
        RECT 38.865 140.105 39.035 140.275 ;
        RECT 39.325 140.105 39.495 140.275 ;
        RECT 39.785 140.105 39.955 140.275 ;
        RECT 40.245 140.105 40.415 140.275 ;
        RECT 40.705 140.105 40.875 140.275 ;
        RECT 41.165 140.105 41.335 140.275 ;
        RECT 41.625 140.105 41.795 140.275 ;
        RECT 42.085 140.105 42.255 140.275 ;
        RECT 42.545 140.105 42.715 140.275 ;
        RECT 43.005 140.105 43.175 140.275 ;
        RECT 43.465 140.105 43.635 140.275 ;
        RECT 43.925 140.105 44.095 140.275 ;
        RECT 44.385 140.105 44.555 140.275 ;
        RECT 44.845 140.105 45.015 140.275 ;
        RECT 45.305 140.105 45.475 140.275 ;
        RECT 45.765 140.105 45.935 140.275 ;
        RECT 46.225 140.105 46.395 140.275 ;
        RECT 46.685 140.105 46.855 140.275 ;
        RECT 47.145 140.105 47.315 140.275 ;
        RECT 47.605 140.105 47.775 140.275 ;
        RECT 48.065 140.105 48.235 140.275 ;
        RECT 48.525 140.105 48.695 140.275 ;
        RECT 48.985 140.105 49.155 140.275 ;
        RECT 49.445 140.105 49.615 140.275 ;
        RECT 49.905 140.105 50.075 140.275 ;
        RECT 50.365 140.105 50.535 140.275 ;
        RECT 50.825 140.105 50.995 140.275 ;
        RECT 51.285 140.105 51.455 140.275 ;
        RECT 51.745 140.105 51.915 140.275 ;
        RECT 52.205 140.105 52.375 140.275 ;
        RECT 52.665 140.105 52.835 140.275 ;
        RECT 53.125 140.105 53.295 140.275 ;
        RECT 53.585 140.105 53.755 140.275 ;
        RECT 54.045 140.105 54.215 140.275 ;
        RECT 54.505 140.105 54.675 140.275 ;
        RECT 54.965 140.105 55.135 140.275 ;
        RECT 55.425 140.105 55.595 140.275 ;
        RECT 55.885 140.105 56.055 140.275 ;
        RECT 56.345 140.105 56.515 140.275 ;
        RECT 56.805 140.105 56.975 140.275 ;
        RECT 57.265 140.105 57.435 140.275 ;
        RECT 57.725 140.105 57.895 140.275 ;
        RECT 58.185 140.105 58.355 140.275 ;
        RECT 58.645 140.105 58.815 140.275 ;
        RECT 59.105 140.105 59.275 140.275 ;
        RECT 59.565 140.105 59.735 140.275 ;
        RECT 60.025 140.105 60.195 140.275 ;
        RECT 60.485 140.105 60.655 140.275 ;
        RECT 60.945 140.105 61.115 140.275 ;
        RECT 61.405 140.105 61.575 140.275 ;
        RECT 61.865 140.105 62.035 140.275 ;
        RECT 62.325 140.105 62.495 140.275 ;
        RECT 62.785 140.105 62.955 140.275 ;
        RECT 63.245 140.105 63.415 140.275 ;
        RECT 63.705 140.105 63.875 140.275 ;
        RECT 64.165 140.105 64.335 140.275 ;
        RECT 64.625 140.105 64.795 140.275 ;
        RECT 65.085 140.105 65.255 140.275 ;
        RECT 65.545 140.105 65.715 140.275 ;
        RECT 66.005 140.105 66.175 140.275 ;
        RECT 66.465 140.105 66.635 140.275 ;
        RECT 66.925 140.105 67.095 140.275 ;
        RECT 67.385 140.105 67.555 140.275 ;
        RECT 67.845 140.105 68.015 140.275 ;
        RECT 68.305 140.105 68.475 140.275 ;
        RECT 68.765 140.105 68.935 140.275 ;
        RECT 69.225 140.105 69.395 140.275 ;
        RECT 69.685 140.105 69.855 140.275 ;
        RECT 70.145 140.105 70.315 140.275 ;
        RECT 70.605 140.105 70.775 140.275 ;
        RECT 71.065 140.105 71.235 140.275 ;
        RECT 71.525 140.105 71.695 140.275 ;
        RECT 71.985 140.105 72.155 140.275 ;
        RECT 72.445 140.105 72.615 140.275 ;
        RECT 72.905 140.105 73.075 140.275 ;
        RECT 73.365 140.105 73.535 140.275 ;
        RECT 73.825 140.105 73.995 140.275 ;
        RECT 74.285 140.105 74.455 140.275 ;
        RECT 74.745 140.105 74.915 140.275 ;
        RECT 75.205 140.105 75.375 140.275 ;
        RECT 75.665 140.105 75.835 140.275 ;
        RECT 76.125 140.105 76.295 140.275 ;
        RECT 76.585 140.105 76.755 140.275 ;
        RECT 77.045 140.105 77.215 140.275 ;
        RECT 77.505 140.105 77.675 140.275 ;
        RECT 77.965 140.105 78.135 140.275 ;
        RECT 78.425 140.105 78.595 140.275 ;
        RECT 78.885 140.105 79.055 140.275 ;
        RECT 79.345 140.105 79.515 140.275 ;
        RECT 79.805 140.105 79.975 140.275 ;
        RECT 80.265 140.105 80.435 140.275 ;
        RECT 80.725 140.105 80.895 140.275 ;
        RECT 81.185 140.105 81.355 140.275 ;
        RECT 81.645 140.105 81.815 140.275 ;
        RECT 82.105 140.105 82.275 140.275 ;
        RECT 82.565 140.105 82.735 140.275 ;
        RECT 83.025 140.105 83.195 140.275 ;
        RECT 83.485 140.105 83.655 140.275 ;
        RECT 83.945 140.105 84.115 140.275 ;
        RECT 84.405 140.105 84.575 140.275 ;
        RECT 84.865 140.105 85.035 140.275 ;
        RECT 85.325 140.105 85.495 140.275 ;
        RECT 85.785 140.105 85.955 140.275 ;
        RECT 86.245 140.105 86.415 140.275 ;
        RECT 86.705 140.105 86.875 140.275 ;
        RECT 87.165 140.105 87.335 140.275 ;
        RECT 87.625 140.105 87.795 140.275 ;
        RECT 88.085 140.105 88.255 140.275 ;
        RECT 88.545 140.105 88.715 140.275 ;
        RECT 89.005 140.105 89.175 140.275 ;
        RECT 89.465 140.105 89.635 140.275 ;
        RECT 89.925 140.105 90.095 140.275 ;
        RECT 90.385 140.105 90.555 140.275 ;
        RECT 90.845 140.105 91.015 140.275 ;
        RECT 91.305 140.105 91.475 140.275 ;
        RECT 91.765 140.105 91.935 140.275 ;
        RECT 92.225 140.105 92.395 140.275 ;
        RECT 92.685 140.105 92.855 140.275 ;
        RECT 93.145 140.105 93.315 140.275 ;
        RECT 93.605 140.105 93.775 140.275 ;
        RECT 94.065 140.105 94.235 140.275 ;
        RECT 94.525 140.105 94.695 140.275 ;
        RECT 94.985 140.105 95.155 140.275 ;
        RECT 95.445 140.105 95.615 140.275 ;
        RECT 95.905 140.105 96.075 140.275 ;
        RECT 96.365 140.105 96.535 140.275 ;
        RECT 96.825 140.105 96.995 140.275 ;
        RECT 97.285 140.105 97.455 140.275 ;
        RECT 97.745 140.105 97.915 140.275 ;
        RECT 98.205 140.105 98.375 140.275 ;
        RECT 98.665 140.105 98.835 140.275 ;
        RECT 99.125 140.105 99.295 140.275 ;
        RECT 99.585 140.105 99.755 140.275 ;
        RECT 100.045 140.105 100.215 140.275 ;
        RECT 100.505 140.105 100.675 140.275 ;
        RECT 100.965 140.105 101.135 140.275 ;
        RECT 101.425 140.105 101.595 140.275 ;
        RECT 101.885 140.105 102.055 140.275 ;
        RECT 102.345 140.105 102.515 140.275 ;
        RECT 102.805 140.105 102.975 140.275 ;
        RECT 103.265 140.105 103.435 140.275 ;
        RECT 103.725 140.105 103.895 140.275 ;
        RECT 104.185 140.105 104.355 140.275 ;
        RECT 104.645 140.105 104.815 140.275 ;
        RECT 105.105 140.105 105.275 140.275 ;
        RECT 105.565 140.105 105.735 140.275 ;
        RECT 106.025 140.105 106.195 140.275 ;
        RECT 106.485 140.105 106.655 140.275 ;
        RECT 106.945 140.105 107.115 140.275 ;
        RECT 107.405 140.105 107.575 140.275 ;
        RECT 107.865 140.105 108.035 140.275 ;
        RECT 108.325 140.105 108.495 140.275 ;
        RECT 108.785 140.105 108.955 140.275 ;
        RECT 109.245 140.105 109.415 140.275 ;
        RECT 109.705 140.105 109.875 140.275 ;
        RECT 110.165 140.105 110.335 140.275 ;
        RECT 110.625 140.105 110.795 140.275 ;
        RECT 111.085 140.105 111.255 140.275 ;
        RECT 111.545 140.105 111.715 140.275 ;
        RECT 112.005 140.105 112.175 140.275 ;
        RECT 112.465 140.105 112.635 140.275 ;
        RECT 112.925 140.105 113.095 140.275 ;
        RECT 113.385 140.105 113.555 140.275 ;
        RECT 113.845 140.105 114.015 140.275 ;
        RECT 114.305 140.105 114.475 140.275 ;
        RECT 114.765 140.105 114.935 140.275 ;
        RECT 115.225 140.105 115.395 140.275 ;
        RECT 115.685 140.105 115.855 140.275 ;
        RECT 116.145 140.105 116.315 140.275 ;
        RECT 116.605 140.105 116.775 140.275 ;
        RECT 117.065 140.105 117.235 140.275 ;
        RECT 117.525 140.105 117.695 140.275 ;
        RECT 117.985 140.105 118.155 140.275 ;
        RECT 118.445 140.105 118.615 140.275 ;
        RECT 118.905 140.105 119.075 140.275 ;
        RECT 119.365 140.105 119.535 140.275 ;
        RECT 119.825 140.105 119.995 140.275 ;
        RECT 120.285 140.105 120.455 140.275 ;
        RECT 120.745 140.105 120.915 140.275 ;
        RECT 121.205 140.105 121.375 140.275 ;
        RECT 121.665 140.105 121.835 140.275 ;
        RECT 122.125 140.105 122.295 140.275 ;
        RECT 122.585 140.105 122.755 140.275 ;
        RECT 123.045 140.105 123.215 140.275 ;
        RECT 123.505 140.105 123.675 140.275 ;
        RECT 123.965 140.105 124.135 140.275 ;
        RECT 124.425 140.105 124.595 140.275 ;
        RECT 124.885 140.105 125.055 140.275 ;
        RECT 125.345 140.105 125.515 140.275 ;
        RECT 125.805 140.105 125.975 140.275 ;
        RECT 126.265 140.105 126.435 140.275 ;
        RECT 126.725 140.105 126.895 140.275 ;
        RECT 127.185 140.105 127.355 140.275 ;
        RECT 127.645 140.105 127.815 140.275 ;
        RECT 128.105 140.105 128.275 140.275 ;
        RECT 128.565 140.105 128.735 140.275 ;
        RECT 129.025 140.105 129.195 140.275 ;
        RECT 129.485 140.105 129.655 140.275 ;
        RECT 129.945 140.105 130.115 140.275 ;
        RECT 130.405 140.105 130.575 140.275 ;
        RECT 130.865 140.105 131.035 140.275 ;
        RECT 131.325 140.105 131.495 140.275 ;
        RECT 131.785 140.105 131.955 140.275 ;
        RECT 132.245 140.105 132.415 140.275 ;
        RECT 132.705 140.105 132.875 140.275 ;
        RECT 133.165 140.105 133.335 140.275 ;
        RECT 133.625 140.105 133.795 140.275 ;
        RECT 134.085 140.105 134.255 140.275 ;
        RECT 134.545 140.105 134.715 140.275 ;
        RECT 135.005 140.105 135.175 140.275 ;
        RECT 135.465 140.105 135.635 140.275 ;
        RECT 135.925 140.105 136.095 140.275 ;
        RECT 136.385 140.105 136.555 140.275 ;
        RECT 136.845 140.105 137.015 140.275 ;
        RECT 137.305 140.105 137.475 140.275 ;
        RECT 137.765 140.105 137.935 140.275 ;
        RECT 138.225 140.105 138.395 140.275 ;
        RECT 138.685 140.105 138.855 140.275 ;
        RECT 139.145 140.105 139.315 140.275 ;
        RECT 139.605 140.105 139.775 140.275 ;
        RECT 140.065 140.105 140.235 140.275 ;
        RECT 140.525 140.105 140.695 140.275 ;
        RECT 140.985 140.105 141.155 140.275 ;
        RECT 141.445 140.105 141.615 140.275 ;
        RECT 141.905 140.105 142.075 140.275 ;
        RECT 142.365 140.105 142.535 140.275 ;
        RECT 142.825 140.105 142.995 140.275 ;
        RECT 143.285 140.105 143.455 140.275 ;
        RECT 143.745 140.105 143.915 140.275 ;
        RECT 144.205 140.105 144.375 140.275 ;
        RECT 144.665 140.105 144.835 140.275 ;
        RECT 145.125 140.105 145.295 140.275 ;
        RECT 145.585 140.105 145.755 140.275 ;
        RECT 146.045 140.105 146.215 140.275 ;
        RECT 146.505 140.105 146.675 140.275 ;
        RECT 146.965 140.105 147.135 140.275 ;
        RECT 147.425 140.105 147.595 140.275 ;
        RECT 147.885 140.105 148.055 140.275 ;
        RECT 148.345 140.105 148.515 140.275 ;
        RECT 148.805 140.105 148.975 140.275 ;
        RECT 149.265 140.105 149.435 140.275 ;
        RECT 149.725 140.105 149.895 140.275 ;
        RECT 150.185 140.105 150.355 140.275 ;
        RECT 15.865 138.915 16.035 139.085 ;
        RECT 16.350 138.235 16.520 138.405 ;
        RECT 16.745 138.575 16.915 138.745 ;
        RECT 17.200 138.915 17.370 139.085 ;
        RECT 17.935 138.575 18.105 138.745 ;
        RECT 18.450 138.235 18.620 138.405 ;
        RECT 20.020 138.235 20.190 138.405 ;
        RECT 20.455 138.575 20.625 138.745 ;
        RECT 22.765 138.235 22.935 138.405 ;
        RECT 24.145 138.915 24.315 139.085 ;
        RECT 24.605 138.575 24.775 138.745 ;
        RECT 27.825 138.915 27.995 139.085 ;
        RECT 28.745 138.575 28.915 138.745 ;
        RECT 29.665 139.255 29.835 139.425 ;
        RECT 25.985 138.235 26.155 138.405 ;
        RECT 27.825 138.235 27.995 138.405 ;
        RECT 31.505 139.255 31.675 139.425 ;
        RECT 31.045 138.915 31.215 139.085 ;
        RECT 38.865 139.595 39.035 139.765 ;
        RECT 31.965 138.915 32.135 139.085 ;
        RECT 32.885 138.915 33.055 139.085 ;
        RECT 30.125 137.895 30.295 138.065 ;
        RECT 46.225 139.255 46.395 139.425 ;
        RECT 47.605 139.255 47.775 139.425 ;
        RECT 56.345 139.255 56.515 139.425 ;
        RECT 58.645 139.595 58.815 139.765 ;
        RECT 61.405 139.595 61.575 139.765 ;
        RECT 57.725 138.915 57.895 139.085 ;
        RECT 59.105 138.915 59.275 139.085 ;
        RECT 59.565 138.915 59.735 139.085 ;
        RECT 56.805 137.895 56.975 138.065 ;
        RECT 60.025 138.575 60.195 138.745 ;
        RECT 60.485 137.895 60.655 138.065 ;
        RECT 65.545 139.255 65.715 139.425 ;
        RECT 66.925 137.895 67.095 138.065 ;
        RECT 75.665 139.595 75.835 139.765 ;
        RECT 73.825 138.915 73.995 139.085 ;
        RECT 73.365 138.575 73.535 138.745 ;
        RECT 77.045 139.255 77.215 139.425 ;
        RECT 77.965 139.255 78.135 139.425 ;
        RECT 78.885 139.255 79.055 139.425 ;
        RECT 76.125 137.895 76.295 138.065 ;
        RECT 81.415 139.255 81.585 139.425 ;
        RECT 82.105 138.575 82.275 138.745 ;
        RECT 84.405 138.915 84.575 139.085 ;
        RECT 85.325 138.915 85.495 139.085 ;
        RECT 87.165 139.595 87.335 139.765 ;
        RECT 86.705 138.915 86.875 139.085 ;
        RECT 87.625 138.915 87.795 139.085 ;
        RECT 89.005 138.915 89.175 139.085 ;
        RECT 86.245 137.895 86.415 138.065 ;
        RECT 89.925 138.915 90.095 139.085 ;
        RECT 89.005 137.895 89.175 138.065 ;
        RECT 91.765 137.895 91.935 138.065 ;
        RECT 94.075 138.575 94.245 138.745 ;
        RECT 94.510 138.235 94.680 138.405 ;
        RECT 96.595 138.575 96.765 138.745 ;
        RECT 96.080 138.235 96.250 138.405 ;
        RECT 97.330 139.255 97.500 139.425 ;
        RECT 97.785 138.575 97.955 138.745 ;
        RECT 98.665 138.575 98.835 138.745 ;
        RECT 98.180 138.235 98.350 138.405 ;
        RECT 100.505 137.895 100.675 138.065 ;
        RECT 101.425 138.575 101.595 138.745 ;
        RECT 101.885 138.915 102.055 139.085 ;
        RECT 102.345 138.575 102.515 138.745 ;
        RECT 102.805 138.575 102.975 138.745 ;
        RECT 103.725 139.255 103.895 139.425 ;
        RECT 106.025 139.595 106.195 139.765 ;
        RECT 106.485 139.255 106.655 139.425 ;
        RECT 107.405 139.595 107.575 139.765 ;
        RECT 107.865 138.915 108.035 139.085 ;
        RECT 116.605 139.595 116.775 139.765 ;
        RECT 105.105 138.235 105.275 138.405 ;
        RECT 106.485 137.895 106.655 138.065 ;
        RECT 115.685 138.915 115.855 139.085 ;
        RECT 114.765 138.575 114.935 138.745 ;
        RECT 11.265 137.385 11.435 137.555 ;
        RECT 11.725 137.385 11.895 137.555 ;
        RECT 12.185 137.385 12.355 137.555 ;
        RECT 12.645 137.385 12.815 137.555 ;
        RECT 13.105 137.385 13.275 137.555 ;
        RECT 13.565 137.385 13.735 137.555 ;
        RECT 14.025 137.385 14.195 137.555 ;
        RECT 14.485 137.385 14.655 137.555 ;
        RECT 14.945 137.385 15.115 137.555 ;
        RECT 15.405 137.385 15.575 137.555 ;
        RECT 15.865 137.385 16.035 137.555 ;
        RECT 16.325 137.385 16.495 137.555 ;
        RECT 16.785 137.385 16.955 137.555 ;
        RECT 17.245 137.385 17.415 137.555 ;
        RECT 17.705 137.385 17.875 137.555 ;
        RECT 18.165 137.385 18.335 137.555 ;
        RECT 18.625 137.385 18.795 137.555 ;
        RECT 19.085 137.385 19.255 137.555 ;
        RECT 19.545 137.385 19.715 137.555 ;
        RECT 20.005 137.385 20.175 137.555 ;
        RECT 20.465 137.385 20.635 137.555 ;
        RECT 20.925 137.385 21.095 137.555 ;
        RECT 21.385 137.385 21.555 137.555 ;
        RECT 21.845 137.385 22.015 137.555 ;
        RECT 22.305 137.385 22.475 137.555 ;
        RECT 22.765 137.385 22.935 137.555 ;
        RECT 23.225 137.385 23.395 137.555 ;
        RECT 23.685 137.385 23.855 137.555 ;
        RECT 24.145 137.385 24.315 137.555 ;
        RECT 24.605 137.385 24.775 137.555 ;
        RECT 25.065 137.385 25.235 137.555 ;
        RECT 25.525 137.385 25.695 137.555 ;
        RECT 25.985 137.385 26.155 137.555 ;
        RECT 26.445 137.385 26.615 137.555 ;
        RECT 26.905 137.385 27.075 137.555 ;
        RECT 27.365 137.385 27.535 137.555 ;
        RECT 27.825 137.385 27.995 137.555 ;
        RECT 28.285 137.385 28.455 137.555 ;
        RECT 28.745 137.385 28.915 137.555 ;
        RECT 29.205 137.385 29.375 137.555 ;
        RECT 29.665 137.385 29.835 137.555 ;
        RECT 30.125 137.385 30.295 137.555 ;
        RECT 30.585 137.385 30.755 137.555 ;
        RECT 31.045 137.385 31.215 137.555 ;
        RECT 31.505 137.385 31.675 137.555 ;
        RECT 31.965 137.385 32.135 137.555 ;
        RECT 32.425 137.385 32.595 137.555 ;
        RECT 32.885 137.385 33.055 137.555 ;
        RECT 33.345 137.385 33.515 137.555 ;
        RECT 33.805 137.385 33.975 137.555 ;
        RECT 34.265 137.385 34.435 137.555 ;
        RECT 34.725 137.385 34.895 137.555 ;
        RECT 35.185 137.385 35.355 137.555 ;
        RECT 35.645 137.385 35.815 137.555 ;
        RECT 36.105 137.385 36.275 137.555 ;
        RECT 36.565 137.385 36.735 137.555 ;
        RECT 37.025 137.385 37.195 137.555 ;
        RECT 37.485 137.385 37.655 137.555 ;
        RECT 37.945 137.385 38.115 137.555 ;
        RECT 38.405 137.385 38.575 137.555 ;
        RECT 38.865 137.385 39.035 137.555 ;
        RECT 39.325 137.385 39.495 137.555 ;
        RECT 39.785 137.385 39.955 137.555 ;
        RECT 40.245 137.385 40.415 137.555 ;
        RECT 40.705 137.385 40.875 137.555 ;
        RECT 41.165 137.385 41.335 137.555 ;
        RECT 41.625 137.385 41.795 137.555 ;
        RECT 42.085 137.385 42.255 137.555 ;
        RECT 42.545 137.385 42.715 137.555 ;
        RECT 43.005 137.385 43.175 137.555 ;
        RECT 43.465 137.385 43.635 137.555 ;
        RECT 43.925 137.385 44.095 137.555 ;
        RECT 44.385 137.385 44.555 137.555 ;
        RECT 44.845 137.385 45.015 137.555 ;
        RECT 45.305 137.385 45.475 137.555 ;
        RECT 45.765 137.385 45.935 137.555 ;
        RECT 46.225 137.385 46.395 137.555 ;
        RECT 46.685 137.385 46.855 137.555 ;
        RECT 47.145 137.385 47.315 137.555 ;
        RECT 47.605 137.385 47.775 137.555 ;
        RECT 48.065 137.385 48.235 137.555 ;
        RECT 48.525 137.385 48.695 137.555 ;
        RECT 48.985 137.385 49.155 137.555 ;
        RECT 49.445 137.385 49.615 137.555 ;
        RECT 49.905 137.385 50.075 137.555 ;
        RECT 50.365 137.385 50.535 137.555 ;
        RECT 50.825 137.385 50.995 137.555 ;
        RECT 51.285 137.385 51.455 137.555 ;
        RECT 51.745 137.385 51.915 137.555 ;
        RECT 52.205 137.385 52.375 137.555 ;
        RECT 52.665 137.385 52.835 137.555 ;
        RECT 53.125 137.385 53.295 137.555 ;
        RECT 53.585 137.385 53.755 137.555 ;
        RECT 54.045 137.385 54.215 137.555 ;
        RECT 54.505 137.385 54.675 137.555 ;
        RECT 54.965 137.385 55.135 137.555 ;
        RECT 55.425 137.385 55.595 137.555 ;
        RECT 55.885 137.385 56.055 137.555 ;
        RECT 56.345 137.385 56.515 137.555 ;
        RECT 56.805 137.385 56.975 137.555 ;
        RECT 57.265 137.385 57.435 137.555 ;
        RECT 57.725 137.385 57.895 137.555 ;
        RECT 58.185 137.385 58.355 137.555 ;
        RECT 58.645 137.385 58.815 137.555 ;
        RECT 59.105 137.385 59.275 137.555 ;
        RECT 59.565 137.385 59.735 137.555 ;
        RECT 60.025 137.385 60.195 137.555 ;
        RECT 60.485 137.385 60.655 137.555 ;
        RECT 60.945 137.385 61.115 137.555 ;
        RECT 61.405 137.385 61.575 137.555 ;
        RECT 61.865 137.385 62.035 137.555 ;
        RECT 62.325 137.385 62.495 137.555 ;
        RECT 62.785 137.385 62.955 137.555 ;
        RECT 63.245 137.385 63.415 137.555 ;
        RECT 63.705 137.385 63.875 137.555 ;
        RECT 64.165 137.385 64.335 137.555 ;
        RECT 64.625 137.385 64.795 137.555 ;
        RECT 65.085 137.385 65.255 137.555 ;
        RECT 65.545 137.385 65.715 137.555 ;
        RECT 66.005 137.385 66.175 137.555 ;
        RECT 66.465 137.385 66.635 137.555 ;
        RECT 66.925 137.385 67.095 137.555 ;
        RECT 67.385 137.385 67.555 137.555 ;
        RECT 67.845 137.385 68.015 137.555 ;
        RECT 68.305 137.385 68.475 137.555 ;
        RECT 68.765 137.385 68.935 137.555 ;
        RECT 69.225 137.385 69.395 137.555 ;
        RECT 69.685 137.385 69.855 137.555 ;
        RECT 70.145 137.385 70.315 137.555 ;
        RECT 70.605 137.385 70.775 137.555 ;
        RECT 71.065 137.385 71.235 137.555 ;
        RECT 71.525 137.385 71.695 137.555 ;
        RECT 71.985 137.385 72.155 137.555 ;
        RECT 72.445 137.385 72.615 137.555 ;
        RECT 72.905 137.385 73.075 137.555 ;
        RECT 73.365 137.385 73.535 137.555 ;
        RECT 73.825 137.385 73.995 137.555 ;
        RECT 74.285 137.385 74.455 137.555 ;
        RECT 74.745 137.385 74.915 137.555 ;
        RECT 75.205 137.385 75.375 137.555 ;
        RECT 75.665 137.385 75.835 137.555 ;
        RECT 76.125 137.385 76.295 137.555 ;
        RECT 76.585 137.385 76.755 137.555 ;
        RECT 77.045 137.385 77.215 137.555 ;
        RECT 77.505 137.385 77.675 137.555 ;
        RECT 77.965 137.385 78.135 137.555 ;
        RECT 78.425 137.385 78.595 137.555 ;
        RECT 78.885 137.385 79.055 137.555 ;
        RECT 79.345 137.385 79.515 137.555 ;
        RECT 79.805 137.385 79.975 137.555 ;
        RECT 80.265 137.385 80.435 137.555 ;
        RECT 80.725 137.385 80.895 137.555 ;
        RECT 81.185 137.385 81.355 137.555 ;
        RECT 81.645 137.385 81.815 137.555 ;
        RECT 82.105 137.385 82.275 137.555 ;
        RECT 82.565 137.385 82.735 137.555 ;
        RECT 83.025 137.385 83.195 137.555 ;
        RECT 83.485 137.385 83.655 137.555 ;
        RECT 83.945 137.385 84.115 137.555 ;
        RECT 84.405 137.385 84.575 137.555 ;
        RECT 84.865 137.385 85.035 137.555 ;
        RECT 85.325 137.385 85.495 137.555 ;
        RECT 85.785 137.385 85.955 137.555 ;
        RECT 86.245 137.385 86.415 137.555 ;
        RECT 86.705 137.385 86.875 137.555 ;
        RECT 87.165 137.385 87.335 137.555 ;
        RECT 87.625 137.385 87.795 137.555 ;
        RECT 88.085 137.385 88.255 137.555 ;
        RECT 88.545 137.385 88.715 137.555 ;
        RECT 89.005 137.385 89.175 137.555 ;
        RECT 89.465 137.385 89.635 137.555 ;
        RECT 89.925 137.385 90.095 137.555 ;
        RECT 90.385 137.385 90.555 137.555 ;
        RECT 90.845 137.385 91.015 137.555 ;
        RECT 91.305 137.385 91.475 137.555 ;
        RECT 91.765 137.385 91.935 137.555 ;
        RECT 92.225 137.385 92.395 137.555 ;
        RECT 92.685 137.385 92.855 137.555 ;
        RECT 93.145 137.385 93.315 137.555 ;
        RECT 93.605 137.385 93.775 137.555 ;
        RECT 94.065 137.385 94.235 137.555 ;
        RECT 94.525 137.385 94.695 137.555 ;
        RECT 94.985 137.385 95.155 137.555 ;
        RECT 95.445 137.385 95.615 137.555 ;
        RECT 95.905 137.385 96.075 137.555 ;
        RECT 96.365 137.385 96.535 137.555 ;
        RECT 96.825 137.385 96.995 137.555 ;
        RECT 97.285 137.385 97.455 137.555 ;
        RECT 97.745 137.385 97.915 137.555 ;
        RECT 98.205 137.385 98.375 137.555 ;
        RECT 98.665 137.385 98.835 137.555 ;
        RECT 99.125 137.385 99.295 137.555 ;
        RECT 99.585 137.385 99.755 137.555 ;
        RECT 100.045 137.385 100.215 137.555 ;
        RECT 100.505 137.385 100.675 137.555 ;
        RECT 100.965 137.385 101.135 137.555 ;
        RECT 101.425 137.385 101.595 137.555 ;
        RECT 101.885 137.385 102.055 137.555 ;
        RECT 102.345 137.385 102.515 137.555 ;
        RECT 102.805 137.385 102.975 137.555 ;
        RECT 103.265 137.385 103.435 137.555 ;
        RECT 103.725 137.385 103.895 137.555 ;
        RECT 104.185 137.385 104.355 137.555 ;
        RECT 104.645 137.385 104.815 137.555 ;
        RECT 105.105 137.385 105.275 137.555 ;
        RECT 105.565 137.385 105.735 137.555 ;
        RECT 106.025 137.385 106.195 137.555 ;
        RECT 106.485 137.385 106.655 137.555 ;
        RECT 106.945 137.385 107.115 137.555 ;
        RECT 107.405 137.385 107.575 137.555 ;
        RECT 107.865 137.385 108.035 137.555 ;
        RECT 108.325 137.385 108.495 137.555 ;
        RECT 108.785 137.385 108.955 137.555 ;
        RECT 109.245 137.385 109.415 137.555 ;
        RECT 109.705 137.385 109.875 137.555 ;
        RECT 110.165 137.385 110.335 137.555 ;
        RECT 110.625 137.385 110.795 137.555 ;
        RECT 111.085 137.385 111.255 137.555 ;
        RECT 111.545 137.385 111.715 137.555 ;
        RECT 112.005 137.385 112.175 137.555 ;
        RECT 112.465 137.385 112.635 137.555 ;
        RECT 112.925 137.385 113.095 137.555 ;
        RECT 113.385 137.385 113.555 137.555 ;
        RECT 113.845 137.385 114.015 137.555 ;
        RECT 114.305 137.385 114.475 137.555 ;
        RECT 114.765 137.385 114.935 137.555 ;
        RECT 115.225 137.385 115.395 137.555 ;
        RECT 115.685 137.385 115.855 137.555 ;
        RECT 116.145 137.385 116.315 137.555 ;
        RECT 116.605 137.385 116.775 137.555 ;
        RECT 117.065 137.385 117.235 137.555 ;
        RECT 117.525 137.385 117.695 137.555 ;
        RECT 117.985 137.385 118.155 137.555 ;
        RECT 118.445 137.385 118.615 137.555 ;
        RECT 118.905 137.385 119.075 137.555 ;
        RECT 119.365 137.385 119.535 137.555 ;
        RECT 119.825 137.385 119.995 137.555 ;
        RECT 120.285 137.385 120.455 137.555 ;
        RECT 120.745 137.385 120.915 137.555 ;
        RECT 121.205 137.385 121.375 137.555 ;
        RECT 121.665 137.385 121.835 137.555 ;
        RECT 122.125 137.385 122.295 137.555 ;
        RECT 122.585 137.385 122.755 137.555 ;
        RECT 123.045 137.385 123.215 137.555 ;
        RECT 123.505 137.385 123.675 137.555 ;
        RECT 123.965 137.385 124.135 137.555 ;
        RECT 124.425 137.385 124.595 137.555 ;
        RECT 124.885 137.385 125.055 137.555 ;
        RECT 125.345 137.385 125.515 137.555 ;
        RECT 125.805 137.385 125.975 137.555 ;
        RECT 126.265 137.385 126.435 137.555 ;
        RECT 126.725 137.385 126.895 137.555 ;
        RECT 127.185 137.385 127.355 137.555 ;
        RECT 127.645 137.385 127.815 137.555 ;
        RECT 128.105 137.385 128.275 137.555 ;
        RECT 128.565 137.385 128.735 137.555 ;
        RECT 129.025 137.385 129.195 137.555 ;
        RECT 129.485 137.385 129.655 137.555 ;
        RECT 129.945 137.385 130.115 137.555 ;
        RECT 130.405 137.385 130.575 137.555 ;
        RECT 130.865 137.385 131.035 137.555 ;
        RECT 131.325 137.385 131.495 137.555 ;
        RECT 131.785 137.385 131.955 137.555 ;
        RECT 132.245 137.385 132.415 137.555 ;
        RECT 132.705 137.385 132.875 137.555 ;
        RECT 133.165 137.385 133.335 137.555 ;
        RECT 133.625 137.385 133.795 137.555 ;
        RECT 134.085 137.385 134.255 137.555 ;
        RECT 134.545 137.385 134.715 137.555 ;
        RECT 135.005 137.385 135.175 137.555 ;
        RECT 135.465 137.385 135.635 137.555 ;
        RECT 135.925 137.385 136.095 137.555 ;
        RECT 136.385 137.385 136.555 137.555 ;
        RECT 136.845 137.385 137.015 137.555 ;
        RECT 137.305 137.385 137.475 137.555 ;
        RECT 137.765 137.385 137.935 137.555 ;
        RECT 138.225 137.385 138.395 137.555 ;
        RECT 138.685 137.385 138.855 137.555 ;
        RECT 139.145 137.385 139.315 137.555 ;
        RECT 139.605 137.385 139.775 137.555 ;
        RECT 140.065 137.385 140.235 137.555 ;
        RECT 140.525 137.385 140.695 137.555 ;
        RECT 140.985 137.385 141.155 137.555 ;
        RECT 141.445 137.385 141.615 137.555 ;
        RECT 141.905 137.385 142.075 137.555 ;
        RECT 142.365 137.385 142.535 137.555 ;
        RECT 142.825 137.385 142.995 137.555 ;
        RECT 143.285 137.385 143.455 137.555 ;
        RECT 143.745 137.385 143.915 137.555 ;
        RECT 144.205 137.385 144.375 137.555 ;
        RECT 144.665 137.385 144.835 137.555 ;
        RECT 145.125 137.385 145.295 137.555 ;
        RECT 145.585 137.385 145.755 137.555 ;
        RECT 146.045 137.385 146.215 137.555 ;
        RECT 146.505 137.385 146.675 137.555 ;
        RECT 146.965 137.385 147.135 137.555 ;
        RECT 147.425 137.385 147.595 137.555 ;
        RECT 147.885 137.385 148.055 137.555 ;
        RECT 148.345 137.385 148.515 137.555 ;
        RECT 148.805 137.385 148.975 137.555 ;
        RECT 149.265 137.385 149.435 137.555 ;
        RECT 149.725 137.385 149.895 137.555 ;
        RECT 150.185 137.385 150.355 137.555 ;
        RECT 18.625 136.875 18.795 137.045 ;
        RECT 19.545 135.855 19.715 136.025 ;
        RECT 20.465 135.855 20.635 136.025 ;
        RECT 26.905 136.195 27.075 136.365 ;
        RECT 27.365 135.855 27.535 136.025 ;
        RECT 29.205 136.535 29.375 136.705 ;
        RECT 37.485 136.875 37.655 137.045 ;
        RECT 39.785 136.195 39.955 136.365 ;
        RECT 39.325 135.855 39.495 136.025 ;
        RECT 41.625 135.855 41.795 136.025 ;
        RECT 43.005 135.855 43.175 136.025 ;
        RECT 42.085 135.515 42.255 135.685 ;
        RECT 46.685 136.875 46.855 137.045 ;
        RECT 47.605 136.875 47.775 137.045 ;
        RECT 45.765 136.195 45.935 136.365 ;
        RECT 48.065 136.535 48.235 136.705 ;
        RECT 44.385 135.515 44.555 135.685 ;
        RECT 46.685 135.855 46.855 136.025 ;
        RECT 43.925 135.175 44.095 135.345 ;
        RECT 48.065 135.855 48.235 136.025 ;
        RECT 53.585 136.875 53.755 137.045 ;
        RECT 48.985 135.855 49.155 136.025 ;
        RECT 52.205 136.195 52.375 136.365 ;
        RECT 51.745 135.855 51.915 136.025 ;
        RECT 60.025 136.875 60.195 137.045 ;
        RECT 57.265 135.855 57.435 136.025 ;
        RECT 58.645 136.195 58.815 136.365 ;
        RECT 58.185 135.855 58.355 136.025 ;
        RECT 57.725 135.515 57.895 135.685 ;
        RECT 62.325 136.875 62.495 137.045 ;
        RECT 60.945 135.855 61.115 136.025 ;
        RECT 65.110 136.535 65.280 136.705 ;
        RECT 61.405 135.175 61.575 135.345 ;
        RECT 62.245 135.175 62.415 135.345 ;
        RECT 64.625 136.195 64.795 136.365 ;
        RECT 63.245 135.515 63.415 135.685 ;
        RECT 65.505 136.195 65.675 136.365 ;
        RECT 65.960 135.515 66.130 135.685 ;
        RECT 67.210 136.535 67.380 136.705 ;
        RECT 66.695 136.195 66.865 136.365 ;
        RECT 68.780 136.535 68.950 136.705 ;
        RECT 69.215 136.195 69.385 136.365 ;
        RECT 71.525 136.875 71.695 137.045 ;
        RECT 73.365 136.875 73.535 137.045 ;
        RECT 77.045 136.875 77.215 137.045 ;
        RECT 72.445 135.175 72.615 135.345 ;
        RECT 73.285 135.175 73.455 135.345 ;
        RECT 74.285 135.515 74.455 135.685 ;
        RECT 76.965 135.515 77.135 135.685 ;
        RECT 76.125 135.175 76.295 135.345 ;
        RECT 77.965 135.515 78.135 135.685 ;
        RECT 83.485 136.875 83.655 137.045 ;
        RECT 82.105 135.855 82.275 136.025 ;
        RECT 82.565 135.515 82.735 135.685 ;
        RECT 83.485 135.855 83.655 136.025 ;
        RECT 83.945 135.855 84.115 136.025 ;
        RECT 84.865 135.855 85.035 136.025 ;
        RECT 84.405 135.175 84.575 135.345 ;
        RECT 89.005 136.195 89.175 136.365 ;
        RECT 88.545 135.855 88.715 136.025 ;
        RECT 90.385 136.195 90.555 136.365 ;
        RECT 94.985 136.535 95.155 136.705 ;
        RECT 92.225 135.855 92.395 136.025 ;
        RECT 93.145 135.855 93.315 136.025 ;
        RECT 93.605 135.855 93.775 136.025 ;
        RECT 94.065 135.855 94.235 136.025 ;
        RECT 95.445 135.855 95.615 136.025 ;
        RECT 96.365 135.855 96.535 136.025 ;
        RECT 97.285 135.855 97.455 136.025 ;
        RECT 97.745 136.875 97.915 137.045 ;
        RECT 98.665 135.855 98.835 136.025 ;
        RECT 11.265 134.665 11.435 134.835 ;
        RECT 11.725 134.665 11.895 134.835 ;
        RECT 12.185 134.665 12.355 134.835 ;
        RECT 12.645 134.665 12.815 134.835 ;
        RECT 13.105 134.665 13.275 134.835 ;
        RECT 13.565 134.665 13.735 134.835 ;
        RECT 14.025 134.665 14.195 134.835 ;
        RECT 14.485 134.665 14.655 134.835 ;
        RECT 14.945 134.665 15.115 134.835 ;
        RECT 15.405 134.665 15.575 134.835 ;
        RECT 15.865 134.665 16.035 134.835 ;
        RECT 16.325 134.665 16.495 134.835 ;
        RECT 16.785 134.665 16.955 134.835 ;
        RECT 17.245 134.665 17.415 134.835 ;
        RECT 17.705 134.665 17.875 134.835 ;
        RECT 18.165 134.665 18.335 134.835 ;
        RECT 18.625 134.665 18.795 134.835 ;
        RECT 19.085 134.665 19.255 134.835 ;
        RECT 19.545 134.665 19.715 134.835 ;
        RECT 20.005 134.665 20.175 134.835 ;
        RECT 20.465 134.665 20.635 134.835 ;
        RECT 20.925 134.665 21.095 134.835 ;
        RECT 21.385 134.665 21.555 134.835 ;
        RECT 21.845 134.665 22.015 134.835 ;
        RECT 22.305 134.665 22.475 134.835 ;
        RECT 22.765 134.665 22.935 134.835 ;
        RECT 23.225 134.665 23.395 134.835 ;
        RECT 23.685 134.665 23.855 134.835 ;
        RECT 24.145 134.665 24.315 134.835 ;
        RECT 24.605 134.665 24.775 134.835 ;
        RECT 25.065 134.665 25.235 134.835 ;
        RECT 25.525 134.665 25.695 134.835 ;
        RECT 25.985 134.665 26.155 134.835 ;
        RECT 26.445 134.665 26.615 134.835 ;
        RECT 26.905 134.665 27.075 134.835 ;
        RECT 27.365 134.665 27.535 134.835 ;
        RECT 27.825 134.665 27.995 134.835 ;
        RECT 28.285 134.665 28.455 134.835 ;
        RECT 28.745 134.665 28.915 134.835 ;
        RECT 29.205 134.665 29.375 134.835 ;
        RECT 29.665 134.665 29.835 134.835 ;
        RECT 30.125 134.665 30.295 134.835 ;
        RECT 30.585 134.665 30.755 134.835 ;
        RECT 31.045 134.665 31.215 134.835 ;
        RECT 31.505 134.665 31.675 134.835 ;
        RECT 31.965 134.665 32.135 134.835 ;
        RECT 32.425 134.665 32.595 134.835 ;
        RECT 32.885 134.665 33.055 134.835 ;
        RECT 33.345 134.665 33.515 134.835 ;
        RECT 33.805 134.665 33.975 134.835 ;
        RECT 34.265 134.665 34.435 134.835 ;
        RECT 34.725 134.665 34.895 134.835 ;
        RECT 35.185 134.665 35.355 134.835 ;
        RECT 35.645 134.665 35.815 134.835 ;
        RECT 36.105 134.665 36.275 134.835 ;
        RECT 36.565 134.665 36.735 134.835 ;
        RECT 37.025 134.665 37.195 134.835 ;
        RECT 37.485 134.665 37.655 134.835 ;
        RECT 37.945 134.665 38.115 134.835 ;
        RECT 38.405 134.665 38.575 134.835 ;
        RECT 38.865 134.665 39.035 134.835 ;
        RECT 39.325 134.665 39.495 134.835 ;
        RECT 39.785 134.665 39.955 134.835 ;
        RECT 40.245 134.665 40.415 134.835 ;
        RECT 40.705 134.665 40.875 134.835 ;
        RECT 41.165 134.665 41.335 134.835 ;
        RECT 41.625 134.665 41.795 134.835 ;
        RECT 42.085 134.665 42.255 134.835 ;
        RECT 42.545 134.665 42.715 134.835 ;
        RECT 43.005 134.665 43.175 134.835 ;
        RECT 43.465 134.665 43.635 134.835 ;
        RECT 43.925 134.665 44.095 134.835 ;
        RECT 44.385 134.665 44.555 134.835 ;
        RECT 44.845 134.665 45.015 134.835 ;
        RECT 45.305 134.665 45.475 134.835 ;
        RECT 45.765 134.665 45.935 134.835 ;
        RECT 46.225 134.665 46.395 134.835 ;
        RECT 46.685 134.665 46.855 134.835 ;
        RECT 47.145 134.665 47.315 134.835 ;
        RECT 47.605 134.665 47.775 134.835 ;
        RECT 48.065 134.665 48.235 134.835 ;
        RECT 48.525 134.665 48.695 134.835 ;
        RECT 48.985 134.665 49.155 134.835 ;
        RECT 49.445 134.665 49.615 134.835 ;
        RECT 49.905 134.665 50.075 134.835 ;
        RECT 50.365 134.665 50.535 134.835 ;
        RECT 50.825 134.665 50.995 134.835 ;
        RECT 51.285 134.665 51.455 134.835 ;
        RECT 51.745 134.665 51.915 134.835 ;
        RECT 52.205 134.665 52.375 134.835 ;
        RECT 52.665 134.665 52.835 134.835 ;
        RECT 53.125 134.665 53.295 134.835 ;
        RECT 53.585 134.665 53.755 134.835 ;
        RECT 54.045 134.665 54.215 134.835 ;
        RECT 54.505 134.665 54.675 134.835 ;
        RECT 54.965 134.665 55.135 134.835 ;
        RECT 55.425 134.665 55.595 134.835 ;
        RECT 55.885 134.665 56.055 134.835 ;
        RECT 56.345 134.665 56.515 134.835 ;
        RECT 56.805 134.665 56.975 134.835 ;
        RECT 57.265 134.665 57.435 134.835 ;
        RECT 57.725 134.665 57.895 134.835 ;
        RECT 58.185 134.665 58.355 134.835 ;
        RECT 58.645 134.665 58.815 134.835 ;
        RECT 59.105 134.665 59.275 134.835 ;
        RECT 59.565 134.665 59.735 134.835 ;
        RECT 60.025 134.665 60.195 134.835 ;
        RECT 60.485 134.665 60.655 134.835 ;
        RECT 60.945 134.665 61.115 134.835 ;
        RECT 61.405 134.665 61.575 134.835 ;
        RECT 61.865 134.665 62.035 134.835 ;
        RECT 62.325 134.665 62.495 134.835 ;
        RECT 62.785 134.665 62.955 134.835 ;
        RECT 63.245 134.665 63.415 134.835 ;
        RECT 63.705 134.665 63.875 134.835 ;
        RECT 64.165 134.665 64.335 134.835 ;
        RECT 64.625 134.665 64.795 134.835 ;
        RECT 65.085 134.665 65.255 134.835 ;
        RECT 65.545 134.665 65.715 134.835 ;
        RECT 66.005 134.665 66.175 134.835 ;
        RECT 66.465 134.665 66.635 134.835 ;
        RECT 66.925 134.665 67.095 134.835 ;
        RECT 67.385 134.665 67.555 134.835 ;
        RECT 67.845 134.665 68.015 134.835 ;
        RECT 68.305 134.665 68.475 134.835 ;
        RECT 68.765 134.665 68.935 134.835 ;
        RECT 69.225 134.665 69.395 134.835 ;
        RECT 69.685 134.665 69.855 134.835 ;
        RECT 70.145 134.665 70.315 134.835 ;
        RECT 70.605 134.665 70.775 134.835 ;
        RECT 71.065 134.665 71.235 134.835 ;
        RECT 71.525 134.665 71.695 134.835 ;
        RECT 71.985 134.665 72.155 134.835 ;
        RECT 72.445 134.665 72.615 134.835 ;
        RECT 72.905 134.665 73.075 134.835 ;
        RECT 73.365 134.665 73.535 134.835 ;
        RECT 73.825 134.665 73.995 134.835 ;
        RECT 74.285 134.665 74.455 134.835 ;
        RECT 74.745 134.665 74.915 134.835 ;
        RECT 75.205 134.665 75.375 134.835 ;
        RECT 75.665 134.665 75.835 134.835 ;
        RECT 76.125 134.665 76.295 134.835 ;
        RECT 76.585 134.665 76.755 134.835 ;
        RECT 77.045 134.665 77.215 134.835 ;
        RECT 77.505 134.665 77.675 134.835 ;
        RECT 77.965 134.665 78.135 134.835 ;
        RECT 78.425 134.665 78.595 134.835 ;
        RECT 78.885 134.665 79.055 134.835 ;
        RECT 79.345 134.665 79.515 134.835 ;
        RECT 79.805 134.665 79.975 134.835 ;
        RECT 80.265 134.665 80.435 134.835 ;
        RECT 80.725 134.665 80.895 134.835 ;
        RECT 81.185 134.665 81.355 134.835 ;
        RECT 81.645 134.665 81.815 134.835 ;
        RECT 82.105 134.665 82.275 134.835 ;
        RECT 82.565 134.665 82.735 134.835 ;
        RECT 83.025 134.665 83.195 134.835 ;
        RECT 83.485 134.665 83.655 134.835 ;
        RECT 83.945 134.665 84.115 134.835 ;
        RECT 84.405 134.665 84.575 134.835 ;
        RECT 84.865 134.665 85.035 134.835 ;
        RECT 85.325 134.665 85.495 134.835 ;
        RECT 85.785 134.665 85.955 134.835 ;
        RECT 86.245 134.665 86.415 134.835 ;
        RECT 86.705 134.665 86.875 134.835 ;
        RECT 87.165 134.665 87.335 134.835 ;
        RECT 87.625 134.665 87.795 134.835 ;
        RECT 88.085 134.665 88.255 134.835 ;
        RECT 88.545 134.665 88.715 134.835 ;
        RECT 89.005 134.665 89.175 134.835 ;
        RECT 89.465 134.665 89.635 134.835 ;
        RECT 89.925 134.665 90.095 134.835 ;
        RECT 90.385 134.665 90.555 134.835 ;
        RECT 90.845 134.665 91.015 134.835 ;
        RECT 91.305 134.665 91.475 134.835 ;
        RECT 91.765 134.665 91.935 134.835 ;
        RECT 92.225 134.665 92.395 134.835 ;
        RECT 92.685 134.665 92.855 134.835 ;
        RECT 93.145 134.665 93.315 134.835 ;
        RECT 93.605 134.665 93.775 134.835 ;
        RECT 94.065 134.665 94.235 134.835 ;
        RECT 94.525 134.665 94.695 134.835 ;
        RECT 94.985 134.665 95.155 134.835 ;
        RECT 95.445 134.665 95.615 134.835 ;
        RECT 95.905 134.665 96.075 134.835 ;
        RECT 96.365 134.665 96.535 134.835 ;
        RECT 96.825 134.665 96.995 134.835 ;
        RECT 97.285 134.665 97.455 134.835 ;
        RECT 97.745 134.665 97.915 134.835 ;
        RECT 98.205 134.665 98.375 134.835 ;
        RECT 98.665 134.665 98.835 134.835 ;
        RECT 99.125 134.665 99.295 134.835 ;
        RECT 99.585 134.665 99.755 134.835 ;
        RECT 100.045 134.665 100.215 134.835 ;
        RECT 100.505 134.665 100.675 134.835 ;
        RECT 100.965 134.665 101.135 134.835 ;
        RECT 101.425 134.665 101.595 134.835 ;
        RECT 101.885 134.665 102.055 134.835 ;
        RECT 102.345 134.665 102.515 134.835 ;
        RECT 102.805 134.665 102.975 134.835 ;
        RECT 103.265 134.665 103.435 134.835 ;
        RECT 103.725 134.665 103.895 134.835 ;
        RECT 104.185 134.665 104.355 134.835 ;
        RECT 104.645 134.665 104.815 134.835 ;
        RECT 105.105 134.665 105.275 134.835 ;
        RECT 105.565 134.665 105.735 134.835 ;
        RECT 106.025 134.665 106.195 134.835 ;
        RECT 106.485 134.665 106.655 134.835 ;
        RECT 106.945 134.665 107.115 134.835 ;
        RECT 107.405 134.665 107.575 134.835 ;
        RECT 107.865 134.665 108.035 134.835 ;
        RECT 108.325 134.665 108.495 134.835 ;
        RECT 108.785 134.665 108.955 134.835 ;
        RECT 109.245 134.665 109.415 134.835 ;
        RECT 109.705 134.665 109.875 134.835 ;
        RECT 110.165 134.665 110.335 134.835 ;
        RECT 110.625 134.665 110.795 134.835 ;
        RECT 111.085 134.665 111.255 134.835 ;
        RECT 111.545 134.665 111.715 134.835 ;
        RECT 112.005 134.665 112.175 134.835 ;
        RECT 112.465 134.665 112.635 134.835 ;
        RECT 112.925 134.665 113.095 134.835 ;
        RECT 113.385 134.665 113.555 134.835 ;
        RECT 113.845 134.665 114.015 134.835 ;
        RECT 114.305 134.665 114.475 134.835 ;
        RECT 114.765 134.665 114.935 134.835 ;
        RECT 115.225 134.665 115.395 134.835 ;
        RECT 115.685 134.665 115.855 134.835 ;
        RECT 116.145 134.665 116.315 134.835 ;
        RECT 116.605 134.665 116.775 134.835 ;
        RECT 117.065 134.665 117.235 134.835 ;
        RECT 117.525 134.665 117.695 134.835 ;
        RECT 117.985 134.665 118.155 134.835 ;
        RECT 118.445 134.665 118.615 134.835 ;
        RECT 118.905 134.665 119.075 134.835 ;
        RECT 119.365 134.665 119.535 134.835 ;
        RECT 119.825 134.665 119.995 134.835 ;
        RECT 120.285 134.665 120.455 134.835 ;
        RECT 120.745 134.665 120.915 134.835 ;
        RECT 121.205 134.665 121.375 134.835 ;
        RECT 121.665 134.665 121.835 134.835 ;
        RECT 122.125 134.665 122.295 134.835 ;
        RECT 122.585 134.665 122.755 134.835 ;
        RECT 123.045 134.665 123.215 134.835 ;
        RECT 123.505 134.665 123.675 134.835 ;
        RECT 123.965 134.665 124.135 134.835 ;
        RECT 124.425 134.665 124.595 134.835 ;
        RECT 124.885 134.665 125.055 134.835 ;
        RECT 125.345 134.665 125.515 134.835 ;
        RECT 125.805 134.665 125.975 134.835 ;
        RECT 126.265 134.665 126.435 134.835 ;
        RECT 126.725 134.665 126.895 134.835 ;
        RECT 127.185 134.665 127.355 134.835 ;
        RECT 127.645 134.665 127.815 134.835 ;
        RECT 128.105 134.665 128.275 134.835 ;
        RECT 128.565 134.665 128.735 134.835 ;
        RECT 129.025 134.665 129.195 134.835 ;
        RECT 129.485 134.665 129.655 134.835 ;
        RECT 129.945 134.665 130.115 134.835 ;
        RECT 130.405 134.665 130.575 134.835 ;
        RECT 130.865 134.665 131.035 134.835 ;
        RECT 131.325 134.665 131.495 134.835 ;
        RECT 131.785 134.665 131.955 134.835 ;
        RECT 132.245 134.665 132.415 134.835 ;
        RECT 132.705 134.665 132.875 134.835 ;
        RECT 133.165 134.665 133.335 134.835 ;
        RECT 133.625 134.665 133.795 134.835 ;
        RECT 134.085 134.665 134.255 134.835 ;
        RECT 134.545 134.665 134.715 134.835 ;
        RECT 135.005 134.665 135.175 134.835 ;
        RECT 135.465 134.665 135.635 134.835 ;
        RECT 135.925 134.665 136.095 134.835 ;
        RECT 136.385 134.665 136.555 134.835 ;
        RECT 136.845 134.665 137.015 134.835 ;
        RECT 137.305 134.665 137.475 134.835 ;
        RECT 137.765 134.665 137.935 134.835 ;
        RECT 138.225 134.665 138.395 134.835 ;
        RECT 138.685 134.665 138.855 134.835 ;
        RECT 139.145 134.665 139.315 134.835 ;
        RECT 139.605 134.665 139.775 134.835 ;
        RECT 140.065 134.665 140.235 134.835 ;
        RECT 140.525 134.665 140.695 134.835 ;
        RECT 140.985 134.665 141.155 134.835 ;
        RECT 141.445 134.665 141.615 134.835 ;
        RECT 141.905 134.665 142.075 134.835 ;
        RECT 142.365 134.665 142.535 134.835 ;
        RECT 142.825 134.665 142.995 134.835 ;
        RECT 143.285 134.665 143.455 134.835 ;
        RECT 143.745 134.665 143.915 134.835 ;
        RECT 144.205 134.665 144.375 134.835 ;
        RECT 144.665 134.665 144.835 134.835 ;
        RECT 145.125 134.665 145.295 134.835 ;
        RECT 145.585 134.665 145.755 134.835 ;
        RECT 146.045 134.665 146.215 134.835 ;
        RECT 146.505 134.665 146.675 134.835 ;
        RECT 146.965 134.665 147.135 134.835 ;
        RECT 147.425 134.665 147.595 134.835 ;
        RECT 147.885 134.665 148.055 134.835 ;
        RECT 148.345 134.665 148.515 134.835 ;
        RECT 148.805 134.665 148.975 134.835 ;
        RECT 149.265 134.665 149.435 134.835 ;
        RECT 149.725 134.665 149.895 134.835 ;
        RECT 150.185 134.665 150.355 134.835 ;
        RECT 31.965 134.155 32.135 134.325 ;
        RECT 32.425 133.475 32.595 133.645 ;
        RECT 35.645 133.475 35.815 133.645 ;
        RECT 36.565 133.525 36.735 133.695 ;
        RECT 36.105 132.795 36.275 132.965 ;
        RECT 38.865 133.475 39.035 133.645 ;
        RECT 39.325 133.475 39.495 133.645 ;
        RECT 39.785 133.475 39.955 133.645 ;
        RECT 40.705 133.475 40.875 133.645 ;
        RECT 41.625 133.475 41.795 133.645 ;
        RECT 42.545 133.475 42.715 133.645 ;
        RECT 37.485 132.455 37.655 132.625 ;
        RECT 42.545 132.455 42.715 132.625 ;
        RECT 43.005 133.135 43.175 133.305 ;
        RECT 44.845 133.475 45.015 133.645 ;
        RECT 44.385 133.135 44.555 133.305 ;
        RECT 46.685 133.815 46.855 133.985 ;
        RECT 46.225 133.475 46.395 133.645 ;
        RECT 47.605 133.475 47.775 133.645 ;
        RECT 54.505 134.155 54.675 134.325 ;
        RECT 52.205 133.475 52.375 133.645 ;
        RECT 48.525 132.455 48.695 132.625 ;
        RECT 53.125 132.455 53.295 132.625 ;
        RECT 65.545 133.475 65.715 133.645 ;
        RECT 66.465 133.475 66.635 133.645 ;
        RECT 66.005 132.455 66.175 132.625 ;
        RECT 68.765 133.475 68.935 133.645 ;
        RECT 70.145 133.475 70.315 133.645 ;
        RECT 67.845 132.455 68.015 132.625 ;
        RECT 69.685 133.135 69.855 133.305 ;
        RECT 104.185 134.155 104.355 134.325 ;
        RECT 102.345 133.475 102.515 133.645 ;
        RECT 102.805 133.135 102.975 133.305 ;
        RECT 105.105 133.815 105.275 133.985 ;
        RECT 104.645 133.475 104.815 133.645 ;
        RECT 107.405 133.815 107.575 133.985 ;
        RECT 106.485 133.475 106.655 133.645 ;
        RECT 107.865 133.475 108.035 133.645 ;
        RECT 108.325 133.475 108.495 133.645 ;
        RECT 110.165 133.475 110.335 133.645 ;
        RECT 110.625 133.475 110.795 133.645 ;
        RECT 111.545 133.475 111.715 133.645 ;
        RECT 109.245 132.795 109.415 132.965 ;
        RECT 112.005 133.475 112.175 133.645 ;
        RECT 112.925 132.455 113.095 132.625 ;
        RECT 11.265 131.945 11.435 132.115 ;
        RECT 11.725 131.945 11.895 132.115 ;
        RECT 12.185 131.945 12.355 132.115 ;
        RECT 12.645 131.945 12.815 132.115 ;
        RECT 13.105 131.945 13.275 132.115 ;
        RECT 13.565 131.945 13.735 132.115 ;
        RECT 14.025 131.945 14.195 132.115 ;
        RECT 14.485 131.945 14.655 132.115 ;
        RECT 14.945 131.945 15.115 132.115 ;
        RECT 15.405 131.945 15.575 132.115 ;
        RECT 15.865 131.945 16.035 132.115 ;
        RECT 16.325 131.945 16.495 132.115 ;
        RECT 16.785 131.945 16.955 132.115 ;
        RECT 17.245 131.945 17.415 132.115 ;
        RECT 17.705 131.945 17.875 132.115 ;
        RECT 18.165 131.945 18.335 132.115 ;
        RECT 18.625 131.945 18.795 132.115 ;
        RECT 19.085 131.945 19.255 132.115 ;
        RECT 19.545 131.945 19.715 132.115 ;
        RECT 20.005 131.945 20.175 132.115 ;
        RECT 20.465 131.945 20.635 132.115 ;
        RECT 20.925 131.945 21.095 132.115 ;
        RECT 21.385 131.945 21.555 132.115 ;
        RECT 21.845 131.945 22.015 132.115 ;
        RECT 22.305 131.945 22.475 132.115 ;
        RECT 22.765 131.945 22.935 132.115 ;
        RECT 23.225 131.945 23.395 132.115 ;
        RECT 23.685 131.945 23.855 132.115 ;
        RECT 24.145 131.945 24.315 132.115 ;
        RECT 24.605 131.945 24.775 132.115 ;
        RECT 25.065 131.945 25.235 132.115 ;
        RECT 25.525 131.945 25.695 132.115 ;
        RECT 25.985 131.945 26.155 132.115 ;
        RECT 26.445 131.945 26.615 132.115 ;
        RECT 26.905 131.945 27.075 132.115 ;
        RECT 27.365 131.945 27.535 132.115 ;
        RECT 27.825 131.945 27.995 132.115 ;
        RECT 28.285 131.945 28.455 132.115 ;
        RECT 28.745 131.945 28.915 132.115 ;
        RECT 29.205 131.945 29.375 132.115 ;
        RECT 29.665 131.945 29.835 132.115 ;
        RECT 30.125 131.945 30.295 132.115 ;
        RECT 30.585 131.945 30.755 132.115 ;
        RECT 31.045 131.945 31.215 132.115 ;
        RECT 31.505 131.945 31.675 132.115 ;
        RECT 31.965 131.945 32.135 132.115 ;
        RECT 32.425 131.945 32.595 132.115 ;
        RECT 32.885 131.945 33.055 132.115 ;
        RECT 33.345 131.945 33.515 132.115 ;
        RECT 33.805 131.945 33.975 132.115 ;
        RECT 34.265 131.945 34.435 132.115 ;
        RECT 34.725 131.945 34.895 132.115 ;
        RECT 35.185 131.945 35.355 132.115 ;
        RECT 35.645 131.945 35.815 132.115 ;
        RECT 36.105 131.945 36.275 132.115 ;
        RECT 36.565 131.945 36.735 132.115 ;
        RECT 37.025 131.945 37.195 132.115 ;
        RECT 37.485 131.945 37.655 132.115 ;
        RECT 37.945 131.945 38.115 132.115 ;
        RECT 38.405 131.945 38.575 132.115 ;
        RECT 38.865 131.945 39.035 132.115 ;
        RECT 39.325 131.945 39.495 132.115 ;
        RECT 39.785 131.945 39.955 132.115 ;
        RECT 40.245 131.945 40.415 132.115 ;
        RECT 40.705 131.945 40.875 132.115 ;
        RECT 41.165 131.945 41.335 132.115 ;
        RECT 41.625 131.945 41.795 132.115 ;
        RECT 42.085 131.945 42.255 132.115 ;
        RECT 42.545 131.945 42.715 132.115 ;
        RECT 43.005 131.945 43.175 132.115 ;
        RECT 43.465 131.945 43.635 132.115 ;
        RECT 43.925 131.945 44.095 132.115 ;
        RECT 44.385 131.945 44.555 132.115 ;
        RECT 44.845 131.945 45.015 132.115 ;
        RECT 45.305 131.945 45.475 132.115 ;
        RECT 45.765 131.945 45.935 132.115 ;
        RECT 46.225 131.945 46.395 132.115 ;
        RECT 46.685 131.945 46.855 132.115 ;
        RECT 47.145 131.945 47.315 132.115 ;
        RECT 47.605 131.945 47.775 132.115 ;
        RECT 48.065 131.945 48.235 132.115 ;
        RECT 48.525 131.945 48.695 132.115 ;
        RECT 48.985 131.945 49.155 132.115 ;
        RECT 49.445 131.945 49.615 132.115 ;
        RECT 49.905 131.945 50.075 132.115 ;
        RECT 50.365 131.945 50.535 132.115 ;
        RECT 50.825 131.945 50.995 132.115 ;
        RECT 51.285 131.945 51.455 132.115 ;
        RECT 51.745 131.945 51.915 132.115 ;
        RECT 52.205 131.945 52.375 132.115 ;
        RECT 52.665 131.945 52.835 132.115 ;
        RECT 53.125 131.945 53.295 132.115 ;
        RECT 53.585 131.945 53.755 132.115 ;
        RECT 54.045 131.945 54.215 132.115 ;
        RECT 54.505 131.945 54.675 132.115 ;
        RECT 54.965 131.945 55.135 132.115 ;
        RECT 55.425 131.945 55.595 132.115 ;
        RECT 55.885 131.945 56.055 132.115 ;
        RECT 56.345 131.945 56.515 132.115 ;
        RECT 56.805 131.945 56.975 132.115 ;
        RECT 57.265 131.945 57.435 132.115 ;
        RECT 57.725 131.945 57.895 132.115 ;
        RECT 58.185 131.945 58.355 132.115 ;
        RECT 58.645 131.945 58.815 132.115 ;
        RECT 59.105 131.945 59.275 132.115 ;
        RECT 59.565 131.945 59.735 132.115 ;
        RECT 60.025 131.945 60.195 132.115 ;
        RECT 60.485 131.945 60.655 132.115 ;
        RECT 60.945 131.945 61.115 132.115 ;
        RECT 61.405 131.945 61.575 132.115 ;
        RECT 61.865 131.945 62.035 132.115 ;
        RECT 62.325 131.945 62.495 132.115 ;
        RECT 62.785 131.945 62.955 132.115 ;
        RECT 63.245 131.945 63.415 132.115 ;
        RECT 63.705 131.945 63.875 132.115 ;
        RECT 64.165 131.945 64.335 132.115 ;
        RECT 64.625 131.945 64.795 132.115 ;
        RECT 65.085 131.945 65.255 132.115 ;
        RECT 65.545 131.945 65.715 132.115 ;
        RECT 66.005 131.945 66.175 132.115 ;
        RECT 66.465 131.945 66.635 132.115 ;
        RECT 66.925 131.945 67.095 132.115 ;
        RECT 67.385 131.945 67.555 132.115 ;
        RECT 67.845 131.945 68.015 132.115 ;
        RECT 68.305 131.945 68.475 132.115 ;
        RECT 68.765 131.945 68.935 132.115 ;
        RECT 69.225 131.945 69.395 132.115 ;
        RECT 69.685 131.945 69.855 132.115 ;
        RECT 70.145 131.945 70.315 132.115 ;
        RECT 70.605 131.945 70.775 132.115 ;
        RECT 71.065 131.945 71.235 132.115 ;
        RECT 71.525 131.945 71.695 132.115 ;
        RECT 71.985 131.945 72.155 132.115 ;
        RECT 72.445 131.945 72.615 132.115 ;
        RECT 72.905 131.945 73.075 132.115 ;
        RECT 73.365 131.945 73.535 132.115 ;
        RECT 73.825 131.945 73.995 132.115 ;
        RECT 74.285 131.945 74.455 132.115 ;
        RECT 74.745 131.945 74.915 132.115 ;
        RECT 75.205 131.945 75.375 132.115 ;
        RECT 75.665 131.945 75.835 132.115 ;
        RECT 76.125 131.945 76.295 132.115 ;
        RECT 76.585 131.945 76.755 132.115 ;
        RECT 77.045 131.945 77.215 132.115 ;
        RECT 77.505 131.945 77.675 132.115 ;
        RECT 77.965 131.945 78.135 132.115 ;
        RECT 78.425 131.945 78.595 132.115 ;
        RECT 78.885 131.945 79.055 132.115 ;
        RECT 79.345 131.945 79.515 132.115 ;
        RECT 79.805 131.945 79.975 132.115 ;
        RECT 80.265 131.945 80.435 132.115 ;
        RECT 80.725 131.945 80.895 132.115 ;
        RECT 81.185 131.945 81.355 132.115 ;
        RECT 81.645 131.945 81.815 132.115 ;
        RECT 82.105 131.945 82.275 132.115 ;
        RECT 82.565 131.945 82.735 132.115 ;
        RECT 83.025 131.945 83.195 132.115 ;
        RECT 83.485 131.945 83.655 132.115 ;
        RECT 83.945 131.945 84.115 132.115 ;
        RECT 84.405 131.945 84.575 132.115 ;
        RECT 84.865 131.945 85.035 132.115 ;
        RECT 85.325 131.945 85.495 132.115 ;
        RECT 85.785 131.945 85.955 132.115 ;
        RECT 86.245 131.945 86.415 132.115 ;
        RECT 86.705 131.945 86.875 132.115 ;
        RECT 87.165 131.945 87.335 132.115 ;
        RECT 87.625 131.945 87.795 132.115 ;
        RECT 88.085 131.945 88.255 132.115 ;
        RECT 88.545 131.945 88.715 132.115 ;
        RECT 89.005 131.945 89.175 132.115 ;
        RECT 89.465 131.945 89.635 132.115 ;
        RECT 89.925 131.945 90.095 132.115 ;
        RECT 90.385 131.945 90.555 132.115 ;
        RECT 90.845 131.945 91.015 132.115 ;
        RECT 91.305 131.945 91.475 132.115 ;
        RECT 91.765 131.945 91.935 132.115 ;
        RECT 92.225 131.945 92.395 132.115 ;
        RECT 92.685 131.945 92.855 132.115 ;
        RECT 93.145 131.945 93.315 132.115 ;
        RECT 93.605 131.945 93.775 132.115 ;
        RECT 94.065 131.945 94.235 132.115 ;
        RECT 94.525 131.945 94.695 132.115 ;
        RECT 94.985 131.945 95.155 132.115 ;
        RECT 95.445 131.945 95.615 132.115 ;
        RECT 95.905 131.945 96.075 132.115 ;
        RECT 96.365 131.945 96.535 132.115 ;
        RECT 96.825 131.945 96.995 132.115 ;
        RECT 97.285 131.945 97.455 132.115 ;
        RECT 97.745 131.945 97.915 132.115 ;
        RECT 98.205 131.945 98.375 132.115 ;
        RECT 98.665 131.945 98.835 132.115 ;
        RECT 99.125 131.945 99.295 132.115 ;
        RECT 99.585 131.945 99.755 132.115 ;
        RECT 100.045 131.945 100.215 132.115 ;
        RECT 100.505 131.945 100.675 132.115 ;
        RECT 100.965 131.945 101.135 132.115 ;
        RECT 101.425 131.945 101.595 132.115 ;
        RECT 101.885 131.945 102.055 132.115 ;
        RECT 102.345 131.945 102.515 132.115 ;
        RECT 102.805 131.945 102.975 132.115 ;
        RECT 103.265 131.945 103.435 132.115 ;
        RECT 103.725 131.945 103.895 132.115 ;
        RECT 104.185 131.945 104.355 132.115 ;
        RECT 104.645 131.945 104.815 132.115 ;
        RECT 105.105 131.945 105.275 132.115 ;
        RECT 105.565 131.945 105.735 132.115 ;
        RECT 106.025 131.945 106.195 132.115 ;
        RECT 106.485 131.945 106.655 132.115 ;
        RECT 106.945 131.945 107.115 132.115 ;
        RECT 107.405 131.945 107.575 132.115 ;
        RECT 107.865 131.945 108.035 132.115 ;
        RECT 108.325 131.945 108.495 132.115 ;
        RECT 108.785 131.945 108.955 132.115 ;
        RECT 109.245 131.945 109.415 132.115 ;
        RECT 109.705 131.945 109.875 132.115 ;
        RECT 110.165 131.945 110.335 132.115 ;
        RECT 110.625 131.945 110.795 132.115 ;
        RECT 111.085 131.945 111.255 132.115 ;
        RECT 111.545 131.945 111.715 132.115 ;
        RECT 112.005 131.945 112.175 132.115 ;
        RECT 112.465 131.945 112.635 132.115 ;
        RECT 112.925 131.945 113.095 132.115 ;
        RECT 113.385 131.945 113.555 132.115 ;
        RECT 113.845 131.945 114.015 132.115 ;
        RECT 114.305 131.945 114.475 132.115 ;
        RECT 114.765 131.945 114.935 132.115 ;
        RECT 115.225 131.945 115.395 132.115 ;
        RECT 115.685 131.945 115.855 132.115 ;
        RECT 116.145 131.945 116.315 132.115 ;
        RECT 116.605 131.945 116.775 132.115 ;
        RECT 117.065 131.945 117.235 132.115 ;
        RECT 117.525 131.945 117.695 132.115 ;
        RECT 117.985 131.945 118.155 132.115 ;
        RECT 118.445 131.945 118.615 132.115 ;
        RECT 118.905 131.945 119.075 132.115 ;
        RECT 119.365 131.945 119.535 132.115 ;
        RECT 119.825 131.945 119.995 132.115 ;
        RECT 120.285 131.945 120.455 132.115 ;
        RECT 120.745 131.945 120.915 132.115 ;
        RECT 121.205 131.945 121.375 132.115 ;
        RECT 121.665 131.945 121.835 132.115 ;
        RECT 122.125 131.945 122.295 132.115 ;
        RECT 122.585 131.945 122.755 132.115 ;
        RECT 123.045 131.945 123.215 132.115 ;
        RECT 123.505 131.945 123.675 132.115 ;
        RECT 123.965 131.945 124.135 132.115 ;
        RECT 124.425 131.945 124.595 132.115 ;
        RECT 124.885 131.945 125.055 132.115 ;
        RECT 125.345 131.945 125.515 132.115 ;
        RECT 125.805 131.945 125.975 132.115 ;
        RECT 126.265 131.945 126.435 132.115 ;
        RECT 126.725 131.945 126.895 132.115 ;
        RECT 127.185 131.945 127.355 132.115 ;
        RECT 127.645 131.945 127.815 132.115 ;
        RECT 128.105 131.945 128.275 132.115 ;
        RECT 128.565 131.945 128.735 132.115 ;
        RECT 129.025 131.945 129.195 132.115 ;
        RECT 129.485 131.945 129.655 132.115 ;
        RECT 129.945 131.945 130.115 132.115 ;
        RECT 130.405 131.945 130.575 132.115 ;
        RECT 130.865 131.945 131.035 132.115 ;
        RECT 131.325 131.945 131.495 132.115 ;
        RECT 131.785 131.945 131.955 132.115 ;
        RECT 132.245 131.945 132.415 132.115 ;
        RECT 132.705 131.945 132.875 132.115 ;
        RECT 133.165 131.945 133.335 132.115 ;
        RECT 133.625 131.945 133.795 132.115 ;
        RECT 134.085 131.945 134.255 132.115 ;
        RECT 134.545 131.945 134.715 132.115 ;
        RECT 135.005 131.945 135.175 132.115 ;
        RECT 135.465 131.945 135.635 132.115 ;
        RECT 135.925 131.945 136.095 132.115 ;
        RECT 136.385 131.945 136.555 132.115 ;
        RECT 136.845 131.945 137.015 132.115 ;
        RECT 137.305 131.945 137.475 132.115 ;
        RECT 137.765 131.945 137.935 132.115 ;
        RECT 138.225 131.945 138.395 132.115 ;
        RECT 138.685 131.945 138.855 132.115 ;
        RECT 139.145 131.945 139.315 132.115 ;
        RECT 139.605 131.945 139.775 132.115 ;
        RECT 140.065 131.945 140.235 132.115 ;
        RECT 140.525 131.945 140.695 132.115 ;
        RECT 140.985 131.945 141.155 132.115 ;
        RECT 141.445 131.945 141.615 132.115 ;
        RECT 141.905 131.945 142.075 132.115 ;
        RECT 142.365 131.945 142.535 132.115 ;
        RECT 142.825 131.945 142.995 132.115 ;
        RECT 143.285 131.945 143.455 132.115 ;
        RECT 143.745 131.945 143.915 132.115 ;
        RECT 144.205 131.945 144.375 132.115 ;
        RECT 144.665 131.945 144.835 132.115 ;
        RECT 145.125 131.945 145.295 132.115 ;
        RECT 145.585 131.945 145.755 132.115 ;
        RECT 146.045 131.945 146.215 132.115 ;
        RECT 146.505 131.945 146.675 132.115 ;
        RECT 146.965 131.945 147.135 132.115 ;
        RECT 147.425 131.945 147.595 132.115 ;
        RECT 147.885 131.945 148.055 132.115 ;
        RECT 148.345 131.945 148.515 132.115 ;
        RECT 148.805 131.945 148.975 132.115 ;
        RECT 149.265 131.945 149.435 132.115 ;
        RECT 149.725 131.945 149.895 132.115 ;
        RECT 150.185 131.945 150.355 132.115 ;
        RECT 27.365 131.435 27.535 131.605 ;
        RECT 29.675 130.755 29.845 130.925 ;
        RECT 30.110 131.095 30.280 131.265 ;
        RECT 31.680 131.095 31.850 131.265 ;
        RECT 32.195 130.755 32.365 130.925 ;
        RECT 32.985 130.415 33.155 130.585 ;
        RECT 33.385 130.755 33.555 130.925 ;
        RECT 33.780 131.095 33.950 131.265 ;
        RECT 34.265 130.415 34.435 130.585 ;
        RECT 44.385 131.095 44.555 131.265 ;
        RECT 43.005 130.415 43.175 130.585 ;
        RECT 44.845 130.415 45.015 130.585 ;
        RECT 42.085 129.735 42.255 129.905 ;
        RECT 52.665 131.435 52.835 131.605 ;
        RECT 52.665 130.415 52.835 130.585 ;
        RECT 54.045 130.415 54.215 130.585 ;
        RECT 53.585 130.075 53.755 130.245 ;
        RECT 55.425 130.755 55.595 130.925 ;
        RECT 55.885 130.755 56.055 130.925 ;
        RECT 56.345 130.415 56.515 130.585 ;
        RECT 56.805 130.415 56.975 130.585 ;
        RECT 60.485 131.435 60.655 131.605 ;
        RECT 60.025 130.755 60.195 130.925 ;
        RECT 58.645 130.415 58.815 130.585 ;
        RECT 54.505 129.735 54.675 129.905 ;
        RECT 61.405 129.735 61.575 129.905 ;
        RECT 68.305 130.075 68.475 130.245 ;
        RECT 69.225 130.415 69.395 130.585 ;
        RECT 73.825 131.095 73.995 131.265 ;
        RECT 67.385 129.735 67.555 129.905 ;
        RECT 73.825 130.075 73.995 130.245 ;
        RECT 74.745 130.415 74.915 130.585 ;
        RECT 75.205 130.415 75.375 130.585 ;
        RECT 78.885 131.095 79.055 131.265 ;
        RECT 76.750 130.415 76.920 130.585 ;
        RECT 76.125 129.735 76.295 129.905 ;
        RECT 79.345 130.755 79.515 130.925 ;
        RECT 80.725 130.415 80.895 130.585 ;
        RECT 81.645 129.735 81.815 129.905 ;
        RECT 83.485 131.095 83.655 131.265 ;
        RECT 84.405 130.415 84.575 130.585 ;
        RECT 84.865 130.075 85.035 130.245 ;
        RECT 85.325 129.735 85.495 129.905 ;
        RECT 86.705 130.415 86.875 130.585 ;
        RECT 86.245 129.735 86.415 129.905 ;
        RECT 87.625 130.075 87.795 130.245 ;
        RECT 88.085 130.415 88.255 130.585 ;
        RECT 88.545 130.415 88.715 130.585 ;
        RECT 100.505 131.095 100.675 131.265 ;
        RECT 89.465 129.735 89.635 129.905 ;
        RECT 99.125 130.755 99.295 130.925 ;
        RECT 98.665 130.415 98.835 130.585 ;
        RECT 107.405 131.095 107.575 131.265 ;
        RECT 109.715 130.755 109.885 130.925 ;
        RECT 110.150 131.095 110.320 131.265 ;
        RECT 111.720 131.095 111.890 131.265 ;
        RECT 112.235 130.755 112.405 130.925 ;
        RECT 112.970 130.415 113.140 130.585 ;
        RECT 113.425 130.755 113.595 130.925 ;
        RECT 113.820 131.095 113.990 131.265 ;
        RECT 114.305 130.755 114.475 130.925 ;
        RECT 11.265 129.225 11.435 129.395 ;
        RECT 11.725 129.225 11.895 129.395 ;
        RECT 12.185 129.225 12.355 129.395 ;
        RECT 12.645 129.225 12.815 129.395 ;
        RECT 13.105 129.225 13.275 129.395 ;
        RECT 13.565 129.225 13.735 129.395 ;
        RECT 14.025 129.225 14.195 129.395 ;
        RECT 14.485 129.225 14.655 129.395 ;
        RECT 14.945 129.225 15.115 129.395 ;
        RECT 15.405 129.225 15.575 129.395 ;
        RECT 15.865 129.225 16.035 129.395 ;
        RECT 16.325 129.225 16.495 129.395 ;
        RECT 16.785 129.225 16.955 129.395 ;
        RECT 17.245 129.225 17.415 129.395 ;
        RECT 17.705 129.225 17.875 129.395 ;
        RECT 18.165 129.225 18.335 129.395 ;
        RECT 18.625 129.225 18.795 129.395 ;
        RECT 19.085 129.225 19.255 129.395 ;
        RECT 19.545 129.225 19.715 129.395 ;
        RECT 20.005 129.225 20.175 129.395 ;
        RECT 20.465 129.225 20.635 129.395 ;
        RECT 20.925 129.225 21.095 129.395 ;
        RECT 21.385 129.225 21.555 129.395 ;
        RECT 21.845 129.225 22.015 129.395 ;
        RECT 22.305 129.225 22.475 129.395 ;
        RECT 22.765 129.225 22.935 129.395 ;
        RECT 23.225 129.225 23.395 129.395 ;
        RECT 23.685 129.225 23.855 129.395 ;
        RECT 24.145 129.225 24.315 129.395 ;
        RECT 24.605 129.225 24.775 129.395 ;
        RECT 25.065 129.225 25.235 129.395 ;
        RECT 25.525 129.225 25.695 129.395 ;
        RECT 25.985 129.225 26.155 129.395 ;
        RECT 26.445 129.225 26.615 129.395 ;
        RECT 26.905 129.225 27.075 129.395 ;
        RECT 27.365 129.225 27.535 129.395 ;
        RECT 27.825 129.225 27.995 129.395 ;
        RECT 28.285 129.225 28.455 129.395 ;
        RECT 28.745 129.225 28.915 129.395 ;
        RECT 29.205 129.225 29.375 129.395 ;
        RECT 29.665 129.225 29.835 129.395 ;
        RECT 30.125 129.225 30.295 129.395 ;
        RECT 30.585 129.225 30.755 129.395 ;
        RECT 31.045 129.225 31.215 129.395 ;
        RECT 31.505 129.225 31.675 129.395 ;
        RECT 31.965 129.225 32.135 129.395 ;
        RECT 32.425 129.225 32.595 129.395 ;
        RECT 32.885 129.225 33.055 129.395 ;
        RECT 33.345 129.225 33.515 129.395 ;
        RECT 33.805 129.225 33.975 129.395 ;
        RECT 34.265 129.225 34.435 129.395 ;
        RECT 34.725 129.225 34.895 129.395 ;
        RECT 35.185 129.225 35.355 129.395 ;
        RECT 35.645 129.225 35.815 129.395 ;
        RECT 36.105 129.225 36.275 129.395 ;
        RECT 36.565 129.225 36.735 129.395 ;
        RECT 37.025 129.225 37.195 129.395 ;
        RECT 37.485 129.225 37.655 129.395 ;
        RECT 37.945 129.225 38.115 129.395 ;
        RECT 38.405 129.225 38.575 129.395 ;
        RECT 38.865 129.225 39.035 129.395 ;
        RECT 39.325 129.225 39.495 129.395 ;
        RECT 39.785 129.225 39.955 129.395 ;
        RECT 40.245 129.225 40.415 129.395 ;
        RECT 40.705 129.225 40.875 129.395 ;
        RECT 41.165 129.225 41.335 129.395 ;
        RECT 41.625 129.225 41.795 129.395 ;
        RECT 42.085 129.225 42.255 129.395 ;
        RECT 42.545 129.225 42.715 129.395 ;
        RECT 43.005 129.225 43.175 129.395 ;
        RECT 43.465 129.225 43.635 129.395 ;
        RECT 43.925 129.225 44.095 129.395 ;
        RECT 44.385 129.225 44.555 129.395 ;
        RECT 44.845 129.225 45.015 129.395 ;
        RECT 45.305 129.225 45.475 129.395 ;
        RECT 45.765 129.225 45.935 129.395 ;
        RECT 46.225 129.225 46.395 129.395 ;
        RECT 46.685 129.225 46.855 129.395 ;
        RECT 47.145 129.225 47.315 129.395 ;
        RECT 47.605 129.225 47.775 129.395 ;
        RECT 48.065 129.225 48.235 129.395 ;
        RECT 48.525 129.225 48.695 129.395 ;
        RECT 48.985 129.225 49.155 129.395 ;
        RECT 49.445 129.225 49.615 129.395 ;
        RECT 49.905 129.225 50.075 129.395 ;
        RECT 50.365 129.225 50.535 129.395 ;
        RECT 50.825 129.225 50.995 129.395 ;
        RECT 51.285 129.225 51.455 129.395 ;
        RECT 51.745 129.225 51.915 129.395 ;
        RECT 52.205 129.225 52.375 129.395 ;
        RECT 52.665 129.225 52.835 129.395 ;
        RECT 53.125 129.225 53.295 129.395 ;
        RECT 53.585 129.225 53.755 129.395 ;
        RECT 54.045 129.225 54.215 129.395 ;
        RECT 54.505 129.225 54.675 129.395 ;
        RECT 54.965 129.225 55.135 129.395 ;
        RECT 55.425 129.225 55.595 129.395 ;
        RECT 55.885 129.225 56.055 129.395 ;
        RECT 56.345 129.225 56.515 129.395 ;
        RECT 56.805 129.225 56.975 129.395 ;
        RECT 57.265 129.225 57.435 129.395 ;
        RECT 57.725 129.225 57.895 129.395 ;
        RECT 58.185 129.225 58.355 129.395 ;
        RECT 58.645 129.225 58.815 129.395 ;
        RECT 59.105 129.225 59.275 129.395 ;
        RECT 59.565 129.225 59.735 129.395 ;
        RECT 60.025 129.225 60.195 129.395 ;
        RECT 60.485 129.225 60.655 129.395 ;
        RECT 60.945 129.225 61.115 129.395 ;
        RECT 61.405 129.225 61.575 129.395 ;
        RECT 61.865 129.225 62.035 129.395 ;
        RECT 62.325 129.225 62.495 129.395 ;
        RECT 62.785 129.225 62.955 129.395 ;
        RECT 63.245 129.225 63.415 129.395 ;
        RECT 63.705 129.225 63.875 129.395 ;
        RECT 64.165 129.225 64.335 129.395 ;
        RECT 64.625 129.225 64.795 129.395 ;
        RECT 65.085 129.225 65.255 129.395 ;
        RECT 65.545 129.225 65.715 129.395 ;
        RECT 66.005 129.225 66.175 129.395 ;
        RECT 66.465 129.225 66.635 129.395 ;
        RECT 66.925 129.225 67.095 129.395 ;
        RECT 67.385 129.225 67.555 129.395 ;
        RECT 67.845 129.225 68.015 129.395 ;
        RECT 68.305 129.225 68.475 129.395 ;
        RECT 68.765 129.225 68.935 129.395 ;
        RECT 69.225 129.225 69.395 129.395 ;
        RECT 69.685 129.225 69.855 129.395 ;
        RECT 70.145 129.225 70.315 129.395 ;
        RECT 70.605 129.225 70.775 129.395 ;
        RECT 71.065 129.225 71.235 129.395 ;
        RECT 71.525 129.225 71.695 129.395 ;
        RECT 71.985 129.225 72.155 129.395 ;
        RECT 72.445 129.225 72.615 129.395 ;
        RECT 72.905 129.225 73.075 129.395 ;
        RECT 73.365 129.225 73.535 129.395 ;
        RECT 73.825 129.225 73.995 129.395 ;
        RECT 74.285 129.225 74.455 129.395 ;
        RECT 74.745 129.225 74.915 129.395 ;
        RECT 75.205 129.225 75.375 129.395 ;
        RECT 75.665 129.225 75.835 129.395 ;
        RECT 76.125 129.225 76.295 129.395 ;
        RECT 76.585 129.225 76.755 129.395 ;
        RECT 77.045 129.225 77.215 129.395 ;
        RECT 77.505 129.225 77.675 129.395 ;
        RECT 77.965 129.225 78.135 129.395 ;
        RECT 78.425 129.225 78.595 129.395 ;
        RECT 78.885 129.225 79.055 129.395 ;
        RECT 79.345 129.225 79.515 129.395 ;
        RECT 79.805 129.225 79.975 129.395 ;
        RECT 80.265 129.225 80.435 129.395 ;
        RECT 80.725 129.225 80.895 129.395 ;
        RECT 81.185 129.225 81.355 129.395 ;
        RECT 81.645 129.225 81.815 129.395 ;
        RECT 82.105 129.225 82.275 129.395 ;
        RECT 82.565 129.225 82.735 129.395 ;
        RECT 83.025 129.225 83.195 129.395 ;
        RECT 83.485 129.225 83.655 129.395 ;
        RECT 83.945 129.225 84.115 129.395 ;
        RECT 84.405 129.225 84.575 129.395 ;
        RECT 84.865 129.225 85.035 129.395 ;
        RECT 85.325 129.225 85.495 129.395 ;
        RECT 85.785 129.225 85.955 129.395 ;
        RECT 86.245 129.225 86.415 129.395 ;
        RECT 86.705 129.225 86.875 129.395 ;
        RECT 87.165 129.225 87.335 129.395 ;
        RECT 87.625 129.225 87.795 129.395 ;
        RECT 88.085 129.225 88.255 129.395 ;
        RECT 88.545 129.225 88.715 129.395 ;
        RECT 89.005 129.225 89.175 129.395 ;
        RECT 89.465 129.225 89.635 129.395 ;
        RECT 89.925 129.225 90.095 129.395 ;
        RECT 90.385 129.225 90.555 129.395 ;
        RECT 90.845 129.225 91.015 129.395 ;
        RECT 91.305 129.225 91.475 129.395 ;
        RECT 91.765 129.225 91.935 129.395 ;
        RECT 92.225 129.225 92.395 129.395 ;
        RECT 92.685 129.225 92.855 129.395 ;
        RECT 93.145 129.225 93.315 129.395 ;
        RECT 93.605 129.225 93.775 129.395 ;
        RECT 94.065 129.225 94.235 129.395 ;
        RECT 94.525 129.225 94.695 129.395 ;
        RECT 94.985 129.225 95.155 129.395 ;
        RECT 95.445 129.225 95.615 129.395 ;
        RECT 95.905 129.225 96.075 129.395 ;
        RECT 96.365 129.225 96.535 129.395 ;
        RECT 96.825 129.225 96.995 129.395 ;
        RECT 97.285 129.225 97.455 129.395 ;
        RECT 97.745 129.225 97.915 129.395 ;
        RECT 98.205 129.225 98.375 129.395 ;
        RECT 98.665 129.225 98.835 129.395 ;
        RECT 99.125 129.225 99.295 129.395 ;
        RECT 99.585 129.225 99.755 129.395 ;
        RECT 100.045 129.225 100.215 129.395 ;
        RECT 100.505 129.225 100.675 129.395 ;
        RECT 100.965 129.225 101.135 129.395 ;
        RECT 101.425 129.225 101.595 129.395 ;
        RECT 101.885 129.225 102.055 129.395 ;
        RECT 102.345 129.225 102.515 129.395 ;
        RECT 102.805 129.225 102.975 129.395 ;
        RECT 103.265 129.225 103.435 129.395 ;
        RECT 103.725 129.225 103.895 129.395 ;
        RECT 104.185 129.225 104.355 129.395 ;
        RECT 104.645 129.225 104.815 129.395 ;
        RECT 105.105 129.225 105.275 129.395 ;
        RECT 105.565 129.225 105.735 129.395 ;
        RECT 106.025 129.225 106.195 129.395 ;
        RECT 106.485 129.225 106.655 129.395 ;
        RECT 106.945 129.225 107.115 129.395 ;
        RECT 107.405 129.225 107.575 129.395 ;
        RECT 107.865 129.225 108.035 129.395 ;
        RECT 108.325 129.225 108.495 129.395 ;
        RECT 108.785 129.225 108.955 129.395 ;
        RECT 109.245 129.225 109.415 129.395 ;
        RECT 109.705 129.225 109.875 129.395 ;
        RECT 110.165 129.225 110.335 129.395 ;
        RECT 110.625 129.225 110.795 129.395 ;
        RECT 111.085 129.225 111.255 129.395 ;
        RECT 111.545 129.225 111.715 129.395 ;
        RECT 112.005 129.225 112.175 129.395 ;
        RECT 112.465 129.225 112.635 129.395 ;
        RECT 112.925 129.225 113.095 129.395 ;
        RECT 113.385 129.225 113.555 129.395 ;
        RECT 113.845 129.225 114.015 129.395 ;
        RECT 114.305 129.225 114.475 129.395 ;
        RECT 114.765 129.225 114.935 129.395 ;
        RECT 115.225 129.225 115.395 129.395 ;
        RECT 115.685 129.225 115.855 129.395 ;
        RECT 116.145 129.225 116.315 129.395 ;
        RECT 116.605 129.225 116.775 129.395 ;
        RECT 117.065 129.225 117.235 129.395 ;
        RECT 117.525 129.225 117.695 129.395 ;
        RECT 117.985 129.225 118.155 129.395 ;
        RECT 118.445 129.225 118.615 129.395 ;
        RECT 118.905 129.225 119.075 129.395 ;
        RECT 119.365 129.225 119.535 129.395 ;
        RECT 119.825 129.225 119.995 129.395 ;
        RECT 120.285 129.225 120.455 129.395 ;
        RECT 120.745 129.225 120.915 129.395 ;
        RECT 121.205 129.225 121.375 129.395 ;
        RECT 121.665 129.225 121.835 129.395 ;
        RECT 122.125 129.225 122.295 129.395 ;
        RECT 122.585 129.225 122.755 129.395 ;
        RECT 123.045 129.225 123.215 129.395 ;
        RECT 123.505 129.225 123.675 129.395 ;
        RECT 123.965 129.225 124.135 129.395 ;
        RECT 124.425 129.225 124.595 129.395 ;
        RECT 124.885 129.225 125.055 129.395 ;
        RECT 125.345 129.225 125.515 129.395 ;
        RECT 125.805 129.225 125.975 129.395 ;
        RECT 126.265 129.225 126.435 129.395 ;
        RECT 126.725 129.225 126.895 129.395 ;
        RECT 127.185 129.225 127.355 129.395 ;
        RECT 127.645 129.225 127.815 129.395 ;
        RECT 128.105 129.225 128.275 129.395 ;
        RECT 128.565 129.225 128.735 129.395 ;
        RECT 129.025 129.225 129.195 129.395 ;
        RECT 129.485 129.225 129.655 129.395 ;
        RECT 129.945 129.225 130.115 129.395 ;
        RECT 130.405 129.225 130.575 129.395 ;
        RECT 130.865 129.225 131.035 129.395 ;
        RECT 131.325 129.225 131.495 129.395 ;
        RECT 131.785 129.225 131.955 129.395 ;
        RECT 132.245 129.225 132.415 129.395 ;
        RECT 132.705 129.225 132.875 129.395 ;
        RECT 133.165 129.225 133.335 129.395 ;
        RECT 133.625 129.225 133.795 129.395 ;
        RECT 134.085 129.225 134.255 129.395 ;
        RECT 134.545 129.225 134.715 129.395 ;
        RECT 135.005 129.225 135.175 129.395 ;
        RECT 135.465 129.225 135.635 129.395 ;
        RECT 135.925 129.225 136.095 129.395 ;
        RECT 136.385 129.225 136.555 129.395 ;
        RECT 136.845 129.225 137.015 129.395 ;
        RECT 137.305 129.225 137.475 129.395 ;
        RECT 137.765 129.225 137.935 129.395 ;
        RECT 138.225 129.225 138.395 129.395 ;
        RECT 138.685 129.225 138.855 129.395 ;
        RECT 139.145 129.225 139.315 129.395 ;
        RECT 139.605 129.225 139.775 129.395 ;
        RECT 140.065 129.225 140.235 129.395 ;
        RECT 140.525 129.225 140.695 129.395 ;
        RECT 140.985 129.225 141.155 129.395 ;
        RECT 141.445 129.225 141.615 129.395 ;
        RECT 141.905 129.225 142.075 129.395 ;
        RECT 142.365 129.225 142.535 129.395 ;
        RECT 142.825 129.225 142.995 129.395 ;
        RECT 143.285 129.225 143.455 129.395 ;
        RECT 143.745 129.225 143.915 129.395 ;
        RECT 144.205 129.225 144.375 129.395 ;
        RECT 144.665 129.225 144.835 129.395 ;
        RECT 145.125 129.225 145.295 129.395 ;
        RECT 145.585 129.225 145.755 129.395 ;
        RECT 146.045 129.225 146.215 129.395 ;
        RECT 146.505 129.225 146.675 129.395 ;
        RECT 146.965 129.225 147.135 129.395 ;
        RECT 147.425 129.225 147.595 129.395 ;
        RECT 147.885 129.225 148.055 129.395 ;
        RECT 148.345 129.225 148.515 129.395 ;
        RECT 148.805 129.225 148.975 129.395 ;
        RECT 149.265 129.225 149.435 129.395 ;
        RECT 149.725 129.225 149.895 129.395 ;
        RECT 150.185 129.225 150.355 129.395 ;
        RECT 42.085 128.035 42.255 128.205 ;
        RECT 43.005 128.035 43.175 128.205 ;
        RECT 43.925 128.035 44.095 128.205 ;
        RECT 44.385 128.035 44.555 128.205 ;
        RECT 48.985 128.035 49.155 128.205 ;
        RECT 49.905 128.035 50.075 128.205 ;
        RECT 45.305 127.015 45.475 127.185 ;
        RECT 49.445 127.695 49.615 127.865 ;
        RECT 51.730 128.035 51.900 128.205 ;
        RECT 50.825 127.355 50.995 127.525 ;
        RECT 53.585 127.695 53.755 127.865 ;
        RECT 59.105 128.375 59.275 128.545 ;
        RECT 54.045 127.695 54.215 127.865 ;
        RECT 60.025 128.715 60.195 128.885 ;
        RECT 61.405 128.715 61.575 128.885 ;
        RECT 60.485 128.035 60.655 128.205 ;
        RECT 60.945 128.035 61.115 128.205 ;
        RECT 61.865 128.035 62.035 128.205 ;
        RECT 63.245 128.035 63.415 128.205 ;
        RECT 59.105 127.015 59.275 127.185 ;
        RECT 66.925 128.035 67.095 128.205 ;
        RECT 67.410 127.355 67.580 127.525 ;
        RECT 67.805 127.695 67.975 127.865 ;
        RECT 68.205 128.035 68.375 128.205 ;
        RECT 68.995 127.695 69.165 127.865 ;
        RECT 69.510 127.355 69.680 127.525 ;
        RECT 71.080 127.355 71.250 127.525 ;
        RECT 71.515 127.695 71.685 127.865 ;
        RECT 73.825 128.715 73.995 128.885 ;
        RECT 75.665 128.715 75.835 128.885 ;
        RECT 77.505 128.035 77.675 128.205 ;
        RECT 77.045 127.695 77.215 127.865 ;
        RECT 84.405 128.715 84.575 128.885 ;
        RECT 81.645 128.375 81.815 128.545 ;
        RECT 81.185 128.035 81.355 128.205 ;
        RECT 82.105 128.035 82.275 128.205 ;
        RECT 82.565 128.035 82.735 128.205 ;
        RECT 83.485 128.035 83.655 128.205 ;
        RECT 86.245 128.035 86.415 128.205 ;
        RECT 88.085 128.035 88.255 128.205 ;
        RECT 89.005 128.035 89.175 128.205 ;
        RECT 89.465 128.035 89.635 128.205 ;
        RECT 85.325 127.355 85.495 127.525 ;
        RECT 87.625 127.015 87.795 127.185 ;
        RECT 90.385 128.375 90.555 128.545 ;
        RECT 90.385 127.355 90.555 127.525 ;
        RECT 91.305 127.015 91.475 127.185 ;
        RECT 93.615 127.695 93.785 127.865 ;
        RECT 94.050 127.355 94.220 127.525 ;
        RECT 96.135 127.695 96.305 127.865 ;
        RECT 95.620 127.355 95.790 127.525 ;
        RECT 96.870 128.035 97.040 128.205 ;
        RECT 97.325 127.695 97.495 127.865 ;
        RECT 98.205 128.035 98.375 128.205 ;
        RECT 97.720 127.355 97.890 127.525 ;
        RECT 11.265 126.505 11.435 126.675 ;
        RECT 11.725 126.505 11.895 126.675 ;
        RECT 12.185 126.505 12.355 126.675 ;
        RECT 12.645 126.505 12.815 126.675 ;
        RECT 13.105 126.505 13.275 126.675 ;
        RECT 13.565 126.505 13.735 126.675 ;
        RECT 14.025 126.505 14.195 126.675 ;
        RECT 14.485 126.505 14.655 126.675 ;
        RECT 14.945 126.505 15.115 126.675 ;
        RECT 15.405 126.505 15.575 126.675 ;
        RECT 15.865 126.505 16.035 126.675 ;
        RECT 16.325 126.505 16.495 126.675 ;
        RECT 16.785 126.505 16.955 126.675 ;
        RECT 17.245 126.505 17.415 126.675 ;
        RECT 17.705 126.505 17.875 126.675 ;
        RECT 18.165 126.505 18.335 126.675 ;
        RECT 18.625 126.505 18.795 126.675 ;
        RECT 19.085 126.505 19.255 126.675 ;
        RECT 19.545 126.505 19.715 126.675 ;
        RECT 20.005 126.505 20.175 126.675 ;
        RECT 20.465 126.505 20.635 126.675 ;
        RECT 20.925 126.505 21.095 126.675 ;
        RECT 21.385 126.505 21.555 126.675 ;
        RECT 21.845 126.505 22.015 126.675 ;
        RECT 22.305 126.505 22.475 126.675 ;
        RECT 22.765 126.505 22.935 126.675 ;
        RECT 23.225 126.505 23.395 126.675 ;
        RECT 23.685 126.505 23.855 126.675 ;
        RECT 24.145 126.505 24.315 126.675 ;
        RECT 24.605 126.505 24.775 126.675 ;
        RECT 25.065 126.505 25.235 126.675 ;
        RECT 25.525 126.505 25.695 126.675 ;
        RECT 25.985 126.505 26.155 126.675 ;
        RECT 26.445 126.505 26.615 126.675 ;
        RECT 26.905 126.505 27.075 126.675 ;
        RECT 27.365 126.505 27.535 126.675 ;
        RECT 27.825 126.505 27.995 126.675 ;
        RECT 28.285 126.505 28.455 126.675 ;
        RECT 28.745 126.505 28.915 126.675 ;
        RECT 29.205 126.505 29.375 126.675 ;
        RECT 29.665 126.505 29.835 126.675 ;
        RECT 30.125 126.505 30.295 126.675 ;
        RECT 30.585 126.505 30.755 126.675 ;
        RECT 31.045 126.505 31.215 126.675 ;
        RECT 31.505 126.505 31.675 126.675 ;
        RECT 31.965 126.505 32.135 126.675 ;
        RECT 32.425 126.505 32.595 126.675 ;
        RECT 32.885 126.505 33.055 126.675 ;
        RECT 33.345 126.505 33.515 126.675 ;
        RECT 33.805 126.505 33.975 126.675 ;
        RECT 34.265 126.505 34.435 126.675 ;
        RECT 34.725 126.505 34.895 126.675 ;
        RECT 35.185 126.505 35.355 126.675 ;
        RECT 35.645 126.505 35.815 126.675 ;
        RECT 36.105 126.505 36.275 126.675 ;
        RECT 36.565 126.505 36.735 126.675 ;
        RECT 37.025 126.505 37.195 126.675 ;
        RECT 37.485 126.505 37.655 126.675 ;
        RECT 37.945 126.505 38.115 126.675 ;
        RECT 38.405 126.505 38.575 126.675 ;
        RECT 38.865 126.505 39.035 126.675 ;
        RECT 39.325 126.505 39.495 126.675 ;
        RECT 39.785 126.505 39.955 126.675 ;
        RECT 40.245 126.505 40.415 126.675 ;
        RECT 40.705 126.505 40.875 126.675 ;
        RECT 41.165 126.505 41.335 126.675 ;
        RECT 41.625 126.505 41.795 126.675 ;
        RECT 42.085 126.505 42.255 126.675 ;
        RECT 42.545 126.505 42.715 126.675 ;
        RECT 43.005 126.505 43.175 126.675 ;
        RECT 43.465 126.505 43.635 126.675 ;
        RECT 43.925 126.505 44.095 126.675 ;
        RECT 44.385 126.505 44.555 126.675 ;
        RECT 44.845 126.505 45.015 126.675 ;
        RECT 45.305 126.505 45.475 126.675 ;
        RECT 45.765 126.505 45.935 126.675 ;
        RECT 46.225 126.505 46.395 126.675 ;
        RECT 46.685 126.505 46.855 126.675 ;
        RECT 47.145 126.505 47.315 126.675 ;
        RECT 47.605 126.505 47.775 126.675 ;
        RECT 48.065 126.505 48.235 126.675 ;
        RECT 48.525 126.505 48.695 126.675 ;
        RECT 48.985 126.505 49.155 126.675 ;
        RECT 49.445 126.505 49.615 126.675 ;
        RECT 49.905 126.505 50.075 126.675 ;
        RECT 50.365 126.505 50.535 126.675 ;
        RECT 50.825 126.505 50.995 126.675 ;
        RECT 51.285 126.505 51.455 126.675 ;
        RECT 51.745 126.505 51.915 126.675 ;
        RECT 52.205 126.505 52.375 126.675 ;
        RECT 52.665 126.505 52.835 126.675 ;
        RECT 53.125 126.505 53.295 126.675 ;
        RECT 53.585 126.505 53.755 126.675 ;
        RECT 54.045 126.505 54.215 126.675 ;
        RECT 54.505 126.505 54.675 126.675 ;
        RECT 54.965 126.505 55.135 126.675 ;
        RECT 55.425 126.505 55.595 126.675 ;
        RECT 55.885 126.505 56.055 126.675 ;
        RECT 56.345 126.505 56.515 126.675 ;
        RECT 56.805 126.505 56.975 126.675 ;
        RECT 57.265 126.505 57.435 126.675 ;
        RECT 57.725 126.505 57.895 126.675 ;
        RECT 58.185 126.505 58.355 126.675 ;
        RECT 58.645 126.505 58.815 126.675 ;
        RECT 59.105 126.505 59.275 126.675 ;
        RECT 59.565 126.505 59.735 126.675 ;
        RECT 60.025 126.505 60.195 126.675 ;
        RECT 60.485 126.505 60.655 126.675 ;
        RECT 60.945 126.505 61.115 126.675 ;
        RECT 61.405 126.505 61.575 126.675 ;
        RECT 61.865 126.505 62.035 126.675 ;
        RECT 62.325 126.505 62.495 126.675 ;
        RECT 62.785 126.505 62.955 126.675 ;
        RECT 63.245 126.505 63.415 126.675 ;
        RECT 63.705 126.505 63.875 126.675 ;
        RECT 64.165 126.505 64.335 126.675 ;
        RECT 64.625 126.505 64.795 126.675 ;
        RECT 65.085 126.505 65.255 126.675 ;
        RECT 65.545 126.505 65.715 126.675 ;
        RECT 66.005 126.505 66.175 126.675 ;
        RECT 66.465 126.505 66.635 126.675 ;
        RECT 66.925 126.505 67.095 126.675 ;
        RECT 67.385 126.505 67.555 126.675 ;
        RECT 67.845 126.505 68.015 126.675 ;
        RECT 68.305 126.505 68.475 126.675 ;
        RECT 68.765 126.505 68.935 126.675 ;
        RECT 69.225 126.505 69.395 126.675 ;
        RECT 69.685 126.505 69.855 126.675 ;
        RECT 70.145 126.505 70.315 126.675 ;
        RECT 70.605 126.505 70.775 126.675 ;
        RECT 71.065 126.505 71.235 126.675 ;
        RECT 71.525 126.505 71.695 126.675 ;
        RECT 71.985 126.505 72.155 126.675 ;
        RECT 72.445 126.505 72.615 126.675 ;
        RECT 72.905 126.505 73.075 126.675 ;
        RECT 73.365 126.505 73.535 126.675 ;
        RECT 73.825 126.505 73.995 126.675 ;
        RECT 74.285 126.505 74.455 126.675 ;
        RECT 74.745 126.505 74.915 126.675 ;
        RECT 75.205 126.505 75.375 126.675 ;
        RECT 75.665 126.505 75.835 126.675 ;
        RECT 76.125 126.505 76.295 126.675 ;
        RECT 76.585 126.505 76.755 126.675 ;
        RECT 77.045 126.505 77.215 126.675 ;
        RECT 77.505 126.505 77.675 126.675 ;
        RECT 77.965 126.505 78.135 126.675 ;
        RECT 78.425 126.505 78.595 126.675 ;
        RECT 78.885 126.505 79.055 126.675 ;
        RECT 79.345 126.505 79.515 126.675 ;
        RECT 79.805 126.505 79.975 126.675 ;
        RECT 80.265 126.505 80.435 126.675 ;
        RECT 80.725 126.505 80.895 126.675 ;
        RECT 81.185 126.505 81.355 126.675 ;
        RECT 81.645 126.505 81.815 126.675 ;
        RECT 82.105 126.505 82.275 126.675 ;
        RECT 82.565 126.505 82.735 126.675 ;
        RECT 83.025 126.505 83.195 126.675 ;
        RECT 83.485 126.505 83.655 126.675 ;
        RECT 83.945 126.505 84.115 126.675 ;
        RECT 84.405 126.505 84.575 126.675 ;
        RECT 84.865 126.505 85.035 126.675 ;
        RECT 85.325 126.505 85.495 126.675 ;
        RECT 85.785 126.505 85.955 126.675 ;
        RECT 86.245 126.505 86.415 126.675 ;
        RECT 86.705 126.505 86.875 126.675 ;
        RECT 87.165 126.505 87.335 126.675 ;
        RECT 87.625 126.505 87.795 126.675 ;
        RECT 88.085 126.505 88.255 126.675 ;
        RECT 88.545 126.505 88.715 126.675 ;
        RECT 89.005 126.505 89.175 126.675 ;
        RECT 89.465 126.505 89.635 126.675 ;
        RECT 89.925 126.505 90.095 126.675 ;
        RECT 90.385 126.505 90.555 126.675 ;
        RECT 90.845 126.505 91.015 126.675 ;
        RECT 91.305 126.505 91.475 126.675 ;
        RECT 91.765 126.505 91.935 126.675 ;
        RECT 92.225 126.505 92.395 126.675 ;
        RECT 92.685 126.505 92.855 126.675 ;
        RECT 93.145 126.505 93.315 126.675 ;
        RECT 93.605 126.505 93.775 126.675 ;
        RECT 94.065 126.505 94.235 126.675 ;
        RECT 94.525 126.505 94.695 126.675 ;
        RECT 94.985 126.505 95.155 126.675 ;
        RECT 95.445 126.505 95.615 126.675 ;
        RECT 95.905 126.505 96.075 126.675 ;
        RECT 96.365 126.505 96.535 126.675 ;
        RECT 96.825 126.505 96.995 126.675 ;
        RECT 97.285 126.505 97.455 126.675 ;
        RECT 97.745 126.505 97.915 126.675 ;
        RECT 98.205 126.505 98.375 126.675 ;
        RECT 98.665 126.505 98.835 126.675 ;
        RECT 99.125 126.505 99.295 126.675 ;
        RECT 99.585 126.505 99.755 126.675 ;
        RECT 100.045 126.505 100.215 126.675 ;
        RECT 100.505 126.505 100.675 126.675 ;
        RECT 100.965 126.505 101.135 126.675 ;
        RECT 101.425 126.505 101.595 126.675 ;
        RECT 101.885 126.505 102.055 126.675 ;
        RECT 102.345 126.505 102.515 126.675 ;
        RECT 102.805 126.505 102.975 126.675 ;
        RECT 103.265 126.505 103.435 126.675 ;
        RECT 103.725 126.505 103.895 126.675 ;
        RECT 104.185 126.505 104.355 126.675 ;
        RECT 104.645 126.505 104.815 126.675 ;
        RECT 105.105 126.505 105.275 126.675 ;
        RECT 105.565 126.505 105.735 126.675 ;
        RECT 106.025 126.505 106.195 126.675 ;
        RECT 106.485 126.505 106.655 126.675 ;
        RECT 106.945 126.505 107.115 126.675 ;
        RECT 107.405 126.505 107.575 126.675 ;
        RECT 107.865 126.505 108.035 126.675 ;
        RECT 108.325 126.505 108.495 126.675 ;
        RECT 108.785 126.505 108.955 126.675 ;
        RECT 109.245 126.505 109.415 126.675 ;
        RECT 109.705 126.505 109.875 126.675 ;
        RECT 110.165 126.505 110.335 126.675 ;
        RECT 110.625 126.505 110.795 126.675 ;
        RECT 111.085 126.505 111.255 126.675 ;
        RECT 111.545 126.505 111.715 126.675 ;
        RECT 112.005 126.505 112.175 126.675 ;
        RECT 112.465 126.505 112.635 126.675 ;
        RECT 112.925 126.505 113.095 126.675 ;
        RECT 113.385 126.505 113.555 126.675 ;
        RECT 113.845 126.505 114.015 126.675 ;
        RECT 114.305 126.505 114.475 126.675 ;
        RECT 114.765 126.505 114.935 126.675 ;
        RECT 115.225 126.505 115.395 126.675 ;
        RECT 115.685 126.505 115.855 126.675 ;
        RECT 116.145 126.505 116.315 126.675 ;
        RECT 116.605 126.505 116.775 126.675 ;
        RECT 117.065 126.505 117.235 126.675 ;
        RECT 117.525 126.505 117.695 126.675 ;
        RECT 117.985 126.505 118.155 126.675 ;
        RECT 118.445 126.505 118.615 126.675 ;
        RECT 118.905 126.505 119.075 126.675 ;
        RECT 119.365 126.505 119.535 126.675 ;
        RECT 119.825 126.505 119.995 126.675 ;
        RECT 120.285 126.505 120.455 126.675 ;
        RECT 120.745 126.505 120.915 126.675 ;
        RECT 121.205 126.505 121.375 126.675 ;
        RECT 121.665 126.505 121.835 126.675 ;
        RECT 122.125 126.505 122.295 126.675 ;
        RECT 122.585 126.505 122.755 126.675 ;
        RECT 123.045 126.505 123.215 126.675 ;
        RECT 123.505 126.505 123.675 126.675 ;
        RECT 123.965 126.505 124.135 126.675 ;
        RECT 124.425 126.505 124.595 126.675 ;
        RECT 124.885 126.505 125.055 126.675 ;
        RECT 125.345 126.505 125.515 126.675 ;
        RECT 125.805 126.505 125.975 126.675 ;
        RECT 126.265 126.505 126.435 126.675 ;
        RECT 126.725 126.505 126.895 126.675 ;
        RECT 127.185 126.505 127.355 126.675 ;
        RECT 127.645 126.505 127.815 126.675 ;
        RECT 128.105 126.505 128.275 126.675 ;
        RECT 128.565 126.505 128.735 126.675 ;
        RECT 129.025 126.505 129.195 126.675 ;
        RECT 129.485 126.505 129.655 126.675 ;
        RECT 129.945 126.505 130.115 126.675 ;
        RECT 130.405 126.505 130.575 126.675 ;
        RECT 130.865 126.505 131.035 126.675 ;
        RECT 131.325 126.505 131.495 126.675 ;
        RECT 131.785 126.505 131.955 126.675 ;
        RECT 132.245 126.505 132.415 126.675 ;
        RECT 132.705 126.505 132.875 126.675 ;
        RECT 133.165 126.505 133.335 126.675 ;
        RECT 133.625 126.505 133.795 126.675 ;
        RECT 134.085 126.505 134.255 126.675 ;
        RECT 134.545 126.505 134.715 126.675 ;
        RECT 135.005 126.505 135.175 126.675 ;
        RECT 135.465 126.505 135.635 126.675 ;
        RECT 135.925 126.505 136.095 126.675 ;
        RECT 136.385 126.505 136.555 126.675 ;
        RECT 136.845 126.505 137.015 126.675 ;
        RECT 137.305 126.505 137.475 126.675 ;
        RECT 137.765 126.505 137.935 126.675 ;
        RECT 138.225 126.505 138.395 126.675 ;
        RECT 138.685 126.505 138.855 126.675 ;
        RECT 139.145 126.505 139.315 126.675 ;
        RECT 139.605 126.505 139.775 126.675 ;
        RECT 140.065 126.505 140.235 126.675 ;
        RECT 140.525 126.505 140.695 126.675 ;
        RECT 140.985 126.505 141.155 126.675 ;
        RECT 141.445 126.505 141.615 126.675 ;
        RECT 141.905 126.505 142.075 126.675 ;
        RECT 142.365 126.505 142.535 126.675 ;
        RECT 142.825 126.505 142.995 126.675 ;
        RECT 143.285 126.505 143.455 126.675 ;
        RECT 143.745 126.505 143.915 126.675 ;
        RECT 144.205 126.505 144.375 126.675 ;
        RECT 144.665 126.505 144.835 126.675 ;
        RECT 145.125 126.505 145.295 126.675 ;
        RECT 145.585 126.505 145.755 126.675 ;
        RECT 146.045 126.505 146.215 126.675 ;
        RECT 146.505 126.505 146.675 126.675 ;
        RECT 146.965 126.505 147.135 126.675 ;
        RECT 147.425 126.505 147.595 126.675 ;
        RECT 147.885 126.505 148.055 126.675 ;
        RECT 148.345 126.505 148.515 126.675 ;
        RECT 148.805 126.505 148.975 126.675 ;
        RECT 149.265 126.505 149.435 126.675 ;
        RECT 149.725 126.505 149.895 126.675 ;
        RECT 150.185 126.505 150.355 126.675 ;
        RECT 39.785 125.995 39.955 126.165 ;
        RECT 42.095 125.315 42.265 125.485 ;
        RECT 42.530 125.655 42.700 125.825 ;
        RECT 44.100 125.655 44.270 125.825 ;
        RECT 44.615 125.315 44.785 125.485 ;
        RECT 45.350 124.635 45.520 124.805 ;
        RECT 45.805 125.315 45.975 125.485 ;
        RECT 46.200 125.655 46.370 125.825 ;
        RECT 46.685 124.975 46.855 125.145 ;
        RECT 58.210 125.655 58.380 125.825 ;
        RECT 57.725 124.975 57.895 125.145 ;
        RECT 58.605 125.315 58.775 125.485 ;
        RECT 59.060 124.635 59.230 124.805 ;
        RECT 60.310 125.655 60.480 125.825 ;
        RECT 59.795 125.315 59.965 125.485 ;
        RECT 61.880 125.655 62.050 125.825 ;
        RECT 62.315 125.315 62.485 125.485 ;
        RECT 64.625 125.995 64.795 126.165 ;
        RECT 66.465 125.995 66.635 126.165 ;
        RECT 65.545 124.975 65.715 125.145 ;
        RECT 91.765 125.315 91.935 125.485 ;
        RECT 95.905 125.995 96.075 126.165 ;
        RECT 94.985 124.975 95.155 125.145 ;
        RECT 95.445 124.975 95.615 125.145 ;
        RECT 96.365 124.975 96.535 125.145 ;
        RECT 11.265 123.785 11.435 123.955 ;
        RECT 11.725 123.785 11.895 123.955 ;
        RECT 12.185 123.785 12.355 123.955 ;
        RECT 12.645 123.785 12.815 123.955 ;
        RECT 13.105 123.785 13.275 123.955 ;
        RECT 13.565 123.785 13.735 123.955 ;
        RECT 14.025 123.785 14.195 123.955 ;
        RECT 14.485 123.785 14.655 123.955 ;
        RECT 14.945 123.785 15.115 123.955 ;
        RECT 15.405 123.785 15.575 123.955 ;
        RECT 15.865 123.785 16.035 123.955 ;
        RECT 16.325 123.785 16.495 123.955 ;
        RECT 16.785 123.785 16.955 123.955 ;
        RECT 17.245 123.785 17.415 123.955 ;
        RECT 17.705 123.785 17.875 123.955 ;
        RECT 18.165 123.785 18.335 123.955 ;
        RECT 18.625 123.785 18.795 123.955 ;
        RECT 19.085 123.785 19.255 123.955 ;
        RECT 19.545 123.785 19.715 123.955 ;
        RECT 20.005 123.785 20.175 123.955 ;
        RECT 20.465 123.785 20.635 123.955 ;
        RECT 20.925 123.785 21.095 123.955 ;
        RECT 21.385 123.785 21.555 123.955 ;
        RECT 21.845 123.785 22.015 123.955 ;
        RECT 22.305 123.785 22.475 123.955 ;
        RECT 22.765 123.785 22.935 123.955 ;
        RECT 23.225 123.785 23.395 123.955 ;
        RECT 23.685 123.785 23.855 123.955 ;
        RECT 24.145 123.785 24.315 123.955 ;
        RECT 24.605 123.785 24.775 123.955 ;
        RECT 25.065 123.785 25.235 123.955 ;
        RECT 25.525 123.785 25.695 123.955 ;
        RECT 25.985 123.785 26.155 123.955 ;
        RECT 26.445 123.785 26.615 123.955 ;
        RECT 26.905 123.785 27.075 123.955 ;
        RECT 27.365 123.785 27.535 123.955 ;
        RECT 27.825 123.785 27.995 123.955 ;
        RECT 28.285 123.785 28.455 123.955 ;
        RECT 28.745 123.785 28.915 123.955 ;
        RECT 29.205 123.785 29.375 123.955 ;
        RECT 29.665 123.785 29.835 123.955 ;
        RECT 30.125 123.785 30.295 123.955 ;
        RECT 30.585 123.785 30.755 123.955 ;
        RECT 31.045 123.785 31.215 123.955 ;
        RECT 31.505 123.785 31.675 123.955 ;
        RECT 31.965 123.785 32.135 123.955 ;
        RECT 32.425 123.785 32.595 123.955 ;
        RECT 32.885 123.785 33.055 123.955 ;
        RECT 33.345 123.785 33.515 123.955 ;
        RECT 33.805 123.785 33.975 123.955 ;
        RECT 34.265 123.785 34.435 123.955 ;
        RECT 34.725 123.785 34.895 123.955 ;
        RECT 35.185 123.785 35.355 123.955 ;
        RECT 35.645 123.785 35.815 123.955 ;
        RECT 36.105 123.785 36.275 123.955 ;
        RECT 36.565 123.785 36.735 123.955 ;
        RECT 37.025 123.785 37.195 123.955 ;
        RECT 37.485 123.785 37.655 123.955 ;
        RECT 37.945 123.785 38.115 123.955 ;
        RECT 38.405 123.785 38.575 123.955 ;
        RECT 38.865 123.785 39.035 123.955 ;
        RECT 39.325 123.785 39.495 123.955 ;
        RECT 39.785 123.785 39.955 123.955 ;
        RECT 40.245 123.785 40.415 123.955 ;
        RECT 40.705 123.785 40.875 123.955 ;
        RECT 41.165 123.785 41.335 123.955 ;
        RECT 41.625 123.785 41.795 123.955 ;
        RECT 42.085 123.785 42.255 123.955 ;
        RECT 42.545 123.785 42.715 123.955 ;
        RECT 43.005 123.785 43.175 123.955 ;
        RECT 43.465 123.785 43.635 123.955 ;
        RECT 43.925 123.785 44.095 123.955 ;
        RECT 44.385 123.785 44.555 123.955 ;
        RECT 44.845 123.785 45.015 123.955 ;
        RECT 45.305 123.785 45.475 123.955 ;
        RECT 45.765 123.785 45.935 123.955 ;
        RECT 46.225 123.785 46.395 123.955 ;
        RECT 46.685 123.785 46.855 123.955 ;
        RECT 47.145 123.785 47.315 123.955 ;
        RECT 47.605 123.785 47.775 123.955 ;
        RECT 48.065 123.785 48.235 123.955 ;
        RECT 48.525 123.785 48.695 123.955 ;
        RECT 48.985 123.785 49.155 123.955 ;
        RECT 49.445 123.785 49.615 123.955 ;
        RECT 49.905 123.785 50.075 123.955 ;
        RECT 50.365 123.785 50.535 123.955 ;
        RECT 50.825 123.785 50.995 123.955 ;
        RECT 51.285 123.785 51.455 123.955 ;
        RECT 51.745 123.785 51.915 123.955 ;
        RECT 52.205 123.785 52.375 123.955 ;
        RECT 52.665 123.785 52.835 123.955 ;
        RECT 53.125 123.785 53.295 123.955 ;
        RECT 53.585 123.785 53.755 123.955 ;
        RECT 54.045 123.785 54.215 123.955 ;
        RECT 54.505 123.785 54.675 123.955 ;
        RECT 54.965 123.785 55.135 123.955 ;
        RECT 55.425 123.785 55.595 123.955 ;
        RECT 55.885 123.785 56.055 123.955 ;
        RECT 56.345 123.785 56.515 123.955 ;
        RECT 56.805 123.785 56.975 123.955 ;
        RECT 57.265 123.785 57.435 123.955 ;
        RECT 57.725 123.785 57.895 123.955 ;
        RECT 58.185 123.785 58.355 123.955 ;
        RECT 58.645 123.785 58.815 123.955 ;
        RECT 59.105 123.785 59.275 123.955 ;
        RECT 59.565 123.785 59.735 123.955 ;
        RECT 60.025 123.785 60.195 123.955 ;
        RECT 60.485 123.785 60.655 123.955 ;
        RECT 60.945 123.785 61.115 123.955 ;
        RECT 61.405 123.785 61.575 123.955 ;
        RECT 61.865 123.785 62.035 123.955 ;
        RECT 62.325 123.785 62.495 123.955 ;
        RECT 62.785 123.785 62.955 123.955 ;
        RECT 63.245 123.785 63.415 123.955 ;
        RECT 63.705 123.785 63.875 123.955 ;
        RECT 64.165 123.785 64.335 123.955 ;
        RECT 64.625 123.785 64.795 123.955 ;
        RECT 65.085 123.785 65.255 123.955 ;
        RECT 65.545 123.785 65.715 123.955 ;
        RECT 66.005 123.785 66.175 123.955 ;
        RECT 66.465 123.785 66.635 123.955 ;
        RECT 66.925 123.785 67.095 123.955 ;
        RECT 67.385 123.785 67.555 123.955 ;
        RECT 67.845 123.785 68.015 123.955 ;
        RECT 68.305 123.785 68.475 123.955 ;
        RECT 68.765 123.785 68.935 123.955 ;
        RECT 69.225 123.785 69.395 123.955 ;
        RECT 69.685 123.785 69.855 123.955 ;
        RECT 70.145 123.785 70.315 123.955 ;
        RECT 70.605 123.785 70.775 123.955 ;
        RECT 71.065 123.785 71.235 123.955 ;
        RECT 71.525 123.785 71.695 123.955 ;
        RECT 71.985 123.785 72.155 123.955 ;
        RECT 72.445 123.785 72.615 123.955 ;
        RECT 72.905 123.785 73.075 123.955 ;
        RECT 73.365 123.785 73.535 123.955 ;
        RECT 73.825 123.785 73.995 123.955 ;
        RECT 74.285 123.785 74.455 123.955 ;
        RECT 74.745 123.785 74.915 123.955 ;
        RECT 75.205 123.785 75.375 123.955 ;
        RECT 75.665 123.785 75.835 123.955 ;
        RECT 76.125 123.785 76.295 123.955 ;
        RECT 76.585 123.785 76.755 123.955 ;
        RECT 77.045 123.785 77.215 123.955 ;
        RECT 77.505 123.785 77.675 123.955 ;
        RECT 77.965 123.785 78.135 123.955 ;
        RECT 78.425 123.785 78.595 123.955 ;
        RECT 78.885 123.785 79.055 123.955 ;
        RECT 79.345 123.785 79.515 123.955 ;
        RECT 79.805 123.785 79.975 123.955 ;
        RECT 80.265 123.785 80.435 123.955 ;
        RECT 80.725 123.785 80.895 123.955 ;
        RECT 81.185 123.785 81.355 123.955 ;
        RECT 81.645 123.785 81.815 123.955 ;
        RECT 82.105 123.785 82.275 123.955 ;
        RECT 82.565 123.785 82.735 123.955 ;
        RECT 83.025 123.785 83.195 123.955 ;
        RECT 83.485 123.785 83.655 123.955 ;
        RECT 83.945 123.785 84.115 123.955 ;
        RECT 84.405 123.785 84.575 123.955 ;
        RECT 84.865 123.785 85.035 123.955 ;
        RECT 85.325 123.785 85.495 123.955 ;
        RECT 85.785 123.785 85.955 123.955 ;
        RECT 86.245 123.785 86.415 123.955 ;
        RECT 86.705 123.785 86.875 123.955 ;
        RECT 87.165 123.785 87.335 123.955 ;
        RECT 87.625 123.785 87.795 123.955 ;
        RECT 88.085 123.785 88.255 123.955 ;
        RECT 88.545 123.785 88.715 123.955 ;
        RECT 89.005 123.785 89.175 123.955 ;
        RECT 89.465 123.785 89.635 123.955 ;
        RECT 89.925 123.785 90.095 123.955 ;
        RECT 90.385 123.785 90.555 123.955 ;
        RECT 90.845 123.785 91.015 123.955 ;
        RECT 91.305 123.785 91.475 123.955 ;
        RECT 91.765 123.785 91.935 123.955 ;
        RECT 92.225 123.785 92.395 123.955 ;
        RECT 92.685 123.785 92.855 123.955 ;
        RECT 93.145 123.785 93.315 123.955 ;
        RECT 93.605 123.785 93.775 123.955 ;
        RECT 94.065 123.785 94.235 123.955 ;
        RECT 94.525 123.785 94.695 123.955 ;
        RECT 94.985 123.785 95.155 123.955 ;
        RECT 95.445 123.785 95.615 123.955 ;
        RECT 95.905 123.785 96.075 123.955 ;
        RECT 96.365 123.785 96.535 123.955 ;
        RECT 96.825 123.785 96.995 123.955 ;
        RECT 97.285 123.785 97.455 123.955 ;
        RECT 97.745 123.785 97.915 123.955 ;
        RECT 98.205 123.785 98.375 123.955 ;
        RECT 98.665 123.785 98.835 123.955 ;
        RECT 99.125 123.785 99.295 123.955 ;
        RECT 99.585 123.785 99.755 123.955 ;
        RECT 100.045 123.785 100.215 123.955 ;
        RECT 100.505 123.785 100.675 123.955 ;
        RECT 100.965 123.785 101.135 123.955 ;
        RECT 101.425 123.785 101.595 123.955 ;
        RECT 101.885 123.785 102.055 123.955 ;
        RECT 102.345 123.785 102.515 123.955 ;
        RECT 102.805 123.785 102.975 123.955 ;
        RECT 103.265 123.785 103.435 123.955 ;
        RECT 103.725 123.785 103.895 123.955 ;
        RECT 104.185 123.785 104.355 123.955 ;
        RECT 104.645 123.785 104.815 123.955 ;
        RECT 105.105 123.785 105.275 123.955 ;
        RECT 105.565 123.785 105.735 123.955 ;
        RECT 106.025 123.785 106.195 123.955 ;
        RECT 106.485 123.785 106.655 123.955 ;
        RECT 106.945 123.785 107.115 123.955 ;
        RECT 107.405 123.785 107.575 123.955 ;
        RECT 107.865 123.785 108.035 123.955 ;
        RECT 108.325 123.785 108.495 123.955 ;
        RECT 108.785 123.785 108.955 123.955 ;
        RECT 109.245 123.785 109.415 123.955 ;
        RECT 109.705 123.785 109.875 123.955 ;
        RECT 110.165 123.785 110.335 123.955 ;
        RECT 110.625 123.785 110.795 123.955 ;
        RECT 111.085 123.785 111.255 123.955 ;
        RECT 111.545 123.785 111.715 123.955 ;
        RECT 112.005 123.785 112.175 123.955 ;
        RECT 112.465 123.785 112.635 123.955 ;
        RECT 112.925 123.785 113.095 123.955 ;
        RECT 113.385 123.785 113.555 123.955 ;
        RECT 113.845 123.785 114.015 123.955 ;
        RECT 114.305 123.785 114.475 123.955 ;
        RECT 114.765 123.785 114.935 123.955 ;
        RECT 115.225 123.785 115.395 123.955 ;
        RECT 115.685 123.785 115.855 123.955 ;
        RECT 116.145 123.785 116.315 123.955 ;
        RECT 116.605 123.785 116.775 123.955 ;
        RECT 117.065 123.785 117.235 123.955 ;
        RECT 117.525 123.785 117.695 123.955 ;
        RECT 117.985 123.785 118.155 123.955 ;
        RECT 118.445 123.785 118.615 123.955 ;
        RECT 118.905 123.785 119.075 123.955 ;
        RECT 119.365 123.785 119.535 123.955 ;
        RECT 119.825 123.785 119.995 123.955 ;
        RECT 120.285 123.785 120.455 123.955 ;
        RECT 120.745 123.785 120.915 123.955 ;
        RECT 121.205 123.785 121.375 123.955 ;
        RECT 121.665 123.785 121.835 123.955 ;
        RECT 122.125 123.785 122.295 123.955 ;
        RECT 122.585 123.785 122.755 123.955 ;
        RECT 123.045 123.785 123.215 123.955 ;
        RECT 123.505 123.785 123.675 123.955 ;
        RECT 123.965 123.785 124.135 123.955 ;
        RECT 124.425 123.785 124.595 123.955 ;
        RECT 124.885 123.785 125.055 123.955 ;
        RECT 125.345 123.785 125.515 123.955 ;
        RECT 125.805 123.785 125.975 123.955 ;
        RECT 126.265 123.785 126.435 123.955 ;
        RECT 126.725 123.785 126.895 123.955 ;
        RECT 127.185 123.785 127.355 123.955 ;
        RECT 127.645 123.785 127.815 123.955 ;
        RECT 128.105 123.785 128.275 123.955 ;
        RECT 128.565 123.785 128.735 123.955 ;
        RECT 129.025 123.785 129.195 123.955 ;
        RECT 129.485 123.785 129.655 123.955 ;
        RECT 129.945 123.785 130.115 123.955 ;
        RECT 130.405 123.785 130.575 123.955 ;
        RECT 130.865 123.785 131.035 123.955 ;
        RECT 131.325 123.785 131.495 123.955 ;
        RECT 131.785 123.785 131.955 123.955 ;
        RECT 132.245 123.785 132.415 123.955 ;
        RECT 132.705 123.785 132.875 123.955 ;
        RECT 133.165 123.785 133.335 123.955 ;
        RECT 133.625 123.785 133.795 123.955 ;
        RECT 134.085 123.785 134.255 123.955 ;
        RECT 134.545 123.785 134.715 123.955 ;
        RECT 135.005 123.785 135.175 123.955 ;
        RECT 135.465 123.785 135.635 123.955 ;
        RECT 135.925 123.785 136.095 123.955 ;
        RECT 136.385 123.785 136.555 123.955 ;
        RECT 136.845 123.785 137.015 123.955 ;
        RECT 137.305 123.785 137.475 123.955 ;
        RECT 137.765 123.785 137.935 123.955 ;
        RECT 138.225 123.785 138.395 123.955 ;
        RECT 138.685 123.785 138.855 123.955 ;
        RECT 139.145 123.785 139.315 123.955 ;
        RECT 139.605 123.785 139.775 123.955 ;
        RECT 140.065 123.785 140.235 123.955 ;
        RECT 140.525 123.785 140.695 123.955 ;
        RECT 140.985 123.785 141.155 123.955 ;
        RECT 141.445 123.785 141.615 123.955 ;
        RECT 141.905 123.785 142.075 123.955 ;
        RECT 142.365 123.785 142.535 123.955 ;
        RECT 142.825 123.785 142.995 123.955 ;
        RECT 143.285 123.785 143.455 123.955 ;
        RECT 143.745 123.785 143.915 123.955 ;
        RECT 144.205 123.785 144.375 123.955 ;
        RECT 144.665 123.785 144.835 123.955 ;
        RECT 145.125 123.785 145.295 123.955 ;
        RECT 145.585 123.785 145.755 123.955 ;
        RECT 146.045 123.785 146.215 123.955 ;
        RECT 146.505 123.785 146.675 123.955 ;
        RECT 146.965 123.785 147.135 123.955 ;
        RECT 147.425 123.785 147.595 123.955 ;
        RECT 147.885 123.785 148.055 123.955 ;
        RECT 148.345 123.785 148.515 123.955 ;
        RECT 148.805 123.785 148.975 123.955 ;
        RECT 149.265 123.785 149.435 123.955 ;
        RECT 149.725 123.785 149.895 123.955 ;
        RECT 150.185 123.785 150.355 123.955 ;
        RECT 47.605 122.595 47.775 122.765 ;
        RECT 48.090 121.915 48.260 122.085 ;
        RECT 48.485 122.255 48.655 122.425 ;
        RECT 48.940 122.935 49.110 123.105 ;
        RECT 49.675 122.255 49.845 122.425 ;
        RECT 50.190 121.915 50.360 122.085 ;
        RECT 51.760 121.915 51.930 122.085 ;
        RECT 52.195 122.255 52.365 122.425 ;
        RECT 54.505 123.275 54.675 123.445 ;
        RECT 11.265 121.065 11.435 121.235 ;
        RECT 11.725 121.065 11.895 121.235 ;
        RECT 12.185 121.065 12.355 121.235 ;
        RECT 12.645 121.065 12.815 121.235 ;
        RECT 13.105 121.065 13.275 121.235 ;
        RECT 13.565 121.065 13.735 121.235 ;
        RECT 14.025 121.065 14.195 121.235 ;
        RECT 14.485 121.065 14.655 121.235 ;
        RECT 14.945 121.065 15.115 121.235 ;
        RECT 15.405 121.065 15.575 121.235 ;
        RECT 15.865 121.065 16.035 121.235 ;
        RECT 16.325 121.065 16.495 121.235 ;
        RECT 16.785 121.065 16.955 121.235 ;
        RECT 17.245 121.065 17.415 121.235 ;
        RECT 17.705 121.065 17.875 121.235 ;
        RECT 18.165 121.065 18.335 121.235 ;
        RECT 18.625 121.065 18.795 121.235 ;
        RECT 19.085 121.065 19.255 121.235 ;
        RECT 19.545 121.065 19.715 121.235 ;
        RECT 20.005 121.065 20.175 121.235 ;
        RECT 20.465 121.065 20.635 121.235 ;
        RECT 20.925 121.065 21.095 121.235 ;
        RECT 21.385 121.065 21.555 121.235 ;
        RECT 21.845 121.065 22.015 121.235 ;
        RECT 22.305 121.065 22.475 121.235 ;
        RECT 22.765 121.065 22.935 121.235 ;
        RECT 23.225 121.065 23.395 121.235 ;
        RECT 23.685 121.065 23.855 121.235 ;
        RECT 24.145 121.065 24.315 121.235 ;
        RECT 24.605 121.065 24.775 121.235 ;
        RECT 25.065 121.065 25.235 121.235 ;
        RECT 25.525 121.065 25.695 121.235 ;
        RECT 25.985 121.065 26.155 121.235 ;
        RECT 26.445 121.065 26.615 121.235 ;
        RECT 26.905 121.065 27.075 121.235 ;
        RECT 27.365 121.065 27.535 121.235 ;
        RECT 27.825 121.065 27.995 121.235 ;
        RECT 28.285 121.065 28.455 121.235 ;
        RECT 28.745 121.065 28.915 121.235 ;
        RECT 29.205 121.065 29.375 121.235 ;
        RECT 29.665 121.065 29.835 121.235 ;
        RECT 30.125 121.065 30.295 121.235 ;
        RECT 30.585 121.065 30.755 121.235 ;
        RECT 31.045 121.065 31.215 121.235 ;
        RECT 31.505 121.065 31.675 121.235 ;
        RECT 31.965 121.065 32.135 121.235 ;
        RECT 32.425 121.065 32.595 121.235 ;
        RECT 32.885 121.065 33.055 121.235 ;
        RECT 33.345 121.065 33.515 121.235 ;
        RECT 33.805 121.065 33.975 121.235 ;
        RECT 34.265 121.065 34.435 121.235 ;
        RECT 34.725 121.065 34.895 121.235 ;
        RECT 35.185 121.065 35.355 121.235 ;
        RECT 35.645 121.065 35.815 121.235 ;
        RECT 36.105 121.065 36.275 121.235 ;
        RECT 36.565 121.065 36.735 121.235 ;
        RECT 37.025 121.065 37.195 121.235 ;
        RECT 37.485 121.065 37.655 121.235 ;
        RECT 37.945 121.065 38.115 121.235 ;
        RECT 38.405 121.065 38.575 121.235 ;
        RECT 38.865 121.065 39.035 121.235 ;
        RECT 39.325 121.065 39.495 121.235 ;
        RECT 39.785 121.065 39.955 121.235 ;
        RECT 40.245 121.065 40.415 121.235 ;
        RECT 40.705 121.065 40.875 121.235 ;
        RECT 41.165 121.065 41.335 121.235 ;
        RECT 41.625 121.065 41.795 121.235 ;
        RECT 42.085 121.065 42.255 121.235 ;
        RECT 42.545 121.065 42.715 121.235 ;
        RECT 43.005 121.065 43.175 121.235 ;
        RECT 43.465 121.065 43.635 121.235 ;
        RECT 43.925 121.065 44.095 121.235 ;
        RECT 44.385 121.065 44.555 121.235 ;
        RECT 44.845 121.065 45.015 121.235 ;
        RECT 45.305 121.065 45.475 121.235 ;
        RECT 45.765 121.065 45.935 121.235 ;
        RECT 46.225 121.065 46.395 121.235 ;
        RECT 46.685 121.065 46.855 121.235 ;
        RECT 47.145 121.065 47.315 121.235 ;
        RECT 47.605 121.065 47.775 121.235 ;
        RECT 48.065 121.065 48.235 121.235 ;
        RECT 48.525 121.065 48.695 121.235 ;
        RECT 48.985 121.065 49.155 121.235 ;
        RECT 49.445 121.065 49.615 121.235 ;
        RECT 49.905 121.065 50.075 121.235 ;
        RECT 50.365 121.065 50.535 121.235 ;
        RECT 50.825 121.065 50.995 121.235 ;
        RECT 51.285 121.065 51.455 121.235 ;
        RECT 51.745 121.065 51.915 121.235 ;
        RECT 52.205 121.065 52.375 121.235 ;
        RECT 52.665 121.065 52.835 121.235 ;
        RECT 53.125 121.065 53.295 121.235 ;
        RECT 53.585 121.065 53.755 121.235 ;
        RECT 54.045 121.065 54.215 121.235 ;
        RECT 54.505 121.065 54.675 121.235 ;
        RECT 54.965 121.065 55.135 121.235 ;
        RECT 55.425 121.065 55.595 121.235 ;
        RECT 55.885 121.065 56.055 121.235 ;
        RECT 56.345 121.065 56.515 121.235 ;
        RECT 56.805 121.065 56.975 121.235 ;
        RECT 57.265 121.065 57.435 121.235 ;
        RECT 57.725 121.065 57.895 121.235 ;
        RECT 58.185 121.065 58.355 121.235 ;
        RECT 58.645 121.065 58.815 121.235 ;
        RECT 59.105 121.065 59.275 121.235 ;
        RECT 59.565 121.065 59.735 121.235 ;
        RECT 60.025 121.065 60.195 121.235 ;
        RECT 60.485 121.065 60.655 121.235 ;
        RECT 60.945 121.065 61.115 121.235 ;
        RECT 61.405 121.065 61.575 121.235 ;
        RECT 61.865 121.065 62.035 121.235 ;
        RECT 62.325 121.065 62.495 121.235 ;
        RECT 62.785 121.065 62.955 121.235 ;
        RECT 63.245 121.065 63.415 121.235 ;
        RECT 63.705 121.065 63.875 121.235 ;
        RECT 64.165 121.065 64.335 121.235 ;
        RECT 64.625 121.065 64.795 121.235 ;
        RECT 65.085 121.065 65.255 121.235 ;
        RECT 65.545 121.065 65.715 121.235 ;
        RECT 66.005 121.065 66.175 121.235 ;
        RECT 66.465 121.065 66.635 121.235 ;
        RECT 66.925 121.065 67.095 121.235 ;
        RECT 67.385 121.065 67.555 121.235 ;
        RECT 67.845 121.065 68.015 121.235 ;
        RECT 68.305 121.065 68.475 121.235 ;
        RECT 68.765 121.065 68.935 121.235 ;
        RECT 69.225 121.065 69.395 121.235 ;
        RECT 69.685 121.065 69.855 121.235 ;
        RECT 70.145 121.065 70.315 121.235 ;
        RECT 70.605 121.065 70.775 121.235 ;
        RECT 71.065 121.065 71.235 121.235 ;
        RECT 71.525 121.065 71.695 121.235 ;
        RECT 71.985 121.065 72.155 121.235 ;
        RECT 72.445 121.065 72.615 121.235 ;
        RECT 72.905 121.065 73.075 121.235 ;
        RECT 73.365 121.065 73.535 121.235 ;
        RECT 73.825 121.065 73.995 121.235 ;
        RECT 74.285 121.065 74.455 121.235 ;
        RECT 74.745 121.065 74.915 121.235 ;
        RECT 75.205 121.065 75.375 121.235 ;
        RECT 75.665 121.065 75.835 121.235 ;
        RECT 76.125 121.065 76.295 121.235 ;
        RECT 76.585 121.065 76.755 121.235 ;
        RECT 77.045 121.065 77.215 121.235 ;
        RECT 77.505 121.065 77.675 121.235 ;
        RECT 77.965 121.065 78.135 121.235 ;
        RECT 78.425 121.065 78.595 121.235 ;
        RECT 78.885 121.065 79.055 121.235 ;
        RECT 79.345 121.065 79.515 121.235 ;
        RECT 79.805 121.065 79.975 121.235 ;
        RECT 80.265 121.065 80.435 121.235 ;
        RECT 80.725 121.065 80.895 121.235 ;
        RECT 81.185 121.065 81.355 121.235 ;
        RECT 81.645 121.065 81.815 121.235 ;
        RECT 82.105 121.065 82.275 121.235 ;
        RECT 82.565 121.065 82.735 121.235 ;
        RECT 83.025 121.065 83.195 121.235 ;
        RECT 83.485 121.065 83.655 121.235 ;
        RECT 83.945 121.065 84.115 121.235 ;
        RECT 84.405 121.065 84.575 121.235 ;
        RECT 84.865 121.065 85.035 121.235 ;
        RECT 85.325 121.065 85.495 121.235 ;
        RECT 85.785 121.065 85.955 121.235 ;
        RECT 86.245 121.065 86.415 121.235 ;
        RECT 86.705 121.065 86.875 121.235 ;
        RECT 87.165 121.065 87.335 121.235 ;
        RECT 87.625 121.065 87.795 121.235 ;
        RECT 88.085 121.065 88.255 121.235 ;
        RECT 88.545 121.065 88.715 121.235 ;
        RECT 89.005 121.065 89.175 121.235 ;
        RECT 89.465 121.065 89.635 121.235 ;
        RECT 89.925 121.065 90.095 121.235 ;
        RECT 90.385 121.065 90.555 121.235 ;
        RECT 90.845 121.065 91.015 121.235 ;
        RECT 91.305 121.065 91.475 121.235 ;
        RECT 91.765 121.065 91.935 121.235 ;
        RECT 92.225 121.065 92.395 121.235 ;
        RECT 92.685 121.065 92.855 121.235 ;
        RECT 93.145 121.065 93.315 121.235 ;
        RECT 93.605 121.065 93.775 121.235 ;
        RECT 94.065 121.065 94.235 121.235 ;
        RECT 94.525 121.065 94.695 121.235 ;
        RECT 94.985 121.065 95.155 121.235 ;
        RECT 95.445 121.065 95.615 121.235 ;
        RECT 95.905 121.065 96.075 121.235 ;
        RECT 96.365 121.065 96.535 121.235 ;
        RECT 96.825 121.065 96.995 121.235 ;
        RECT 97.285 121.065 97.455 121.235 ;
        RECT 97.745 121.065 97.915 121.235 ;
        RECT 98.205 121.065 98.375 121.235 ;
        RECT 98.665 121.065 98.835 121.235 ;
        RECT 99.125 121.065 99.295 121.235 ;
        RECT 99.585 121.065 99.755 121.235 ;
        RECT 100.045 121.065 100.215 121.235 ;
        RECT 100.505 121.065 100.675 121.235 ;
        RECT 100.965 121.065 101.135 121.235 ;
        RECT 101.425 121.065 101.595 121.235 ;
        RECT 101.885 121.065 102.055 121.235 ;
        RECT 102.345 121.065 102.515 121.235 ;
        RECT 102.805 121.065 102.975 121.235 ;
        RECT 103.265 121.065 103.435 121.235 ;
        RECT 103.725 121.065 103.895 121.235 ;
        RECT 104.185 121.065 104.355 121.235 ;
        RECT 104.645 121.065 104.815 121.235 ;
        RECT 105.105 121.065 105.275 121.235 ;
        RECT 105.565 121.065 105.735 121.235 ;
        RECT 106.025 121.065 106.195 121.235 ;
        RECT 106.485 121.065 106.655 121.235 ;
        RECT 106.945 121.065 107.115 121.235 ;
        RECT 107.405 121.065 107.575 121.235 ;
        RECT 107.865 121.065 108.035 121.235 ;
        RECT 108.325 121.065 108.495 121.235 ;
        RECT 108.785 121.065 108.955 121.235 ;
        RECT 109.245 121.065 109.415 121.235 ;
        RECT 109.705 121.065 109.875 121.235 ;
        RECT 110.165 121.065 110.335 121.235 ;
        RECT 110.625 121.065 110.795 121.235 ;
        RECT 111.085 121.065 111.255 121.235 ;
        RECT 111.545 121.065 111.715 121.235 ;
        RECT 112.005 121.065 112.175 121.235 ;
        RECT 112.465 121.065 112.635 121.235 ;
        RECT 112.925 121.065 113.095 121.235 ;
        RECT 113.385 121.065 113.555 121.235 ;
        RECT 113.845 121.065 114.015 121.235 ;
        RECT 114.305 121.065 114.475 121.235 ;
        RECT 114.765 121.065 114.935 121.235 ;
        RECT 115.225 121.065 115.395 121.235 ;
        RECT 115.685 121.065 115.855 121.235 ;
        RECT 116.145 121.065 116.315 121.235 ;
        RECT 116.605 121.065 116.775 121.235 ;
        RECT 117.065 121.065 117.235 121.235 ;
        RECT 117.525 121.065 117.695 121.235 ;
        RECT 117.985 121.065 118.155 121.235 ;
        RECT 118.445 121.065 118.615 121.235 ;
        RECT 118.905 121.065 119.075 121.235 ;
        RECT 119.365 121.065 119.535 121.235 ;
        RECT 119.825 121.065 119.995 121.235 ;
        RECT 120.285 121.065 120.455 121.235 ;
        RECT 120.745 121.065 120.915 121.235 ;
        RECT 121.205 121.065 121.375 121.235 ;
        RECT 121.665 121.065 121.835 121.235 ;
        RECT 122.125 121.065 122.295 121.235 ;
        RECT 122.585 121.065 122.755 121.235 ;
        RECT 123.045 121.065 123.215 121.235 ;
        RECT 123.505 121.065 123.675 121.235 ;
        RECT 123.965 121.065 124.135 121.235 ;
        RECT 124.425 121.065 124.595 121.235 ;
        RECT 124.885 121.065 125.055 121.235 ;
        RECT 125.345 121.065 125.515 121.235 ;
        RECT 125.805 121.065 125.975 121.235 ;
        RECT 126.265 121.065 126.435 121.235 ;
        RECT 126.725 121.065 126.895 121.235 ;
        RECT 127.185 121.065 127.355 121.235 ;
        RECT 127.645 121.065 127.815 121.235 ;
        RECT 128.105 121.065 128.275 121.235 ;
        RECT 128.565 121.065 128.735 121.235 ;
        RECT 129.025 121.065 129.195 121.235 ;
        RECT 129.485 121.065 129.655 121.235 ;
        RECT 129.945 121.065 130.115 121.235 ;
        RECT 130.405 121.065 130.575 121.235 ;
        RECT 130.865 121.065 131.035 121.235 ;
        RECT 131.325 121.065 131.495 121.235 ;
        RECT 131.785 121.065 131.955 121.235 ;
        RECT 132.245 121.065 132.415 121.235 ;
        RECT 132.705 121.065 132.875 121.235 ;
        RECT 133.165 121.065 133.335 121.235 ;
        RECT 133.625 121.065 133.795 121.235 ;
        RECT 134.085 121.065 134.255 121.235 ;
        RECT 134.545 121.065 134.715 121.235 ;
        RECT 135.005 121.065 135.175 121.235 ;
        RECT 135.465 121.065 135.635 121.235 ;
        RECT 135.925 121.065 136.095 121.235 ;
        RECT 136.385 121.065 136.555 121.235 ;
        RECT 136.845 121.065 137.015 121.235 ;
        RECT 137.305 121.065 137.475 121.235 ;
        RECT 137.765 121.065 137.935 121.235 ;
        RECT 138.225 121.065 138.395 121.235 ;
        RECT 138.685 121.065 138.855 121.235 ;
        RECT 139.145 121.065 139.315 121.235 ;
        RECT 139.605 121.065 139.775 121.235 ;
        RECT 140.065 121.065 140.235 121.235 ;
        RECT 140.525 121.065 140.695 121.235 ;
        RECT 140.985 121.065 141.155 121.235 ;
        RECT 141.445 121.065 141.615 121.235 ;
        RECT 141.905 121.065 142.075 121.235 ;
        RECT 142.365 121.065 142.535 121.235 ;
        RECT 142.825 121.065 142.995 121.235 ;
        RECT 143.285 121.065 143.455 121.235 ;
        RECT 143.745 121.065 143.915 121.235 ;
        RECT 144.205 121.065 144.375 121.235 ;
        RECT 144.665 121.065 144.835 121.235 ;
        RECT 145.125 121.065 145.295 121.235 ;
        RECT 145.585 121.065 145.755 121.235 ;
        RECT 146.045 121.065 146.215 121.235 ;
        RECT 146.505 121.065 146.675 121.235 ;
        RECT 146.965 121.065 147.135 121.235 ;
        RECT 147.425 121.065 147.595 121.235 ;
        RECT 147.885 121.065 148.055 121.235 ;
        RECT 148.345 121.065 148.515 121.235 ;
        RECT 148.805 121.065 148.975 121.235 ;
        RECT 149.265 121.065 149.435 121.235 ;
        RECT 149.725 121.065 149.895 121.235 ;
        RECT 150.185 121.065 150.355 121.235 ;
        RECT 11.265 118.345 11.435 118.515 ;
        RECT 11.725 118.345 11.895 118.515 ;
        RECT 12.185 118.345 12.355 118.515 ;
        RECT 12.645 118.345 12.815 118.515 ;
        RECT 13.105 118.345 13.275 118.515 ;
        RECT 13.565 118.345 13.735 118.515 ;
        RECT 14.025 118.345 14.195 118.515 ;
        RECT 14.485 118.345 14.655 118.515 ;
        RECT 14.945 118.345 15.115 118.515 ;
        RECT 15.405 118.345 15.575 118.515 ;
        RECT 15.865 118.345 16.035 118.515 ;
        RECT 16.325 118.345 16.495 118.515 ;
        RECT 16.785 118.345 16.955 118.515 ;
        RECT 17.245 118.345 17.415 118.515 ;
        RECT 17.705 118.345 17.875 118.515 ;
        RECT 18.165 118.345 18.335 118.515 ;
        RECT 18.625 118.345 18.795 118.515 ;
        RECT 19.085 118.345 19.255 118.515 ;
        RECT 19.545 118.345 19.715 118.515 ;
        RECT 20.005 118.345 20.175 118.515 ;
        RECT 20.465 118.345 20.635 118.515 ;
        RECT 20.925 118.345 21.095 118.515 ;
        RECT 21.385 118.345 21.555 118.515 ;
        RECT 21.845 118.345 22.015 118.515 ;
        RECT 22.305 118.345 22.475 118.515 ;
        RECT 22.765 118.345 22.935 118.515 ;
        RECT 23.225 118.345 23.395 118.515 ;
        RECT 23.685 118.345 23.855 118.515 ;
        RECT 24.145 118.345 24.315 118.515 ;
        RECT 24.605 118.345 24.775 118.515 ;
        RECT 25.065 118.345 25.235 118.515 ;
        RECT 25.525 118.345 25.695 118.515 ;
        RECT 25.985 118.345 26.155 118.515 ;
        RECT 26.445 118.345 26.615 118.515 ;
        RECT 26.905 118.345 27.075 118.515 ;
        RECT 27.365 118.345 27.535 118.515 ;
        RECT 27.825 118.345 27.995 118.515 ;
        RECT 28.285 118.345 28.455 118.515 ;
        RECT 28.745 118.345 28.915 118.515 ;
        RECT 29.205 118.345 29.375 118.515 ;
        RECT 29.665 118.345 29.835 118.515 ;
        RECT 30.125 118.345 30.295 118.515 ;
        RECT 30.585 118.345 30.755 118.515 ;
        RECT 31.045 118.345 31.215 118.515 ;
        RECT 31.505 118.345 31.675 118.515 ;
        RECT 31.965 118.345 32.135 118.515 ;
        RECT 32.425 118.345 32.595 118.515 ;
        RECT 32.885 118.345 33.055 118.515 ;
        RECT 33.345 118.345 33.515 118.515 ;
        RECT 33.805 118.345 33.975 118.515 ;
        RECT 34.265 118.345 34.435 118.515 ;
        RECT 34.725 118.345 34.895 118.515 ;
        RECT 35.185 118.345 35.355 118.515 ;
        RECT 35.645 118.345 35.815 118.515 ;
        RECT 36.105 118.345 36.275 118.515 ;
        RECT 36.565 118.345 36.735 118.515 ;
        RECT 37.025 118.345 37.195 118.515 ;
        RECT 37.485 118.345 37.655 118.515 ;
        RECT 37.945 118.345 38.115 118.515 ;
        RECT 38.405 118.345 38.575 118.515 ;
        RECT 38.865 118.345 39.035 118.515 ;
        RECT 39.325 118.345 39.495 118.515 ;
        RECT 39.785 118.345 39.955 118.515 ;
        RECT 40.245 118.345 40.415 118.515 ;
        RECT 40.705 118.345 40.875 118.515 ;
        RECT 41.165 118.345 41.335 118.515 ;
        RECT 41.625 118.345 41.795 118.515 ;
        RECT 42.085 118.345 42.255 118.515 ;
        RECT 42.545 118.345 42.715 118.515 ;
        RECT 43.005 118.345 43.175 118.515 ;
        RECT 43.465 118.345 43.635 118.515 ;
        RECT 43.925 118.345 44.095 118.515 ;
        RECT 44.385 118.345 44.555 118.515 ;
        RECT 44.845 118.345 45.015 118.515 ;
        RECT 45.305 118.345 45.475 118.515 ;
        RECT 45.765 118.345 45.935 118.515 ;
        RECT 46.225 118.345 46.395 118.515 ;
        RECT 46.685 118.345 46.855 118.515 ;
        RECT 47.145 118.345 47.315 118.515 ;
        RECT 47.605 118.345 47.775 118.515 ;
        RECT 48.065 118.345 48.235 118.515 ;
        RECT 48.525 118.345 48.695 118.515 ;
        RECT 48.985 118.345 49.155 118.515 ;
        RECT 49.445 118.345 49.615 118.515 ;
        RECT 49.905 118.345 50.075 118.515 ;
        RECT 50.365 118.345 50.535 118.515 ;
        RECT 50.825 118.345 50.995 118.515 ;
        RECT 51.285 118.345 51.455 118.515 ;
        RECT 51.745 118.345 51.915 118.515 ;
        RECT 52.205 118.345 52.375 118.515 ;
        RECT 52.665 118.345 52.835 118.515 ;
        RECT 53.125 118.345 53.295 118.515 ;
        RECT 53.585 118.345 53.755 118.515 ;
        RECT 54.045 118.345 54.215 118.515 ;
        RECT 54.505 118.345 54.675 118.515 ;
        RECT 54.965 118.345 55.135 118.515 ;
        RECT 55.425 118.345 55.595 118.515 ;
        RECT 55.885 118.345 56.055 118.515 ;
        RECT 56.345 118.345 56.515 118.515 ;
        RECT 56.805 118.345 56.975 118.515 ;
        RECT 57.265 118.345 57.435 118.515 ;
        RECT 57.725 118.345 57.895 118.515 ;
        RECT 58.185 118.345 58.355 118.515 ;
        RECT 58.645 118.345 58.815 118.515 ;
        RECT 59.105 118.345 59.275 118.515 ;
        RECT 59.565 118.345 59.735 118.515 ;
        RECT 60.025 118.345 60.195 118.515 ;
        RECT 60.485 118.345 60.655 118.515 ;
        RECT 60.945 118.345 61.115 118.515 ;
        RECT 61.405 118.345 61.575 118.515 ;
        RECT 61.865 118.345 62.035 118.515 ;
        RECT 62.325 118.345 62.495 118.515 ;
        RECT 62.785 118.345 62.955 118.515 ;
        RECT 63.245 118.345 63.415 118.515 ;
        RECT 63.705 118.345 63.875 118.515 ;
        RECT 64.165 118.345 64.335 118.515 ;
        RECT 64.625 118.345 64.795 118.515 ;
        RECT 65.085 118.345 65.255 118.515 ;
        RECT 65.545 118.345 65.715 118.515 ;
        RECT 66.005 118.345 66.175 118.515 ;
        RECT 66.465 118.345 66.635 118.515 ;
        RECT 66.925 118.345 67.095 118.515 ;
        RECT 67.385 118.345 67.555 118.515 ;
        RECT 67.845 118.345 68.015 118.515 ;
        RECT 68.305 118.345 68.475 118.515 ;
        RECT 68.765 118.345 68.935 118.515 ;
        RECT 69.225 118.345 69.395 118.515 ;
        RECT 69.685 118.345 69.855 118.515 ;
        RECT 70.145 118.345 70.315 118.515 ;
        RECT 70.605 118.345 70.775 118.515 ;
        RECT 71.065 118.345 71.235 118.515 ;
        RECT 71.525 118.345 71.695 118.515 ;
        RECT 71.985 118.345 72.155 118.515 ;
        RECT 72.445 118.345 72.615 118.515 ;
        RECT 72.905 118.345 73.075 118.515 ;
        RECT 73.365 118.345 73.535 118.515 ;
        RECT 73.825 118.345 73.995 118.515 ;
        RECT 74.285 118.345 74.455 118.515 ;
        RECT 74.745 118.345 74.915 118.515 ;
        RECT 75.205 118.345 75.375 118.515 ;
        RECT 75.665 118.345 75.835 118.515 ;
        RECT 76.125 118.345 76.295 118.515 ;
        RECT 76.585 118.345 76.755 118.515 ;
        RECT 77.045 118.345 77.215 118.515 ;
        RECT 77.505 118.345 77.675 118.515 ;
        RECT 77.965 118.345 78.135 118.515 ;
        RECT 78.425 118.345 78.595 118.515 ;
        RECT 78.885 118.345 79.055 118.515 ;
        RECT 79.345 118.345 79.515 118.515 ;
        RECT 79.805 118.345 79.975 118.515 ;
        RECT 80.265 118.345 80.435 118.515 ;
        RECT 80.725 118.345 80.895 118.515 ;
        RECT 81.185 118.345 81.355 118.515 ;
        RECT 81.645 118.345 81.815 118.515 ;
        RECT 82.105 118.345 82.275 118.515 ;
        RECT 82.565 118.345 82.735 118.515 ;
        RECT 83.025 118.345 83.195 118.515 ;
        RECT 83.485 118.345 83.655 118.515 ;
        RECT 83.945 118.345 84.115 118.515 ;
        RECT 84.405 118.345 84.575 118.515 ;
        RECT 84.865 118.345 85.035 118.515 ;
        RECT 85.325 118.345 85.495 118.515 ;
        RECT 85.785 118.345 85.955 118.515 ;
        RECT 86.245 118.345 86.415 118.515 ;
        RECT 86.705 118.345 86.875 118.515 ;
        RECT 87.165 118.345 87.335 118.515 ;
        RECT 87.625 118.345 87.795 118.515 ;
        RECT 88.085 118.345 88.255 118.515 ;
        RECT 88.545 118.345 88.715 118.515 ;
        RECT 89.005 118.345 89.175 118.515 ;
        RECT 89.465 118.345 89.635 118.515 ;
        RECT 89.925 118.345 90.095 118.515 ;
        RECT 90.385 118.345 90.555 118.515 ;
        RECT 90.845 118.345 91.015 118.515 ;
        RECT 91.305 118.345 91.475 118.515 ;
        RECT 91.765 118.345 91.935 118.515 ;
        RECT 92.225 118.345 92.395 118.515 ;
        RECT 92.685 118.345 92.855 118.515 ;
        RECT 93.145 118.345 93.315 118.515 ;
        RECT 93.605 118.345 93.775 118.515 ;
        RECT 94.065 118.345 94.235 118.515 ;
        RECT 94.525 118.345 94.695 118.515 ;
        RECT 94.985 118.345 95.155 118.515 ;
        RECT 95.445 118.345 95.615 118.515 ;
        RECT 95.905 118.345 96.075 118.515 ;
        RECT 96.365 118.345 96.535 118.515 ;
        RECT 96.825 118.345 96.995 118.515 ;
        RECT 97.285 118.345 97.455 118.515 ;
        RECT 97.745 118.345 97.915 118.515 ;
        RECT 98.205 118.345 98.375 118.515 ;
        RECT 98.665 118.345 98.835 118.515 ;
        RECT 99.125 118.345 99.295 118.515 ;
        RECT 99.585 118.345 99.755 118.515 ;
        RECT 100.045 118.345 100.215 118.515 ;
        RECT 100.505 118.345 100.675 118.515 ;
        RECT 100.965 118.345 101.135 118.515 ;
        RECT 101.425 118.345 101.595 118.515 ;
        RECT 101.885 118.345 102.055 118.515 ;
        RECT 102.345 118.345 102.515 118.515 ;
        RECT 102.805 118.345 102.975 118.515 ;
        RECT 103.265 118.345 103.435 118.515 ;
        RECT 103.725 118.345 103.895 118.515 ;
        RECT 104.185 118.345 104.355 118.515 ;
        RECT 104.645 118.345 104.815 118.515 ;
        RECT 105.105 118.345 105.275 118.515 ;
        RECT 105.565 118.345 105.735 118.515 ;
        RECT 106.025 118.345 106.195 118.515 ;
        RECT 106.485 118.345 106.655 118.515 ;
        RECT 106.945 118.345 107.115 118.515 ;
        RECT 107.405 118.345 107.575 118.515 ;
        RECT 107.865 118.345 108.035 118.515 ;
        RECT 108.325 118.345 108.495 118.515 ;
        RECT 108.785 118.345 108.955 118.515 ;
        RECT 109.245 118.345 109.415 118.515 ;
        RECT 109.705 118.345 109.875 118.515 ;
        RECT 110.165 118.345 110.335 118.515 ;
        RECT 110.625 118.345 110.795 118.515 ;
        RECT 111.085 118.345 111.255 118.515 ;
        RECT 111.545 118.345 111.715 118.515 ;
        RECT 112.005 118.345 112.175 118.515 ;
        RECT 112.465 118.345 112.635 118.515 ;
        RECT 112.925 118.345 113.095 118.515 ;
        RECT 113.385 118.345 113.555 118.515 ;
        RECT 113.845 118.345 114.015 118.515 ;
        RECT 114.305 118.345 114.475 118.515 ;
        RECT 114.765 118.345 114.935 118.515 ;
        RECT 115.225 118.345 115.395 118.515 ;
        RECT 115.685 118.345 115.855 118.515 ;
        RECT 116.145 118.345 116.315 118.515 ;
        RECT 116.605 118.345 116.775 118.515 ;
        RECT 117.065 118.345 117.235 118.515 ;
        RECT 117.525 118.345 117.695 118.515 ;
        RECT 117.985 118.345 118.155 118.515 ;
        RECT 118.445 118.345 118.615 118.515 ;
        RECT 118.905 118.345 119.075 118.515 ;
        RECT 119.365 118.345 119.535 118.515 ;
        RECT 119.825 118.345 119.995 118.515 ;
        RECT 120.285 118.345 120.455 118.515 ;
        RECT 120.745 118.345 120.915 118.515 ;
        RECT 121.205 118.345 121.375 118.515 ;
        RECT 121.665 118.345 121.835 118.515 ;
        RECT 122.125 118.345 122.295 118.515 ;
        RECT 122.585 118.345 122.755 118.515 ;
        RECT 123.045 118.345 123.215 118.515 ;
        RECT 123.505 118.345 123.675 118.515 ;
        RECT 123.965 118.345 124.135 118.515 ;
        RECT 124.425 118.345 124.595 118.515 ;
        RECT 124.885 118.345 125.055 118.515 ;
        RECT 125.345 118.345 125.515 118.515 ;
        RECT 125.805 118.345 125.975 118.515 ;
        RECT 126.265 118.345 126.435 118.515 ;
        RECT 126.725 118.345 126.895 118.515 ;
        RECT 127.185 118.345 127.355 118.515 ;
        RECT 127.645 118.345 127.815 118.515 ;
        RECT 128.105 118.345 128.275 118.515 ;
        RECT 128.565 118.345 128.735 118.515 ;
        RECT 129.025 118.345 129.195 118.515 ;
        RECT 129.485 118.345 129.655 118.515 ;
        RECT 129.945 118.345 130.115 118.515 ;
        RECT 130.405 118.345 130.575 118.515 ;
        RECT 130.865 118.345 131.035 118.515 ;
        RECT 131.325 118.345 131.495 118.515 ;
        RECT 131.785 118.345 131.955 118.515 ;
        RECT 132.245 118.345 132.415 118.515 ;
        RECT 132.705 118.345 132.875 118.515 ;
        RECT 133.165 118.345 133.335 118.515 ;
        RECT 133.625 118.345 133.795 118.515 ;
        RECT 134.085 118.345 134.255 118.515 ;
        RECT 134.545 118.345 134.715 118.515 ;
        RECT 135.005 118.345 135.175 118.515 ;
        RECT 135.465 118.345 135.635 118.515 ;
        RECT 135.925 118.345 136.095 118.515 ;
        RECT 136.385 118.345 136.555 118.515 ;
        RECT 136.845 118.345 137.015 118.515 ;
        RECT 137.305 118.345 137.475 118.515 ;
        RECT 137.765 118.345 137.935 118.515 ;
        RECT 138.225 118.345 138.395 118.515 ;
        RECT 138.685 118.345 138.855 118.515 ;
        RECT 139.145 118.345 139.315 118.515 ;
        RECT 139.605 118.345 139.775 118.515 ;
        RECT 140.065 118.345 140.235 118.515 ;
        RECT 140.525 118.345 140.695 118.515 ;
        RECT 140.985 118.345 141.155 118.515 ;
        RECT 141.445 118.345 141.615 118.515 ;
        RECT 141.905 118.345 142.075 118.515 ;
        RECT 142.365 118.345 142.535 118.515 ;
        RECT 142.825 118.345 142.995 118.515 ;
        RECT 143.285 118.345 143.455 118.515 ;
        RECT 143.745 118.345 143.915 118.515 ;
        RECT 144.205 118.345 144.375 118.515 ;
        RECT 144.665 118.345 144.835 118.515 ;
        RECT 145.125 118.345 145.295 118.515 ;
        RECT 145.585 118.345 145.755 118.515 ;
        RECT 146.045 118.345 146.215 118.515 ;
        RECT 146.505 118.345 146.675 118.515 ;
        RECT 146.965 118.345 147.135 118.515 ;
        RECT 147.425 118.345 147.595 118.515 ;
        RECT 147.885 118.345 148.055 118.515 ;
        RECT 148.345 118.345 148.515 118.515 ;
        RECT 148.805 118.345 148.975 118.515 ;
        RECT 149.265 118.345 149.435 118.515 ;
        RECT 149.725 118.345 149.895 118.515 ;
        RECT 150.185 118.345 150.355 118.515 ;
        RECT 11.265 115.625 11.435 115.795 ;
        RECT 11.725 115.625 11.895 115.795 ;
        RECT 12.185 115.625 12.355 115.795 ;
        RECT 12.645 115.625 12.815 115.795 ;
        RECT 13.105 115.625 13.275 115.795 ;
        RECT 13.565 115.625 13.735 115.795 ;
        RECT 14.025 115.625 14.195 115.795 ;
        RECT 14.485 115.625 14.655 115.795 ;
        RECT 14.945 115.625 15.115 115.795 ;
        RECT 15.405 115.625 15.575 115.795 ;
        RECT 15.865 115.625 16.035 115.795 ;
        RECT 16.325 115.625 16.495 115.795 ;
        RECT 16.785 115.625 16.955 115.795 ;
        RECT 17.245 115.625 17.415 115.795 ;
        RECT 17.705 115.625 17.875 115.795 ;
        RECT 18.165 115.625 18.335 115.795 ;
        RECT 18.625 115.625 18.795 115.795 ;
        RECT 19.085 115.625 19.255 115.795 ;
        RECT 19.545 115.625 19.715 115.795 ;
        RECT 20.005 115.625 20.175 115.795 ;
        RECT 20.465 115.625 20.635 115.795 ;
        RECT 20.925 115.625 21.095 115.795 ;
        RECT 21.385 115.625 21.555 115.795 ;
        RECT 21.845 115.625 22.015 115.795 ;
        RECT 22.305 115.625 22.475 115.795 ;
        RECT 22.765 115.625 22.935 115.795 ;
        RECT 23.225 115.625 23.395 115.795 ;
        RECT 23.685 115.625 23.855 115.795 ;
        RECT 24.145 115.625 24.315 115.795 ;
        RECT 24.605 115.625 24.775 115.795 ;
        RECT 25.065 115.625 25.235 115.795 ;
        RECT 25.525 115.625 25.695 115.795 ;
        RECT 25.985 115.625 26.155 115.795 ;
        RECT 26.445 115.625 26.615 115.795 ;
        RECT 26.905 115.625 27.075 115.795 ;
        RECT 27.365 115.625 27.535 115.795 ;
        RECT 27.825 115.625 27.995 115.795 ;
        RECT 28.285 115.625 28.455 115.795 ;
        RECT 28.745 115.625 28.915 115.795 ;
        RECT 29.205 115.625 29.375 115.795 ;
        RECT 29.665 115.625 29.835 115.795 ;
        RECT 30.125 115.625 30.295 115.795 ;
        RECT 30.585 115.625 30.755 115.795 ;
        RECT 31.045 115.625 31.215 115.795 ;
        RECT 31.505 115.625 31.675 115.795 ;
        RECT 31.965 115.625 32.135 115.795 ;
        RECT 32.425 115.625 32.595 115.795 ;
        RECT 32.885 115.625 33.055 115.795 ;
        RECT 33.345 115.625 33.515 115.795 ;
        RECT 33.805 115.625 33.975 115.795 ;
        RECT 34.265 115.625 34.435 115.795 ;
        RECT 34.725 115.625 34.895 115.795 ;
        RECT 35.185 115.625 35.355 115.795 ;
        RECT 35.645 115.625 35.815 115.795 ;
        RECT 36.105 115.625 36.275 115.795 ;
        RECT 36.565 115.625 36.735 115.795 ;
        RECT 37.025 115.625 37.195 115.795 ;
        RECT 37.485 115.625 37.655 115.795 ;
        RECT 37.945 115.625 38.115 115.795 ;
        RECT 38.405 115.625 38.575 115.795 ;
        RECT 38.865 115.625 39.035 115.795 ;
        RECT 39.325 115.625 39.495 115.795 ;
        RECT 39.785 115.625 39.955 115.795 ;
        RECT 40.245 115.625 40.415 115.795 ;
        RECT 40.705 115.625 40.875 115.795 ;
        RECT 41.165 115.625 41.335 115.795 ;
        RECT 41.625 115.625 41.795 115.795 ;
        RECT 42.085 115.625 42.255 115.795 ;
        RECT 42.545 115.625 42.715 115.795 ;
        RECT 43.005 115.625 43.175 115.795 ;
        RECT 43.465 115.625 43.635 115.795 ;
        RECT 43.925 115.625 44.095 115.795 ;
        RECT 44.385 115.625 44.555 115.795 ;
        RECT 44.845 115.625 45.015 115.795 ;
        RECT 45.305 115.625 45.475 115.795 ;
        RECT 45.765 115.625 45.935 115.795 ;
        RECT 46.225 115.625 46.395 115.795 ;
        RECT 46.685 115.625 46.855 115.795 ;
        RECT 47.145 115.625 47.315 115.795 ;
        RECT 47.605 115.625 47.775 115.795 ;
        RECT 48.065 115.625 48.235 115.795 ;
        RECT 48.525 115.625 48.695 115.795 ;
        RECT 48.985 115.625 49.155 115.795 ;
        RECT 49.445 115.625 49.615 115.795 ;
        RECT 49.905 115.625 50.075 115.795 ;
        RECT 50.365 115.625 50.535 115.795 ;
        RECT 50.825 115.625 50.995 115.795 ;
        RECT 51.285 115.625 51.455 115.795 ;
        RECT 51.745 115.625 51.915 115.795 ;
        RECT 52.205 115.625 52.375 115.795 ;
        RECT 52.665 115.625 52.835 115.795 ;
        RECT 53.125 115.625 53.295 115.795 ;
        RECT 53.585 115.625 53.755 115.795 ;
        RECT 54.045 115.625 54.215 115.795 ;
        RECT 54.505 115.625 54.675 115.795 ;
        RECT 54.965 115.625 55.135 115.795 ;
        RECT 55.425 115.625 55.595 115.795 ;
        RECT 55.885 115.625 56.055 115.795 ;
        RECT 56.345 115.625 56.515 115.795 ;
        RECT 56.805 115.625 56.975 115.795 ;
        RECT 57.265 115.625 57.435 115.795 ;
        RECT 57.725 115.625 57.895 115.795 ;
        RECT 58.185 115.625 58.355 115.795 ;
        RECT 58.645 115.625 58.815 115.795 ;
        RECT 59.105 115.625 59.275 115.795 ;
        RECT 59.565 115.625 59.735 115.795 ;
        RECT 60.025 115.625 60.195 115.795 ;
        RECT 60.485 115.625 60.655 115.795 ;
        RECT 60.945 115.625 61.115 115.795 ;
        RECT 61.405 115.625 61.575 115.795 ;
        RECT 61.865 115.625 62.035 115.795 ;
        RECT 62.325 115.625 62.495 115.795 ;
        RECT 62.785 115.625 62.955 115.795 ;
        RECT 63.245 115.625 63.415 115.795 ;
        RECT 63.705 115.625 63.875 115.795 ;
        RECT 64.165 115.625 64.335 115.795 ;
        RECT 64.625 115.625 64.795 115.795 ;
        RECT 65.085 115.625 65.255 115.795 ;
        RECT 65.545 115.625 65.715 115.795 ;
        RECT 66.005 115.625 66.175 115.795 ;
        RECT 66.465 115.625 66.635 115.795 ;
        RECT 66.925 115.625 67.095 115.795 ;
        RECT 67.385 115.625 67.555 115.795 ;
        RECT 67.845 115.625 68.015 115.795 ;
        RECT 68.305 115.625 68.475 115.795 ;
        RECT 68.765 115.625 68.935 115.795 ;
        RECT 69.225 115.625 69.395 115.795 ;
        RECT 69.685 115.625 69.855 115.795 ;
        RECT 70.145 115.625 70.315 115.795 ;
        RECT 70.605 115.625 70.775 115.795 ;
        RECT 71.065 115.625 71.235 115.795 ;
        RECT 71.525 115.625 71.695 115.795 ;
        RECT 71.985 115.625 72.155 115.795 ;
        RECT 72.445 115.625 72.615 115.795 ;
        RECT 72.905 115.625 73.075 115.795 ;
        RECT 73.365 115.625 73.535 115.795 ;
        RECT 73.825 115.625 73.995 115.795 ;
        RECT 74.285 115.625 74.455 115.795 ;
        RECT 74.745 115.625 74.915 115.795 ;
        RECT 75.205 115.625 75.375 115.795 ;
        RECT 75.665 115.625 75.835 115.795 ;
        RECT 76.125 115.625 76.295 115.795 ;
        RECT 76.585 115.625 76.755 115.795 ;
        RECT 77.045 115.625 77.215 115.795 ;
        RECT 77.505 115.625 77.675 115.795 ;
        RECT 77.965 115.625 78.135 115.795 ;
        RECT 78.425 115.625 78.595 115.795 ;
        RECT 78.885 115.625 79.055 115.795 ;
        RECT 79.345 115.625 79.515 115.795 ;
        RECT 79.805 115.625 79.975 115.795 ;
        RECT 80.265 115.625 80.435 115.795 ;
        RECT 80.725 115.625 80.895 115.795 ;
        RECT 81.185 115.625 81.355 115.795 ;
        RECT 81.645 115.625 81.815 115.795 ;
        RECT 82.105 115.625 82.275 115.795 ;
        RECT 82.565 115.625 82.735 115.795 ;
        RECT 83.025 115.625 83.195 115.795 ;
        RECT 83.485 115.625 83.655 115.795 ;
        RECT 83.945 115.625 84.115 115.795 ;
        RECT 84.405 115.625 84.575 115.795 ;
        RECT 84.865 115.625 85.035 115.795 ;
        RECT 85.325 115.625 85.495 115.795 ;
        RECT 85.785 115.625 85.955 115.795 ;
        RECT 86.245 115.625 86.415 115.795 ;
        RECT 86.705 115.625 86.875 115.795 ;
        RECT 87.165 115.625 87.335 115.795 ;
        RECT 87.625 115.625 87.795 115.795 ;
        RECT 88.085 115.625 88.255 115.795 ;
        RECT 88.545 115.625 88.715 115.795 ;
        RECT 89.005 115.625 89.175 115.795 ;
        RECT 89.465 115.625 89.635 115.795 ;
        RECT 89.925 115.625 90.095 115.795 ;
        RECT 90.385 115.625 90.555 115.795 ;
        RECT 90.845 115.625 91.015 115.795 ;
        RECT 91.305 115.625 91.475 115.795 ;
        RECT 91.765 115.625 91.935 115.795 ;
        RECT 92.225 115.625 92.395 115.795 ;
        RECT 92.685 115.625 92.855 115.795 ;
        RECT 93.145 115.625 93.315 115.795 ;
        RECT 93.605 115.625 93.775 115.795 ;
        RECT 94.065 115.625 94.235 115.795 ;
        RECT 94.525 115.625 94.695 115.795 ;
        RECT 94.985 115.625 95.155 115.795 ;
        RECT 95.445 115.625 95.615 115.795 ;
        RECT 95.905 115.625 96.075 115.795 ;
        RECT 96.365 115.625 96.535 115.795 ;
        RECT 96.825 115.625 96.995 115.795 ;
        RECT 97.285 115.625 97.455 115.795 ;
        RECT 97.745 115.625 97.915 115.795 ;
        RECT 98.205 115.625 98.375 115.795 ;
        RECT 98.665 115.625 98.835 115.795 ;
        RECT 99.125 115.625 99.295 115.795 ;
        RECT 99.585 115.625 99.755 115.795 ;
        RECT 100.045 115.625 100.215 115.795 ;
        RECT 100.505 115.625 100.675 115.795 ;
        RECT 100.965 115.625 101.135 115.795 ;
        RECT 101.425 115.625 101.595 115.795 ;
        RECT 101.885 115.625 102.055 115.795 ;
        RECT 102.345 115.625 102.515 115.795 ;
        RECT 102.805 115.625 102.975 115.795 ;
        RECT 103.265 115.625 103.435 115.795 ;
        RECT 103.725 115.625 103.895 115.795 ;
        RECT 104.185 115.625 104.355 115.795 ;
        RECT 104.645 115.625 104.815 115.795 ;
        RECT 105.105 115.625 105.275 115.795 ;
        RECT 105.565 115.625 105.735 115.795 ;
        RECT 106.025 115.625 106.195 115.795 ;
        RECT 106.485 115.625 106.655 115.795 ;
        RECT 106.945 115.625 107.115 115.795 ;
        RECT 107.405 115.625 107.575 115.795 ;
        RECT 107.865 115.625 108.035 115.795 ;
        RECT 108.325 115.625 108.495 115.795 ;
        RECT 108.785 115.625 108.955 115.795 ;
        RECT 109.245 115.625 109.415 115.795 ;
        RECT 109.705 115.625 109.875 115.795 ;
        RECT 110.165 115.625 110.335 115.795 ;
        RECT 110.625 115.625 110.795 115.795 ;
        RECT 111.085 115.625 111.255 115.795 ;
        RECT 111.545 115.625 111.715 115.795 ;
        RECT 112.005 115.625 112.175 115.795 ;
        RECT 112.465 115.625 112.635 115.795 ;
        RECT 112.925 115.625 113.095 115.795 ;
        RECT 113.385 115.625 113.555 115.795 ;
        RECT 113.845 115.625 114.015 115.795 ;
        RECT 114.305 115.625 114.475 115.795 ;
        RECT 114.765 115.625 114.935 115.795 ;
        RECT 115.225 115.625 115.395 115.795 ;
        RECT 115.685 115.625 115.855 115.795 ;
        RECT 116.145 115.625 116.315 115.795 ;
        RECT 116.605 115.625 116.775 115.795 ;
        RECT 117.065 115.625 117.235 115.795 ;
        RECT 117.525 115.625 117.695 115.795 ;
        RECT 117.985 115.625 118.155 115.795 ;
        RECT 118.445 115.625 118.615 115.795 ;
        RECT 118.905 115.625 119.075 115.795 ;
        RECT 119.365 115.625 119.535 115.795 ;
        RECT 119.825 115.625 119.995 115.795 ;
        RECT 120.285 115.625 120.455 115.795 ;
        RECT 120.745 115.625 120.915 115.795 ;
        RECT 121.205 115.625 121.375 115.795 ;
        RECT 121.665 115.625 121.835 115.795 ;
        RECT 122.125 115.625 122.295 115.795 ;
        RECT 122.585 115.625 122.755 115.795 ;
        RECT 123.045 115.625 123.215 115.795 ;
        RECT 123.505 115.625 123.675 115.795 ;
        RECT 123.965 115.625 124.135 115.795 ;
        RECT 124.425 115.625 124.595 115.795 ;
        RECT 124.885 115.625 125.055 115.795 ;
        RECT 125.345 115.625 125.515 115.795 ;
        RECT 125.805 115.625 125.975 115.795 ;
        RECT 126.265 115.625 126.435 115.795 ;
        RECT 126.725 115.625 126.895 115.795 ;
        RECT 127.185 115.625 127.355 115.795 ;
        RECT 127.645 115.625 127.815 115.795 ;
        RECT 128.105 115.625 128.275 115.795 ;
        RECT 128.565 115.625 128.735 115.795 ;
        RECT 129.025 115.625 129.195 115.795 ;
        RECT 129.485 115.625 129.655 115.795 ;
        RECT 129.945 115.625 130.115 115.795 ;
        RECT 130.405 115.625 130.575 115.795 ;
        RECT 130.865 115.625 131.035 115.795 ;
        RECT 131.325 115.625 131.495 115.795 ;
        RECT 131.785 115.625 131.955 115.795 ;
        RECT 132.245 115.625 132.415 115.795 ;
        RECT 132.705 115.625 132.875 115.795 ;
        RECT 133.165 115.625 133.335 115.795 ;
        RECT 133.625 115.625 133.795 115.795 ;
        RECT 134.085 115.625 134.255 115.795 ;
        RECT 134.545 115.625 134.715 115.795 ;
        RECT 135.005 115.625 135.175 115.795 ;
        RECT 135.465 115.625 135.635 115.795 ;
        RECT 135.925 115.625 136.095 115.795 ;
        RECT 136.385 115.625 136.555 115.795 ;
        RECT 136.845 115.625 137.015 115.795 ;
        RECT 137.305 115.625 137.475 115.795 ;
        RECT 137.765 115.625 137.935 115.795 ;
        RECT 138.225 115.625 138.395 115.795 ;
        RECT 138.685 115.625 138.855 115.795 ;
        RECT 139.145 115.625 139.315 115.795 ;
        RECT 139.605 115.625 139.775 115.795 ;
        RECT 140.065 115.625 140.235 115.795 ;
        RECT 140.525 115.625 140.695 115.795 ;
        RECT 140.985 115.625 141.155 115.795 ;
        RECT 141.445 115.625 141.615 115.795 ;
        RECT 141.905 115.625 142.075 115.795 ;
        RECT 142.365 115.625 142.535 115.795 ;
        RECT 142.825 115.625 142.995 115.795 ;
        RECT 143.285 115.625 143.455 115.795 ;
        RECT 143.745 115.625 143.915 115.795 ;
        RECT 144.205 115.625 144.375 115.795 ;
        RECT 144.665 115.625 144.835 115.795 ;
        RECT 145.125 115.625 145.295 115.795 ;
        RECT 145.585 115.625 145.755 115.795 ;
        RECT 146.045 115.625 146.215 115.795 ;
        RECT 146.505 115.625 146.675 115.795 ;
        RECT 146.965 115.625 147.135 115.795 ;
        RECT 147.425 115.625 147.595 115.795 ;
        RECT 147.885 115.625 148.055 115.795 ;
        RECT 148.345 115.625 148.515 115.795 ;
        RECT 148.805 115.625 148.975 115.795 ;
        RECT 149.265 115.625 149.435 115.795 ;
        RECT 149.725 115.625 149.895 115.795 ;
        RECT 150.185 115.625 150.355 115.795 ;
        RECT 11.265 112.905 11.435 113.075 ;
        RECT 11.725 112.905 11.895 113.075 ;
        RECT 12.185 112.905 12.355 113.075 ;
        RECT 12.645 112.905 12.815 113.075 ;
        RECT 13.105 112.905 13.275 113.075 ;
        RECT 13.565 112.905 13.735 113.075 ;
        RECT 14.025 112.905 14.195 113.075 ;
        RECT 14.485 112.905 14.655 113.075 ;
        RECT 14.945 112.905 15.115 113.075 ;
        RECT 15.405 112.905 15.575 113.075 ;
        RECT 15.865 112.905 16.035 113.075 ;
        RECT 16.325 112.905 16.495 113.075 ;
        RECT 16.785 112.905 16.955 113.075 ;
        RECT 17.245 112.905 17.415 113.075 ;
        RECT 17.705 112.905 17.875 113.075 ;
        RECT 18.165 112.905 18.335 113.075 ;
        RECT 18.625 112.905 18.795 113.075 ;
        RECT 19.085 112.905 19.255 113.075 ;
        RECT 19.545 112.905 19.715 113.075 ;
        RECT 20.005 112.905 20.175 113.075 ;
        RECT 20.465 112.905 20.635 113.075 ;
        RECT 20.925 112.905 21.095 113.075 ;
        RECT 21.385 112.905 21.555 113.075 ;
        RECT 21.845 112.905 22.015 113.075 ;
        RECT 22.305 112.905 22.475 113.075 ;
        RECT 22.765 112.905 22.935 113.075 ;
        RECT 23.225 112.905 23.395 113.075 ;
        RECT 23.685 112.905 23.855 113.075 ;
        RECT 24.145 112.905 24.315 113.075 ;
        RECT 24.605 112.905 24.775 113.075 ;
        RECT 25.065 112.905 25.235 113.075 ;
        RECT 25.525 112.905 25.695 113.075 ;
        RECT 25.985 112.905 26.155 113.075 ;
        RECT 26.445 112.905 26.615 113.075 ;
        RECT 26.905 112.905 27.075 113.075 ;
        RECT 27.365 112.905 27.535 113.075 ;
        RECT 27.825 112.905 27.995 113.075 ;
        RECT 28.285 112.905 28.455 113.075 ;
        RECT 28.745 112.905 28.915 113.075 ;
        RECT 29.205 112.905 29.375 113.075 ;
        RECT 29.665 112.905 29.835 113.075 ;
        RECT 30.125 112.905 30.295 113.075 ;
        RECT 30.585 112.905 30.755 113.075 ;
        RECT 31.045 112.905 31.215 113.075 ;
        RECT 31.505 112.905 31.675 113.075 ;
        RECT 31.965 112.905 32.135 113.075 ;
        RECT 32.425 112.905 32.595 113.075 ;
        RECT 32.885 112.905 33.055 113.075 ;
        RECT 33.345 112.905 33.515 113.075 ;
        RECT 33.805 112.905 33.975 113.075 ;
        RECT 34.265 112.905 34.435 113.075 ;
        RECT 34.725 112.905 34.895 113.075 ;
        RECT 35.185 112.905 35.355 113.075 ;
        RECT 35.645 112.905 35.815 113.075 ;
        RECT 36.105 112.905 36.275 113.075 ;
        RECT 36.565 112.905 36.735 113.075 ;
        RECT 37.025 112.905 37.195 113.075 ;
        RECT 37.485 112.905 37.655 113.075 ;
        RECT 37.945 112.905 38.115 113.075 ;
        RECT 38.405 112.905 38.575 113.075 ;
        RECT 38.865 112.905 39.035 113.075 ;
        RECT 39.325 112.905 39.495 113.075 ;
        RECT 39.785 112.905 39.955 113.075 ;
        RECT 40.245 112.905 40.415 113.075 ;
        RECT 40.705 112.905 40.875 113.075 ;
        RECT 41.165 112.905 41.335 113.075 ;
        RECT 41.625 112.905 41.795 113.075 ;
        RECT 42.085 112.905 42.255 113.075 ;
        RECT 42.545 112.905 42.715 113.075 ;
        RECT 43.005 112.905 43.175 113.075 ;
        RECT 43.465 112.905 43.635 113.075 ;
        RECT 43.925 112.905 44.095 113.075 ;
        RECT 44.385 112.905 44.555 113.075 ;
        RECT 44.845 112.905 45.015 113.075 ;
        RECT 45.305 112.905 45.475 113.075 ;
        RECT 45.765 112.905 45.935 113.075 ;
        RECT 46.225 112.905 46.395 113.075 ;
        RECT 46.685 112.905 46.855 113.075 ;
        RECT 47.145 112.905 47.315 113.075 ;
        RECT 47.605 112.905 47.775 113.075 ;
        RECT 48.065 112.905 48.235 113.075 ;
        RECT 48.525 112.905 48.695 113.075 ;
        RECT 48.985 112.905 49.155 113.075 ;
        RECT 49.445 112.905 49.615 113.075 ;
        RECT 49.905 112.905 50.075 113.075 ;
        RECT 50.365 112.905 50.535 113.075 ;
        RECT 50.825 112.905 50.995 113.075 ;
        RECT 51.285 112.905 51.455 113.075 ;
        RECT 51.745 112.905 51.915 113.075 ;
        RECT 52.205 112.905 52.375 113.075 ;
        RECT 52.665 112.905 52.835 113.075 ;
        RECT 53.125 112.905 53.295 113.075 ;
        RECT 53.585 112.905 53.755 113.075 ;
        RECT 54.045 112.905 54.215 113.075 ;
        RECT 54.505 112.905 54.675 113.075 ;
        RECT 54.965 112.905 55.135 113.075 ;
        RECT 55.425 112.905 55.595 113.075 ;
        RECT 55.885 112.905 56.055 113.075 ;
        RECT 56.345 112.905 56.515 113.075 ;
        RECT 56.805 112.905 56.975 113.075 ;
        RECT 57.265 112.905 57.435 113.075 ;
        RECT 57.725 112.905 57.895 113.075 ;
        RECT 58.185 112.905 58.355 113.075 ;
        RECT 58.645 112.905 58.815 113.075 ;
        RECT 59.105 112.905 59.275 113.075 ;
        RECT 59.565 112.905 59.735 113.075 ;
        RECT 60.025 112.905 60.195 113.075 ;
        RECT 60.485 112.905 60.655 113.075 ;
        RECT 60.945 112.905 61.115 113.075 ;
        RECT 61.405 112.905 61.575 113.075 ;
        RECT 61.865 112.905 62.035 113.075 ;
        RECT 62.325 112.905 62.495 113.075 ;
        RECT 62.785 112.905 62.955 113.075 ;
        RECT 63.245 112.905 63.415 113.075 ;
        RECT 63.705 112.905 63.875 113.075 ;
        RECT 64.165 112.905 64.335 113.075 ;
        RECT 64.625 112.905 64.795 113.075 ;
        RECT 65.085 112.905 65.255 113.075 ;
        RECT 65.545 112.905 65.715 113.075 ;
        RECT 66.005 112.905 66.175 113.075 ;
        RECT 66.465 112.905 66.635 113.075 ;
        RECT 66.925 112.905 67.095 113.075 ;
        RECT 67.385 112.905 67.555 113.075 ;
        RECT 67.845 112.905 68.015 113.075 ;
        RECT 68.305 112.905 68.475 113.075 ;
        RECT 68.765 112.905 68.935 113.075 ;
        RECT 69.225 112.905 69.395 113.075 ;
        RECT 69.685 112.905 69.855 113.075 ;
        RECT 70.145 112.905 70.315 113.075 ;
        RECT 70.605 112.905 70.775 113.075 ;
        RECT 71.065 112.905 71.235 113.075 ;
        RECT 71.525 112.905 71.695 113.075 ;
        RECT 71.985 112.905 72.155 113.075 ;
        RECT 72.445 112.905 72.615 113.075 ;
        RECT 72.905 112.905 73.075 113.075 ;
        RECT 73.365 112.905 73.535 113.075 ;
        RECT 73.825 112.905 73.995 113.075 ;
        RECT 74.285 112.905 74.455 113.075 ;
        RECT 74.745 112.905 74.915 113.075 ;
        RECT 75.205 112.905 75.375 113.075 ;
        RECT 75.665 112.905 75.835 113.075 ;
        RECT 76.125 112.905 76.295 113.075 ;
        RECT 76.585 112.905 76.755 113.075 ;
        RECT 77.045 112.905 77.215 113.075 ;
        RECT 77.505 112.905 77.675 113.075 ;
        RECT 77.965 112.905 78.135 113.075 ;
        RECT 78.425 112.905 78.595 113.075 ;
        RECT 78.885 112.905 79.055 113.075 ;
        RECT 79.345 112.905 79.515 113.075 ;
        RECT 79.805 112.905 79.975 113.075 ;
        RECT 80.265 112.905 80.435 113.075 ;
        RECT 80.725 112.905 80.895 113.075 ;
        RECT 81.185 112.905 81.355 113.075 ;
        RECT 81.645 112.905 81.815 113.075 ;
        RECT 82.105 112.905 82.275 113.075 ;
        RECT 82.565 112.905 82.735 113.075 ;
        RECT 83.025 112.905 83.195 113.075 ;
        RECT 83.485 112.905 83.655 113.075 ;
        RECT 83.945 112.905 84.115 113.075 ;
        RECT 84.405 112.905 84.575 113.075 ;
        RECT 84.865 112.905 85.035 113.075 ;
        RECT 85.325 112.905 85.495 113.075 ;
        RECT 85.785 112.905 85.955 113.075 ;
        RECT 86.245 112.905 86.415 113.075 ;
        RECT 86.705 112.905 86.875 113.075 ;
        RECT 87.165 112.905 87.335 113.075 ;
        RECT 87.625 112.905 87.795 113.075 ;
        RECT 88.085 112.905 88.255 113.075 ;
        RECT 88.545 112.905 88.715 113.075 ;
        RECT 89.005 112.905 89.175 113.075 ;
        RECT 89.465 112.905 89.635 113.075 ;
        RECT 89.925 112.905 90.095 113.075 ;
        RECT 90.385 112.905 90.555 113.075 ;
        RECT 90.845 112.905 91.015 113.075 ;
        RECT 91.305 112.905 91.475 113.075 ;
        RECT 91.765 112.905 91.935 113.075 ;
        RECT 92.225 112.905 92.395 113.075 ;
        RECT 92.685 112.905 92.855 113.075 ;
        RECT 93.145 112.905 93.315 113.075 ;
        RECT 93.605 112.905 93.775 113.075 ;
        RECT 94.065 112.905 94.235 113.075 ;
        RECT 94.525 112.905 94.695 113.075 ;
        RECT 94.985 112.905 95.155 113.075 ;
        RECT 95.445 112.905 95.615 113.075 ;
        RECT 95.905 112.905 96.075 113.075 ;
        RECT 96.365 112.905 96.535 113.075 ;
        RECT 96.825 112.905 96.995 113.075 ;
        RECT 97.285 112.905 97.455 113.075 ;
        RECT 97.745 112.905 97.915 113.075 ;
        RECT 98.205 112.905 98.375 113.075 ;
        RECT 98.665 112.905 98.835 113.075 ;
        RECT 99.125 112.905 99.295 113.075 ;
        RECT 99.585 112.905 99.755 113.075 ;
        RECT 100.045 112.905 100.215 113.075 ;
        RECT 100.505 112.905 100.675 113.075 ;
        RECT 100.965 112.905 101.135 113.075 ;
        RECT 101.425 112.905 101.595 113.075 ;
        RECT 101.885 112.905 102.055 113.075 ;
        RECT 102.345 112.905 102.515 113.075 ;
        RECT 102.805 112.905 102.975 113.075 ;
        RECT 103.265 112.905 103.435 113.075 ;
        RECT 103.725 112.905 103.895 113.075 ;
        RECT 104.185 112.905 104.355 113.075 ;
        RECT 104.645 112.905 104.815 113.075 ;
        RECT 105.105 112.905 105.275 113.075 ;
        RECT 105.565 112.905 105.735 113.075 ;
        RECT 106.025 112.905 106.195 113.075 ;
        RECT 106.485 112.905 106.655 113.075 ;
        RECT 106.945 112.905 107.115 113.075 ;
        RECT 107.405 112.905 107.575 113.075 ;
        RECT 107.865 112.905 108.035 113.075 ;
        RECT 108.325 112.905 108.495 113.075 ;
        RECT 108.785 112.905 108.955 113.075 ;
        RECT 109.245 112.905 109.415 113.075 ;
        RECT 109.705 112.905 109.875 113.075 ;
        RECT 110.165 112.905 110.335 113.075 ;
        RECT 110.625 112.905 110.795 113.075 ;
        RECT 111.085 112.905 111.255 113.075 ;
        RECT 111.545 112.905 111.715 113.075 ;
        RECT 112.005 112.905 112.175 113.075 ;
        RECT 112.465 112.905 112.635 113.075 ;
        RECT 112.925 112.905 113.095 113.075 ;
        RECT 113.385 112.905 113.555 113.075 ;
        RECT 113.845 112.905 114.015 113.075 ;
        RECT 114.305 112.905 114.475 113.075 ;
        RECT 114.765 112.905 114.935 113.075 ;
        RECT 115.225 112.905 115.395 113.075 ;
        RECT 115.685 112.905 115.855 113.075 ;
        RECT 116.145 112.905 116.315 113.075 ;
        RECT 116.605 112.905 116.775 113.075 ;
        RECT 117.065 112.905 117.235 113.075 ;
        RECT 117.525 112.905 117.695 113.075 ;
        RECT 117.985 112.905 118.155 113.075 ;
        RECT 118.445 112.905 118.615 113.075 ;
        RECT 118.905 112.905 119.075 113.075 ;
        RECT 119.365 112.905 119.535 113.075 ;
        RECT 119.825 112.905 119.995 113.075 ;
        RECT 120.285 112.905 120.455 113.075 ;
        RECT 120.745 112.905 120.915 113.075 ;
        RECT 121.205 112.905 121.375 113.075 ;
        RECT 121.665 112.905 121.835 113.075 ;
        RECT 122.125 112.905 122.295 113.075 ;
        RECT 122.585 112.905 122.755 113.075 ;
        RECT 123.045 112.905 123.215 113.075 ;
        RECT 123.505 112.905 123.675 113.075 ;
        RECT 123.965 112.905 124.135 113.075 ;
        RECT 124.425 112.905 124.595 113.075 ;
        RECT 124.885 112.905 125.055 113.075 ;
        RECT 125.345 112.905 125.515 113.075 ;
        RECT 125.805 112.905 125.975 113.075 ;
        RECT 126.265 112.905 126.435 113.075 ;
        RECT 126.725 112.905 126.895 113.075 ;
        RECT 127.185 112.905 127.355 113.075 ;
        RECT 127.645 112.905 127.815 113.075 ;
        RECT 128.105 112.905 128.275 113.075 ;
        RECT 128.565 112.905 128.735 113.075 ;
        RECT 129.025 112.905 129.195 113.075 ;
        RECT 129.485 112.905 129.655 113.075 ;
        RECT 129.945 112.905 130.115 113.075 ;
        RECT 130.405 112.905 130.575 113.075 ;
        RECT 130.865 112.905 131.035 113.075 ;
        RECT 131.325 112.905 131.495 113.075 ;
        RECT 131.785 112.905 131.955 113.075 ;
        RECT 132.245 112.905 132.415 113.075 ;
        RECT 132.705 112.905 132.875 113.075 ;
        RECT 133.165 112.905 133.335 113.075 ;
        RECT 133.625 112.905 133.795 113.075 ;
        RECT 134.085 112.905 134.255 113.075 ;
        RECT 134.545 112.905 134.715 113.075 ;
        RECT 135.005 112.905 135.175 113.075 ;
        RECT 135.465 112.905 135.635 113.075 ;
        RECT 135.925 112.905 136.095 113.075 ;
        RECT 136.385 112.905 136.555 113.075 ;
        RECT 136.845 112.905 137.015 113.075 ;
        RECT 137.305 112.905 137.475 113.075 ;
        RECT 137.765 112.905 137.935 113.075 ;
        RECT 138.225 112.905 138.395 113.075 ;
        RECT 138.685 112.905 138.855 113.075 ;
        RECT 139.145 112.905 139.315 113.075 ;
        RECT 139.605 112.905 139.775 113.075 ;
        RECT 140.065 112.905 140.235 113.075 ;
        RECT 140.525 112.905 140.695 113.075 ;
        RECT 140.985 112.905 141.155 113.075 ;
        RECT 141.445 112.905 141.615 113.075 ;
        RECT 141.905 112.905 142.075 113.075 ;
        RECT 142.365 112.905 142.535 113.075 ;
        RECT 142.825 112.905 142.995 113.075 ;
        RECT 143.285 112.905 143.455 113.075 ;
        RECT 143.745 112.905 143.915 113.075 ;
        RECT 144.205 112.905 144.375 113.075 ;
        RECT 144.665 112.905 144.835 113.075 ;
        RECT 145.125 112.905 145.295 113.075 ;
        RECT 145.585 112.905 145.755 113.075 ;
        RECT 146.045 112.905 146.215 113.075 ;
        RECT 146.505 112.905 146.675 113.075 ;
        RECT 146.965 112.905 147.135 113.075 ;
        RECT 147.425 112.905 147.595 113.075 ;
        RECT 147.885 112.905 148.055 113.075 ;
        RECT 148.345 112.905 148.515 113.075 ;
        RECT 148.805 112.905 148.975 113.075 ;
        RECT 149.265 112.905 149.435 113.075 ;
        RECT 149.725 112.905 149.895 113.075 ;
        RECT 150.185 112.905 150.355 113.075 ;
        RECT 11.265 110.185 11.435 110.355 ;
        RECT 11.725 110.185 11.895 110.355 ;
        RECT 12.185 110.185 12.355 110.355 ;
        RECT 12.645 110.185 12.815 110.355 ;
        RECT 13.105 110.185 13.275 110.355 ;
        RECT 13.565 110.185 13.735 110.355 ;
        RECT 14.025 110.185 14.195 110.355 ;
        RECT 14.485 110.185 14.655 110.355 ;
        RECT 14.945 110.185 15.115 110.355 ;
        RECT 15.405 110.185 15.575 110.355 ;
        RECT 15.865 110.185 16.035 110.355 ;
        RECT 16.325 110.185 16.495 110.355 ;
        RECT 16.785 110.185 16.955 110.355 ;
        RECT 17.245 110.185 17.415 110.355 ;
        RECT 17.705 110.185 17.875 110.355 ;
        RECT 18.165 110.185 18.335 110.355 ;
        RECT 18.625 110.185 18.795 110.355 ;
        RECT 19.085 110.185 19.255 110.355 ;
        RECT 19.545 110.185 19.715 110.355 ;
        RECT 20.005 110.185 20.175 110.355 ;
        RECT 20.465 110.185 20.635 110.355 ;
        RECT 20.925 110.185 21.095 110.355 ;
        RECT 21.385 110.185 21.555 110.355 ;
        RECT 21.845 110.185 22.015 110.355 ;
        RECT 22.305 110.185 22.475 110.355 ;
        RECT 22.765 110.185 22.935 110.355 ;
        RECT 23.225 110.185 23.395 110.355 ;
        RECT 23.685 110.185 23.855 110.355 ;
        RECT 24.145 110.185 24.315 110.355 ;
        RECT 24.605 110.185 24.775 110.355 ;
        RECT 25.065 110.185 25.235 110.355 ;
        RECT 25.525 110.185 25.695 110.355 ;
        RECT 25.985 110.185 26.155 110.355 ;
        RECT 26.445 110.185 26.615 110.355 ;
        RECT 26.905 110.185 27.075 110.355 ;
        RECT 27.365 110.185 27.535 110.355 ;
        RECT 27.825 110.185 27.995 110.355 ;
        RECT 28.285 110.185 28.455 110.355 ;
        RECT 28.745 110.185 28.915 110.355 ;
        RECT 29.205 110.185 29.375 110.355 ;
        RECT 29.665 110.185 29.835 110.355 ;
        RECT 30.125 110.185 30.295 110.355 ;
        RECT 30.585 110.185 30.755 110.355 ;
        RECT 31.045 110.185 31.215 110.355 ;
        RECT 31.505 110.185 31.675 110.355 ;
        RECT 31.965 110.185 32.135 110.355 ;
        RECT 32.425 110.185 32.595 110.355 ;
        RECT 32.885 110.185 33.055 110.355 ;
        RECT 33.345 110.185 33.515 110.355 ;
        RECT 33.805 110.185 33.975 110.355 ;
        RECT 34.265 110.185 34.435 110.355 ;
        RECT 34.725 110.185 34.895 110.355 ;
        RECT 35.185 110.185 35.355 110.355 ;
        RECT 35.645 110.185 35.815 110.355 ;
        RECT 36.105 110.185 36.275 110.355 ;
        RECT 36.565 110.185 36.735 110.355 ;
        RECT 37.025 110.185 37.195 110.355 ;
        RECT 37.485 110.185 37.655 110.355 ;
        RECT 37.945 110.185 38.115 110.355 ;
        RECT 38.405 110.185 38.575 110.355 ;
        RECT 38.865 110.185 39.035 110.355 ;
        RECT 39.325 110.185 39.495 110.355 ;
        RECT 39.785 110.185 39.955 110.355 ;
        RECT 40.245 110.185 40.415 110.355 ;
        RECT 40.705 110.185 40.875 110.355 ;
        RECT 41.165 110.185 41.335 110.355 ;
        RECT 41.625 110.185 41.795 110.355 ;
        RECT 42.085 110.185 42.255 110.355 ;
        RECT 42.545 110.185 42.715 110.355 ;
        RECT 43.005 110.185 43.175 110.355 ;
        RECT 43.465 110.185 43.635 110.355 ;
        RECT 43.925 110.185 44.095 110.355 ;
        RECT 44.385 110.185 44.555 110.355 ;
        RECT 44.845 110.185 45.015 110.355 ;
        RECT 45.305 110.185 45.475 110.355 ;
        RECT 45.765 110.185 45.935 110.355 ;
        RECT 46.225 110.185 46.395 110.355 ;
        RECT 46.685 110.185 46.855 110.355 ;
        RECT 47.145 110.185 47.315 110.355 ;
        RECT 47.605 110.185 47.775 110.355 ;
        RECT 48.065 110.185 48.235 110.355 ;
        RECT 48.525 110.185 48.695 110.355 ;
        RECT 48.985 110.185 49.155 110.355 ;
        RECT 49.445 110.185 49.615 110.355 ;
        RECT 49.905 110.185 50.075 110.355 ;
        RECT 50.365 110.185 50.535 110.355 ;
        RECT 50.825 110.185 50.995 110.355 ;
        RECT 51.285 110.185 51.455 110.355 ;
        RECT 51.745 110.185 51.915 110.355 ;
        RECT 52.205 110.185 52.375 110.355 ;
        RECT 52.665 110.185 52.835 110.355 ;
        RECT 53.125 110.185 53.295 110.355 ;
        RECT 53.585 110.185 53.755 110.355 ;
        RECT 54.045 110.185 54.215 110.355 ;
        RECT 54.505 110.185 54.675 110.355 ;
        RECT 54.965 110.185 55.135 110.355 ;
        RECT 55.425 110.185 55.595 110.355 ;
        RECT 55.885 110.185 56.055 110.355 ;
        RECT 56.345 110.185 56.515 110.355 ;
        RECT 56.805 110.185 56.975 110.355 ;
        RECT 57.265 110.185 57.435 110.355 ;
        RECT 57.725 110.185 57.895 110.355 ;
        RECT 58.185 110.185 58.355 110.355 ;
        RECT 58.645 110.185 58.815 110.355 ;
        RECT 59.105 110.185 59.275 110.355 ;
        RECT 59.565 110.185 59.735 110.355 ;
        RECT 60.025 110.185 60.195 110.355 ;
        RECT 60.485 110.185 60.655 110.355 ;
        RECT 60.945 110.185 61.115 110.355 ;
        RECT 61.405 110.185 61.575 110.355 ;
        RECT 61.865 110.185 62.035 110.355 ;
        RECT 62.325 110.185 62.495 110.355 ;
        RECT 62.785 110.185 62.955 110.355 ;
        RECT 63.245 110.185 63.415 110.355 ;
        RECT 63.705 110.185 63.875 110.355 ;
        RECT 64.165 110.185 64.335 110.355 ;
        RECT 64.625 110.185 64.795 110.355 ;
        RECT 65.085 110.185 65.255 110.355 ;
        RECT 65.545 110.185 65.715 110.355 ;
        RECT 66.005 110.185 66.175 110.355 ;
        RECT 66.465 110.185 66.635 110.355 ;
        RECT 66.925 110.185 67.095 110.355 ;
        RECT 67.385 110.185 67.555 110.355 ;
        RECT 67.845 110.185 68.015 110.355 ;
        RECT 68.305 110.185 68.475 110.355 ;
        RECT 68.765 110.185 68.935 110.355 ;
        RECT 69.225 110.185 69.395 110.355 ;
        RECT 69.685 110.185 69.855 110.355 ;
        RECT 70.145 110.185 70.315 110.355 ;
        RECT 70.605 110.185 70.775 110.355 ;
        RECT 71.065 110.185 71.235 110.355 ;
        RECT 71.525 110.185 71.695 110.355 ;
        RECT 71.985 110.185 72.155 110.355 ;
        RECT 72.445 110.185 72.615 110.355 ;
        RECT 72.905 110.185 73.075 110.355 ;
        RECT 73.365 110.185 73.535 110.355 ;
        RECT 73.825 110.185 73.995 110.355 ;
        RECT 74.285 110.185 74.455 110.355 ;
        RECT 74.745 110.185 74.915 110.355 ;
        RECT 75.205 110.185 75.375 110.355 ;
        RECT 75.665 110.185 75.835 110.355 ;
        RECT 76.125 110.185 76.295 110.355 ;
        RECT 76.585 110.185 76.755 110.355 ;
        RECT 77.045 110.185 77.215 110.355 ;
        RECT 77.505 110.185 77.675 110.355 ;
        RECT 77.965 110.185 78.135 110.355 ;
        RECT 78.425 110.185 78.595 110.355 ;
        RECT 78.885 110.185 79.055 110.355 ;
        RECT 79.345 110.185 79.515 110.355 ;
        RECT 79.805 110.185 79.975 110.355 ;
        RECT 80.265 110.185 80.435 110.355 ;
        RECT 80.725 110.185 80.895 110.355 ;
        RECT 81.185 110.185 81.355 110.355 ;
        RECT 81.645 110.185 81.815 110.355 ;
        RECT 82.105 110.185 82.275 110.355 ;
        RECT 82.565 110.185 82.735 110.355 ;
        RECT 83.025 110.185 83.195 110.355 ;
        RECT 83.485 110.185 83.655 110.355 ;
        RECT 83.945 110.185 84.115 110.355 ;
        RECT 84.405 110.185 84.575 110.355 ;
        RECT 84.865 110.185 85.035 110.355 ;
        RECT 85.325 110.185 85.495 110.355 ;
        RECT 85.785 110.185 85.955 110.355 ;
        RECT 86.245 110.185 86.415 110.355 ;
        RECT 86.705 110.185 86.875 110.355 ;
        RECT 87.165 110.185 87.335 110.355 ;
        RECT 87.625 110.185 87.795 110.355 ;
        RECT 88.085 110.185 88.255 110.355 ;
        RECT 88.545 110.185 88.715 110.355 ;
        RECT 89.005 110.185 89.175 110.355 ;
        RECT 89.465 110.185 89.635 110.355 ;
        RECT 89.925 110.185 90.095 110.355 ;
        RECT 90.385 110.185 90.555 110.355 ;
        RECT 90.845 110.185 91.015 110.355 ;
        RECT 91.305 110.185 91.475 110.355 ;
        RECT 91.765 110.185 91.935 110.355 ;
        RECT 92.225 110.185 92.395 110.355 ;
        RECT 92.685 110.185 92.855 110.355 ;
        RECT 93.145 110.185 93.315 110.355 ;
        RECT 93.605 110.185 93.775 110.355 ;
        RECT 94.065 110.185 94.235 110.355 ;
        RECT 94.525 110.185 94.695 110.355 ;
        RECT 94.985 110.185 95.155 110.355 ;
        RECT 95.445 110.185 95.615 110.355 ;
        RECT 95.905 110.185 96.075 110.355 ;
        RECT 96.365 110.185 96.535 110.355 ;
        RECT 96.825 110.185 96.995 110.355 ;
        RECT 97.285 110.185 97.455 110.355 ;
        RECT 97.745 110.185 97.915 110.355 ;
        RECT 98.205 110.185 98.375 110.355 ;
        RECT 98.665 110.185 98.835 110.355 ;
        RECT 99.125 110.185 99.295 110.355 ;
        RECT 99.585 110.185 99.755 110.355 ;
        RECT 100.045 110.185 100.215 110.355 ;
        RECT 100.505 110.185 100.675 110.355 ;
        RECT 100.965 110.185 101.135 110.355 ;
        RECT 101.425 110.185 101.595 110.355 ;
        RECT 101.885 110.185 102.055 110.355 ;
        RECT 102.345 110.185 102.515 110.355 ;
        RECT 102.805 110.185 102.975 110.355 ;
        RECT 103.265 110.185 103.435 110.355 ;
        RECT 103.725 110.185 103.895 110.355 ;
        RECT 104.185 110.185 104.355 110.355 ;
        RECT 104.645 110.185 104.815 110.355 ;
        RECT 105.105 110.185 105.275 110.355 ;
        RECT 105.565 110.185 105.735 110.355 ;
        RECT 106.025 110.185 106.195 110.355 ;
        RECT 106.485 110.185 106.655 110.355 ;
        RECT 106.945 110.185 107.115 110.355 ;
        RECT 107.405 110.185 107.575 110.355 ;
        RECT 107.865 110.185 108.035 110.355 ;
        RECT 108.325 110.185 108.495 110.355 ;
        RECT 108.785 110.185 108.955 110.355 ;
        RECT 109.245 110.185 109.415 110.355 ;
        RECT 109.705 110.185 109.875 110.355 ;
        RECT 110.165 110.185 110.335 110.355 ;
        RECT 110.625 110.185 110.795 110.355 ;
        RECT 111.085 110.185 111.255 110.355 ;
        RECT 111.545 110.185 111.715 110.355 ;
        RECT 112.005 110.185 112.175 110.355 ;
        RECT 112.465 110.185 112.635 110.355 ;
        RECT 112.925 110.185 113.095 110.355 ;
        RECT 113.385 110.185 113.555 110.355 ;
        RECT 113.845 110.185 114.015 110.355 ;
        RECT 114.305 110.185 114.475 110.355 ;
        RECT 114.765 110.185 114.935 110.355 ;
        RECT 115.225 110.185 115.395 110.355 ;
        RECT 115.685 110.185 115.855 110.355 ;
        RECT 116.145 110.185 116.315 110.355 ;
        RECT 116.605 110.185 116.775 110.355 ;
        RECT 117.065 110.185 117.235 110.355 ;
        RECT 117.525 110.185 117.695 110.355 ;
        RECT 117.985 110.185 118.155 110.355 ;
        RECT 118.445 110.185 118.615 110.355 ;
        RECT 118.905 110.185 119.075 110.355 ;
        RECT 119.365 110.185 119.535 110.355 ;
        RECT 119.825 110.185 119.995 110.355 ;
        RECT 120.285 110.185 120.455 110.355 ;
        RECT 120.745 110.185 120.915 110.355 ;
        RECT 121.205 110.185 121.375 110.355 ;
        RECT 121.665 110.185 121.835 110.355 ;
        RECT 122.125 110.185 122.295 110.355 ;
        RECT 122.585 110.185 122.755 110.355 ;
        RECT 123.045 110.185 123.215 110.355 ;
        RECT 123.505 110.185 123.675 110.355 ;
        RECT 123.965 110.185 124.135 110.355 ;
        RECT 124.425 110.185 124.595 110.355 ;
        RECT 124.885 110.185 125.055 110.355 ;
        RECT 125.345 110.185 125.515 110.355 ;
        RECT 125.805 110.185 125.975 110.355 ;
        RECT 126.265 110.185 126.435 110.355 ;
        RECT 126.725 110.185 126.895 110.355 ;
        RECT 127.185 110.185 127.355 110.355 ;
        RECT 127.645 110.185 127.815 110.355 ;
        RECT 128.105 110.185 128.275 110.355 ;
        RECT 128.565 110.185 128.735 110.355 ;
        RECT 129.025 110.185 129.195 110.355 ;
        RECT 129.485 110.185 129.655 110.355 ;
        RECT 129.945 110.185 130.115 110.355 ;
        RECT 130.405 110.185 130.575 110.355 ;
        RECT 130.865 110.185 131.035 110.355 ;
        RECT 131.325 110.185 131.495 110.355 ;
        RECT 131.785 110.185 131.955 110.355 ;
        RECT 132.245 110.185 132.415 110.355 ;
        RECT 132.705 110.185 132.875 110.355 ;
        RECT 133.165 110.185 133.335 110.355 ;
        RECT 133.625 110.185 133.795 110.355 ;
        RECT 134.085 110.185 134.255 110.355 ;
        RECT 134.545 110.185 134.715 110.355 ;
        RECT 135.005 110.185 135.175 110.355 ;
        RECT 135.465 110.185 135.635 110.355 ;
        RECT 135.925 110.185 136.095 110.355 ;
        RECT 136.385 110.185 136.555 110.355 ;
        RECT 136.845 110.185 137.015 110.355 ;
        RECT 137.305 110.185 137.475 110.355 ;
        RECT 137.765 110.185 137.935 110.355 ;
        RECT 138.225 110.185 138.395 110.355 ;
        RECT 138.685 110.185 138.855 110.355 ;
        RECT 139.145 110.185 139.315 110.355 ;
        RECT 139.605 110.185 139.775 110.355 ;
        RECT 140.065 110.185 140.235 110.355 ;
        RECT 140.525 110.185 140.695 110.355 ;
        RECT 140.985 110.185 141.155 110.355 ;
        RECT 141.445 110.185 141.615 110.355 ;
        RECT 141.905 110.185 142.075 110.355 ;
        RECT 142.365 110.185 142.535 110.355 ;
        RECT 142.825 110.185 142.995 110.355 ;
        RECT 143.285 110.185 143.455 110.355 ;
        RECT 143.745 110.185 143.915 110.355 ;
        RECT 144.205 110.185 144.375 110.355 ;
        RECT 144.665 110.185 144.835 110.355 ;
        RECT 145.125 110.185 145.295 110.355 ;
        RECT 145.585 110.185 145.755 110.355 ;
        RECT 146.045 110.185 146.215 110.355 ;
        RECT 146.505 110.185 146.675 110.355 ;
        RECT 146.965 110.185 147.135 110.355 ;
        RECT 147.425 110.185 147.595 110.355 ;
        RECT 147.885 110.185 148.055 110.355 ;
        RECT 148.345 110.185 148.515 110.355 ;
        RECT 148.805 110.185 148.975 110.355 ;
        RECT 149.265 110.185 149.435 110.355 ;
        RECT 149.725 110.185 149.895 110.355 ;
        RECT 150.185 110.185 150.355 110.355 ;
        RECT 11.265 107.465 11.435 107.635 ;
        RECT 11.725 107.465 11.895 107.635 ;
        RECT 12.185 107.465 12.355 107.635 ;
        RECT 12.645 107.465 12.815 107.635 ;
        RECT 13.105 107.465 13.275 107.635 ;
        RECT 13.565 107.465 13.735 107.635 ;
        RECT 14.025 107.465 14.195 107.635 ;
        RECT 14.485 107.465 14.655 107.635 ;
        RECT 14.945 107.465 15.115 107.635 ;
        RECT 15.405 107.465 15.575 107.635 ;
        RECT 15.865 107.465 16.035 107.635 ;
        RECT 16.325 107.465 16.495 107.635 ;
        RECT 16.785 107.465 16.955 107.635 ;
        RECT 17.245 107.465 17.415 107.635 ;
        RECT 17.705 107.465 17.875 107.635 ;
        RECT 18.165 107.465 18.335 107.635 ;
        RECT 18.625 107.465 18.795 107.635 ;
        RECT 19.085 107.465 19.255 107.635 ;
        RECT 19.545 107.465 19.715 107.635 ;
        RECT 20.005 107.465 20.175 107.635 ;
        RECT 20.465 107.465 20.635 107.635 ;
        RECT 20.925 107.465 21.095 107.635 ;
        RECT 21.385 107.465 21.555 107.635 ;
        RECT 21.845 107.465 22.015 107.635 ;
        RECT 22.305 107.465 22.475 107.635 ;
        RECT 22.765 107.465 22.935 107.635 ;
        RECT 23.225 107.465 23.395 107.635 ;
        RECT 23.685 107.465 23.855 107.635 ;
        RECT 24.145 107.465 24.315 107.635 ;
        RECT 24.605 107.465 24.775 107.635 ;
        RECT 25.065 107.465 25.235 107.635 ;
        RECT 25.525 107.465 25.695 107.635 ;
        RECT 25.985 107.465 26.155 107.635 ;
        RECT 26.445 107.465 26.615 107.635 ;
        RECT 26.905 107.465 27.075 107.635 ;
        RECT 27.365 107.465 27.535 107.635 ;
        RECT 27.825 107.465 27.995 107.635 ;
        RECT 28.285 107.465 28.455 107.635 ;
        RECT 28.745 107.465 28.915 107.635 ;
        RECT 29.205 107.465 29.375 107.635 ;
        RECT 29.665 107.465 29.835 107.635 ;
        RECT 30.125 107.465 30.295 107.635 ;
        RECT 30.585 107.465 30.755 107.635 ;
        RECT 31.045 107.465 31.215 107.635 ;
        RECT 31.505 107.465 31.675 107.635 ;
        RECT 31.965 107.465 32.135 107.635 ;
        RECT 32.425 107.465 32.595 107.635 ;
        RECT 32.885 107.465 33.055 107.635 ;
        RECT 33.345 107.465 33.515 107.635 ;
        RECT 33.805 107.465 33.975 107.635 ;
        RECT 34.265 107.465 34.435 107.635 ;
        RECT 34.725 107.465 34.895 107.635 ;
        RECT 35.185 107.465 35.355 107.635 ;
        RECT 35.645 107.465 35.815 107.635 ;
        RECT 36.105 107.465 36.275 107.635 ;
        RECT 36.565 107.465 36.735 107.635 ;
        RECT 37.025 107.465 37.195 107.635 ;
        RECT 37.485 107.465 37.655 107.635 ;
        RECT 37.945 107.465 38.115 107.635 ;
        RECT 38.405 107.465 38.575 107.635 ;
        RECT 38.865 107.465 39.035 107.635 ;
        RECT 39.325 107.465 39.495 107.635 ;
        RECT 39.785 107.465 39.955 107.635 ;
        RECT 40.245 107.465 40.415 107.635 ;
        RECT 40.705 107.465 40.875 107.635 ;
        RECT 41.165 107.465 41.335 107.635 ;
        RECT 41.625 107.465 41.795 107.635 ;
        RECT 42.085 107.465 42.255 107.635 ;
        RECT 42.545 107.465 42.715 107.635 ;
        RECT 43.005 107.465 43.175 107.635 ;
        RECT 43.465 107.465 43.635 107.635 ;
        RECT 43.925 107.465 44.095 107.635 ;
        RECT 44.385 107.465 44.555 107.635 ;
        RECT 44.845 107.465 45.015 107.635 ;
        RECT 45.305 107.465 45.475 107.635 ;
        RECT 45.765 107.465 45.935 107.635 ;
        RECT 46.225 107.465 46.395 107.635 ;
        RECT 46.685 107.465 46.855 107.635 ;
        RECT 47.145 107.465 47.315 107.635 ;
        RECT 47.605 107.465 47.775 107.635 ;
        RECT 48.065 107.465 48.235 107.635 ;
        RECT 48.525 107.465 48.695 107.635 ;
        RECT 48.985 107.465 49.155 107.635 ;
        RECT 49.445 107.465 49.615 107.635 ;
        RECT 49.905 107.465 50.075 107.635 ;
        RECT 50.365 107.465 50.535 107.635 ;
        RECT 50.825 107.465 50.995 107.635 ;
        RECT 51.285 107.465 51.455 107.635 ;
        RECT 51.745 107.465 51.915 107.635 ;
        RECT 52.205 107.465 52.375 107.635 ;
        RECT 52.665 107.465 52.835 107.635 ;
        RECT 53.125 107.465 53.295 107.635 ;
        RECT 53.585 107.465 53.755 107.635 ;
        RECT 54.045 107.465 54.215 107.635 ;
        RECT 54.505 107.465 54.675 107.635 ;
        RECT 54.965 107.465 55.135 107.635 ;
        RECT 55.425 107.465 55.595 107.635 ;
        RECT 55.885 107.465 56.055 107.635 ;
        RECT 56.345 107.465 56.515 107.635 ;
        RECT 56.805 107.465 56.975 107.635 ;
        RECT 57.265 107.465 57.435 107.635 ;
        RECT 57.725 107.465 57.895 107.635 ;
        RECT 58.185 107.465 58.355 107.635 ;
        RECT 58.645 107.465 58.815 107.635 ;
        RECT 59.105 107.465 59.275 107.635 ;
        RECT 59.565 107.465 59.735 107.635 ;
        RECT 60.025 107.465 60.195 107.635 ;
        RECT 60.485 107.465 60.655 107.635 ;
        RECT 60.945 107.465 61.115 107.635 ;
        RECT 61.405 107.465 61.575 107.635 ;
        RECT 61.865 107.465 62.035 107.635 ;
        RECT 62.325 107.465 62.495 107.635 ;
        RECT 62.785 107.465 62.955 107.635 ;
        RECT 63.245 107.465 63.415 107.635 ;
        RECT 63.705 107.465 63.875 107.635 ;
        RECT 64.165 107.465 64.335 107.635 ;
        RECT 64.625 107.465 64.795 107.635 ;
        RECT 65.085 107.465 65.255 107.635 ;
        RECT 65.545 107.465 65.715 107.635 ;
        RECT 66.005 107.465 66.175 107.635 ;
        RECT 66.465 107.465 66.635 107.635 ;
        RECT 66.925 107.465 67.095 107.635 ;
        RECT 67.385 107.465 67.555 107.635 ;
        RECT 67.845 107.465 68.015 107.635 ;
        RECT 68.305 107.465 68.475 107.635 ;
        RECT 68.765 107.465 68.935 107.635 ;
        RECT 69.225 107.465 69.395 107.635 ;
        RECT 69.685 107.465 69.855 107.635 ;
        RECT 70.145 107.465 70.315 107.635 ;
        RECT 70.605 107.465 70.775 107.635 ;
        RECT 71.065 107.465 71.235 107.635 ;
        RECT 71.525 107.465 71.695 107.635 ;
        RECT 71.985 107.465 72.155 107.635 ;
        RECT 72.445 107.465 72.615 107.635 ;
        RECT 72.905 107.465 73.075 107.635 ;
        RECT 73.365 107.465 73.535 107.635 ;
        RECT 73.825 107.465 73.995 107.635 ;
        RECT 74.285 107.465 74.455 107.635 ;
        RECT 74.745 107.465 74.915 107.635 ;
        RECT 75.205 107.465 75.375 107.635 ;
        RECT 75.665 107.465 75.835 107.635 ;
        RECT 76.125 107.465 76.295 107.635 ;
        RECT 76.585 107.465 76.755 107.635 ;
        RECT 77.045 107.465 77.215 107.635 ;
        RECT 77.505 107.465 77.675 107.635 ;
        RECT 77.965 107.465 78.135 107.635 ;
        RECT 78.425 107.465 78.595 107.635 ;
        RECT 78.885 107.465 79.055 107.635 ;
        RECT 79.345 107.465 79.515 107.635 ;
        RECT 79.805 107.465 79.975 107.635 ;
        RECT 80.265 107.465 80.435 107.635 ;
        RECT 80.725 107.465 80.895 107.635 ;
        RECT 81.185 107.465 81.355 107.635 ;
        RECT 81.645 107.465 81.815 107.635 ;
        RECT 82.105 107.465 82.275 107.635 ;
        RECT 82.565 107.465 82.735 107.635 ;
        RECT 83.025 107.465 83.195 107.635 ;
        RECT 83.485 107.465 83.655 107.635 ;
        RECT 83.945 107.465 84.115 107.635 ;
        RECT 84.405 107.465 84.575 107.635 ;
        RECT 84.865 107.465 85.035 107.635 ;
        RECT 85.325 107.465 85.495 107.635 ;
        RECT 85.785 107.465 85.955 107.635 ;
        RECT 86.245 107.465 86.415 107.635 ;
        RECT 86.705 107.465 86.875 107.635 ;
        RECT 87.165 107.465 87.335 107.635 ;
        RECT 87.625 107.465 87.795 107.635 ;
        RECT 88.085 107.465 88.255 107.635 ;
        RECT 88.545 107.465 88.715 107.635 ;
        RECT 89.005 107.465 89.175 107.635 ;
        RECT 89.465 107.465 89.635 107.635 ;
        RECT 89.925 107.465 90.095 107.635 ;
        RECT 90.385 107.465 90.555 107.635 ;
        RECT 90.845 107.465 91.015 107.635 ;
        RECT 91.305 107.465 91.475 107.635 ;
        RECT 91.765 107.465 91.935 107.635 ;
        RECT 92.225 107.465 92.395 107.635 ;
        RECT 92.685 107.465 92.855 107.635 ;
        RECT 93.145 107.465 93.315 107.635 ;
        RECT 93.605 107.465 93.775 107.635 ;
        RECT 94.065 107.465 94.235 107.635 ;
        RECT 94.525 107.465 94.695 107.635 ;
        RECT 94.985 107.465 95.155 107.635 ;
        RECT 95.445 107.465 95.615 107.635 ;
        RECT 95.905 107.465 96.075 107.635 ;
        RECT 96.365 107.465 96.535 107.635 ;
        RECT 96.825 107.465 96.995 107.635 ;
        RECT 97.285 107.465 97.455 107.635 ;
        RECT 97.745 107.465 97.915 107.635 ;
        RECT 98.205 107.465 98.375 107.635 ;
        RECT 98.665 107.465 98.835 107.635 ;
        RECT 99.125 107.465 99.295 107.635 ;
        RECT 99.585 107.465 99.755 107.635 ;
        RECT 100.045 107.465 100.215 107.635 ;
        RECT 100.505 107.465 100.675 107.635 ;
        RECT 100.965 107.465 101.135 107.635 ;
        RECT 101.425 107.465 101.595 107.635 ;
        RECT 101.885 107.465 102.055 107.635 ;
        RECT 102.345 107.465 102.515 107.635 ;
        RECT 102.805 107.465 102.975 107.635 ;
        RECT 103.265 107.465 103.435 107.635 ;
        RECT 103.725 107.465 103.895 107.635 ;
        RECT 104.185 107.465 104.355 107.635 ;
        RECT 104.645 107.465 104.815 107.635 ;
        RECT 105.105 107.465 105.275 107.635 ;
        RECT 105.565 107.465 105.735 107.635 ;
        RECT 106.025 107.465 106.195 107.635 ;
        RECT 106.485 107.465 106.655 107.635 ;
        RECT 106.945 107.465 107.115 107.635 ;
        RECT 107.405 107.465 107.575 107.635 ;
        RECT 107.865 107.465 108.035 107.635 ;
        RECT 108.325 107.465 108.495 107.635 ;
        RECT 108.785 107.465 108.955 107.635 ;
        RECT 109.245 107.465 109.415 107.635 ;
        RECT 109.705 107.465 109.875 107.635 ;
        RECT 110.165 107.465 110.335 107.635 ;
        RECT 110.625 107.465 110.795 107.635 ;
        RECT 111.085 107.465 111.255 107.635 ;
        RECT 111.545 107.465 111.715 107.635 ;
        RECT 112.005 107.465 112.175 107.635 ;
        RECT 112.465 107.465 112.635 107.635 ;
        RECT 112.925 107.465 113.095 107.635 ;
        RECT 113.385 107.465 113.555 107.635 ;
        RECT 113.845 107.465 114.015 107.635 ;
        RECT 114.305 107.465 114.475 107.635 ;
        RECT 114.765 107.465 114.935 107.635 ;
        RECT 115.225 107.465 115.395 107.635 ;
        RECT 115.685 107.465 115.855 107.635 ;
        RECT 116.145 107.465 116.315 107.635 ;
        RECT 116.605 107.465 116.775 107.635 ;
        RECT 117.065 107.465 117.235 107.635 ;
        RECT 117.525 107.465 117.695 107.635 ;
        RECT 117.985 107.465 118.155 107.635 ;
        RECT 118.445 107.465 118.615 107.635 ;
        RECT 118.905 107.465 119.075 107.635 ;
        RECT 119.365 107.465 119.535 107.635 ;
        RECT 119.825 107.465 119.995 107.635 ;
        RECT 120.285 107.465 120.455 107.635 ;
        RECT 120.745 107.465 120.915 107.635 ;
        RECT 121.205 107.465 121.375 107.635 ;
        RECT 121.665 107.465 121.835 107.635 ;
        RECT 122.125 107.465 122.295 107.635 ;
        RECT 122.585 107.465 122.755 107.635 ;
        RECT 123.045 107.465 123.215 107.635 ;
        RECT 123.505 107.465 123.675 107.635 ;
        RECT 123.965 107.465 124.135 107.635 ;
        RECT 124.425 107.465 124.595 107.635 ;
        RECT 124.885 107.465 125.055 107.635 ;
        RECT 125.345 107.465 125.515 107.635 ;
        RECT 125.805 107.465 125.975 107.635 ;
        RECT 126.265 107.465 126.435 107.635 ;
        RECT 126.725 107.465 126.895 107.635 ;
        RECT 127.185 107.465 127.355 107.635 ;
        RECT 127.645 107.465 127.815 107.635 ;
        RECT 128.105 107.465 128.275 107.635 ;
        RECT 128.565 107.465 128.735 107.635 ;
        RECT 129.025 107.465 129.195 107.635 ;
        RECT 129.485 107.465 129.655 107.635 ;
        RECT 129.945 107.465 130.115 107.635 ;
        RECT 130.405 107.465 130.575 107.635 ;
        RECT 130.865 107.465 131.035 107.635 ;
        RECT 131.325 107.465 131.495 107.635 ;
        RECT 131.785 107.465 131.955 107.635 ;
        RECT 132.245 107.465 132.415 107.635 ;
        RECT 132.705 107.465 132.875 107.635 ;
        RECT 133.165 107.465 133.335 107.635 ;
        RECT 133.625 107.465 133.795 107.635 ;
        RECT 134.085 107.465 134.255 107.635 ;
        RECT 134.545 107.465 134.715 107.635 ;
        RECT 135.005 107.465 135.175 107.635 ;
        RECT 135.465 107.465 135.635 107.635 ;
        RECT 135.925 107.465 136.095 107.635 ;
        RECT 136.385 107.465 136.555 107.635 ;
        RECT 136.845 107.465 137.015 107.635 ;
        RECT 137.305 107.465 137.475 107.635 ;
        RECT 137.765 107.465 137.935 107.635 ;
        RECT 138.225 107.465 138.395 107.635 ;
        RECT 138.685 107.465 138.855 107.635 ;
        RECT 139.145 107.465 139.315 107.635 ;
        RECT 139.605 107.465 139.775 107.635 ;
        RECT 140.065 107.465 140.235 107.635 ;
        RECT 140.525 107.465 140.695 107.635 ;
        RECT 140.985 107.465 141.155 107.635 ;
        RECT 141.445 107.465 141.615 107.635 ;
        RECT 141.905 107.465 142.075 107.635 ;
        RECT 142.365 107.465 142.535 107.635 ;
        RECT 142.825 107.465 142.995 107.635 ;
        RECT 143.285 107.465 143.455 107.635 ;
        RECT 143.745 107.465 143.915 107.635 ;
        RECT 144.205 107.465 144.375 107.635 ;
        RECT 144.665 107.465 144.835 107.635 ;
        RECT 145.125 107.465 145.295 107.635 ;
        RECT 145.585 107.465 145.755 107.635 ;
        RECT 146.045 107.465 146.215 107.635 ;
        RECT 146.505 107.465 146.675 107.635 ;
        RECT 146.965 107.465 147.135 107.635 ;
        RECT 147.425 107.465 147.595 107.635 ;
        RECT 147.885 107.465 148.055 107.635 ;
        RECT 148.345 107.465 148.515 107.635 ;
        RECT 148.805 107.465 148.975 107.635 ;
        RECT 149.265 107.465 149.435 107.635 ;
        RECT 149.725 107.465 149.895 107.635 ;
        RECT 150.185 107.465 150.355 107.635 ;
        RECT 11.265 104.745 11.435 104.915 ;
        RECT 11.725 104.745 11.895 104.915 ;
        RECT 12.185 104.745 12.355 104.915 ;
        RECT 12.645 104.745 12.815 104.915 ;
        RECT 13.105 104.745 13.275 104.915 ;
        RECT 13.565 104.745 13.735 104.915 ;
        RECT 14.025 104.745 14.195 104.915 ;
        RECT 14.485 104.745 14.655 104.915 ;
        RECT 14.945 104.745 15.115 104.915 ;
        RECT 15.405 104.745 15.575 104.915 ;
        RECT 15.865 104.745 16.035 104.915 ;
        RECT 16.325 104.745 16.495 104.915 ;
        RECT 16.785 104.745 16.955 104.915 ;
        RECT 17.245 104.745 17.415 104.915 ;
        RECT 17.705 104.745 17.875 104.915 ;
        RECT 18.165 104.745 18.335 104.915 ;
        RECT 18.625 104.745 18.795 104.915 ;
        RECT 19.085 104.745 19.255 104.915 ;
        RECT 19.545 104.745 19.715 104.915 ;
        RECT 20.005 104.745 20.175 104.915 ;
        RECT 20.465 104.745 20.635 104.915 ;
        RECT 20.925 104.745 21.095 104.915 ;
        RECT 21.385 104.745 21.555 104.915 ;
        RECT 21.845 104.745 22.015 104.915 ;
        RECT 22.305 104.745 22.475 104.915 ;
        RECT 22.765 104.745 22.935 104.915 ;
        RECT 23.225 104.745 23.395 104.915 ;
        RECT 23.685 104.745 23.855 104.915 ;
        RECT 24.145 104.745 24.315 104.915 ;
        RECT 24.605 104.745 24.775 104.915 ;
        RECT 25.065 104.745 25.235 104.915 ;
        RECT 25.525 104.745 25.695 104.915 ;
        RECT 25.985 104.745 26.155 104.915 ;
        RECT 26.445 104.745 26.615 104.915 ;
        RECT 26.905 104.745 27.075 104.915 ;
        RECT 27.365 104.745 27.535 104.915 ;
        RECT 27.825 104.745 27.995 104.915 ;
        RECT 28.285 104.745 28.455 104.915 ;
        RECT 28.745 104.745 28.915 104.915 ;
        RECT 29.205 104.745 29.375 104.915 ;
        RECT 29.665 104.745 29.835 104.915 ;
        RECT 30.125 104.745 30.295 104.915 ;
        RECT 30.585 104.745 30.755 104.915 ;
        RECT 31.045 104.745 31.215 104.915 ;
        RECT 31.505 104.745 31.675 104.915 ;
        RECT 31.965 104.745 32.135 104.915 ;
        RECT 32.425 104.745 32.595 104.915 ;
        RECT 32.885 104.745 33.055 104.915 ;
        RECT 33.345 104.745 33.515 104.915 ;
        RECT 33.805 104.745 33.975 104.915 ;
        RECT 34.265 104.745 34.435 104.915 ;
        RECT 34.725 104.745 34.895 104.915 ;
        RECT 35.185 104.745 35.355 104.915 ;
        RECT 35.645 104.745 35.815 104.915 ;
        RECT 36.105 104.745 36.275 104.915 ;
        RECT 36.565 104.745 36.735 104.915 ;
        RECT 37.025 104.745 37.195 104.915 ;
        RECT 37.485 104.745 37.655 104.915 ;
        RECT 37.945 104.745 38.115 104.915 ;
        RECT 38.405 104.745 38.575 104.915 ;
        RECT 38.865 104.745 39.035 104.915 ;
        RECT 39.325 104.745 39.495 104.915 ;
        RECT 39.785 104.745 39.955 104.915 ;
        RECT 40.245 104.745 40.415 104.915 ;
        RECT 40.705 104.745 40.875 104.915 ;
        RECT 41.165 104.745 41.335 104.915 ;
        RECT 41.625 104.745 41.795 104.915 ;
        RECT 42.085 104.745 42.255 104.915 ;
        RECT 42.545 104.745 42.715 104.915 ;
        RECT 43.005 104.745 43.175 104.915 ;
        RECT 43.465 104.745 43.635 104.915 ;
        RECT 43.925 104.745 44.095 104.915 ;
        RECT 44.385 104.745 44.555 104.915 ;
        RECT 44.845 104.745 45.015 104.915 ;
        RECT 45.305 104.745 45.475 104.915 ;
        RECT 45.765 104.745 45.935 104.915 ;
        RECT 46.225 104.745 46.395 104.915 ;
        RECT 46.685 104.745 46.855 104.915 ;
        RECT 47.145 104.745 47.315 104.915 ;
        RECT 47.605 104.745 47.775 104.915 ;
        RECT 48.065 104.745 48.235 104.915 ;
        RECT 48.525 104.745 48.695 104.915 ;
        RECT 48.985 104.745 49.155 104.915 ;
        RECT 49.445 104.745 49.615 104.915 ;
        RECT 49.905 104.745 50.075 104.915 ;
        RECT 50.365 104.745 50.535 104.915 ;
        RECT 50.825 104.745 50.995 104.915 ;
        RECT 51.285 104.745 51.455 104.915 ;
        RECT 51.745 104.745 51.915 104.915 ;
        RECT 52.205 104.745 52.375 104.915 ;
        RECT 52.665 104.745 52.835 104.915 ;
        RECT 53.125 104.745 53.295 104.915 ;
        RECT 53.585 104.745 53.755 104.915 ;
        RECT 54.045 104.745 54.215 104.915 ;
        RECT 54.505 104.745 54.675 104.915 ;
        RECT 54.965 104.745 55.135 104.915 ;
        RECT 55.425 104.745 55.595 104.915 ;
        RECT 55.885 104.745 56.055 104.915 ;
        RECT 56.345 104.745 56.515 104.915 ;
        RECT 56.805 104.745 56.975 104.915 ;
        RECT 57.265 104.745 57.435 104.915 ;
        RECT 57.725 104.745 57.895 104.915 ;
        RECT 58.185 104.745 58.355 104.915 ;
        RECT 58.645 104.745 58.815 104.915 ;
        RECT 59.105 104.745 59.275 104.915 ;
        RECT 59.565 104.745 59.735 104.915 ;
        RECT 60.025 104.745 60.195 104.915 ;
        RECT 60.485 104.745 60.655 104.915 ;
        RECT 60.945 104.745 61.115 104.915 ;
        RECT 61.405 104.745 61.575 104.915 ;
        RECT 61.865 104.745 62.035 104.915 ;
        RECT 62.325 104.745 62.495 104.915 ;
        RECT 62.785 104.745 62.955 104.915 ;
        RECT 63.245 104.745 63.415 104.915 ;
        RECT 63.705 104.745 63.875 104.915 ;
        RECT 64.165 104.745 64.335 104.915 ;
        RECT 64.625 104.745 64.795 104.915 ;
        RECT 65.085 104.745 65.255 104.915 ;
        RECT 65.545 104.745 65.715 104.915 ;
        RECT 66.005 104.745 66.175 104.915 ;
        RECT 66.465 104.745 66.635 104.915 ;
        RECT 66.925 104.745 67.095 104.915 ;
        RECT 67.385 104.745 67.555 104.915 ;
        RECT 67.845 104.745 68.015 104.915 ;
        RECT 68.305 104.745 68.475 104.915 ;
        RECT 68.765 104.745 68.935 104.915 ;
        RECT 69.225 104.745 69.395 104.915 ;
        RECT 69.685 104.745 69.855 104.915 ;
        RECT 70.145 104.745 70.315 104.915 ;
        RECT 70.605 104.745 70.775 104.915 ;
        RECT 71.065 104.745 71.235 104.915 ;
        RECT 71.525 104.745 71.695 104.915 ;
        RECT 71.985 104.745 72.155 104.915 ;
        RECT 72.445 104.745 72.615 104.915 ;
        RECT 72.905 104.745 73.075 104.915 ;
        RECT 73.365 104.745 73.535 104.915 ;
        RECT 73.825 104.745 73.995 104.915 ;
        RECT 74.285 104.745 74.455 104.915 ;
        RECT 74.745 104.745 74.915 104.915 ;
        RECT 75.205 104.745 75.375 104.915 ;
        RECT 75.665 104.745 75.835 104.915 ;
        RECT 76.125 104.745 76.295 104.915 ;
        RECT 76.585 104.745 76.755 104.915 ;
        RECT 77.045 104.745 77.215 104.915 ;
        RECT 77.505 104.745 77.675 104.915 ;
        RECT 77.965 104.745 78.135 104.915 ;
        RECT 78.425 104.745 78.595 104.915 ;
        RECT 78.885 104.745 79.055 104.915 ;
        RECT 79.345 104.745 79.515 104.915 ;
        RECT 79.805 104.745 79.975 104.915 ;
        RECT 80.265 104.745 80.435 104.915 ;
        RECT 80.725 104.745 80.895 104.915 ;
        RECT 81.185 104.745 81.355 104.915 ;
        RECT 81.645 104.745 81.815 104.915 ;
        RECT 82.105 104.745 82.275 104.915 ;
        RECT 82.565 104.745 82.735 104.915 ;
        RECT 83.025 104.745 83.195 104.915 ;
        RECT 83.485 104.745 83.655 104.915 ;
        RECT 83.945 104.745 84.115 104.915 ;
        RECT 84.405 104.745 84.575 104.915 ;
        RECT 84.865 104.745 85.035 104.915 ;
        RECT 85.325 104.745 85.495 104.915 ;
        RECT 85.785 104.745 85.955 104.915 ;
        RECT 86.245 104.745 86.415 104.915 ;
        RECT 86.705 104.745 86.875 104.915 ;
        RECT 87.165 104.745 87.335 104.915 ;
        RECT 87.625 104.745 87.795 104.915 ;
        RECT 88.085 104.745 88.255 104.915 ;
        RECT 88.545 104.745 88.715 104.915 ;
        RECT 89.005 104.745 89.175 104.915 ;
        RECT 89.465 104.745 89.635 104.915 ;
        RECT 89.925 104.745 90.095 104.915 ;
        RECT 90.385 104.745 90.555 104.915 ;
        RECT 90.845 104.745 91.015 104.915 ;
        RECT 91.305 104.745 91.475 104.915 ;
        RECT 91.765 104.745 91.935 104.915 ;
        RECT 92.225 104.745 92.395 104.915 ;
        RECT 92.685 104.745 92.855 104.915 ;
        RECT 93.145 104.745 93.315 104.915 ;
        RECT 93.605 104.745 93.775 104.915 ;
        RECT 94.065 104.745 94.235 104.915 ;
        RECT 94.525 104.745 94.695 104.915 ;
        RECT 94.985 104.745 95.155 104.915 ;
        RECT 95.445 104.745 95.615 104.915 ;
        RECT 95.905 104.745 96.075 104.915 ;
        RECT 96.365 104.745 96.535 104.915 ;
        RECT 96.825 104.745 96.995 104.915 ;
        RECT 97.285 104.745 97.455 104.915 ;
        RECT 97.745 104.745 97.915 104.915 ;
        RECT 98.205 104.745 98.375 104.915 ;
        RECT 98.665 104.745 98.835 104.915 ;
        RECT 99.125 104.745 99.295 104.915 ;
        RECT 99.585 104.745 99.755 104.915 ;
        RECT 100.045 104.745 100.215 104.915 ;
        RECT 100.505 104.745 100.675 104.915 ;
        RECT 100.965 104.745 101.135 104.915 ;
        RECT 101.425 104.745 101.595 104.915 ;
        RECT 101.885 104.745 102.055 104.915 ;
        RECT 102.345 104.745 102.515 104.915 ;
        RECT 102.805 104.745 102.975 104.915 ;
        RECT 103.265 104.745 103.435 104.915 ;
        RECT 103.725 104.745 103.895 104.915 ;
        RECT 104.185 104.745 104.355 104.915 ;
        RECT 104.645 104.745 104.815 104.915 ;
        RECT 105.105 104.745 105.275 104.915 ;
        RECT 105.565 104.745 105.735 104.915 ;
        RECT 106.025 104.745 106.195 104.915 ;
        RECT 106.485 104.745 106.655 104.915 ;
        RECT 106.945 104.745 107.115 104.915 ;
        RECT 107.405 104.745 107.575 104.915 ;
        RECT 107.865 104.745 108.035 104.915 ;
        RECT 108.325 104.745 108.495 104.915 ;
        RECT 108.785 104.745 108.955 104.915 ;
        RECT 109.245 104.745 109.415 104.915 ;
        RECT 109.705 104.745 109.875 104.915 ;
        RECT 110.165 104.745 110.335 104.915 ;
        RECT 110.625 104.745 110.795 104.915 ;
        RECT 111.085 104.745 111.255 104.915 ;
        RECT 111.545 104.745 111.715 104.915 ;
        RECT 112.005 104.745 112.175 104.915 ;
        RECT 112.465 104.745 112.635 104.915 ;
        RECT 112.925 104.745 113.095 104.915 ;
        RECT 113.385 104.745 113.555 104.915 ;
        RECT 113.845 104.745 114.015 104.915 ;
        RECT 114.305 104.745 114.475 104.915 ;
        RECT 114.765 104.745 114.935 104.915 ;
        RECT 115.225 104.745 115.395 104.915 ;
        RECT 115.685 104.745 115.855 104.915 ;
        RECT 116.145 104.745 116.315 104.915 ;
        RECT 116.605 104.745 116.775 104.915 ;
        RECT 117.065 104.745 117.235 104.915 ;
        RECT 117.525 104.745 117.695 104.915 ;
        RECT 117.985 104.745 118.155 104.915 ;
        RECT 118.445 104.745 118.615 104.915 ;
        RECT 118.905 104.745 119.075 104.915 ;
        RECT 119.365 104.745 119.535 104.915 ;
        RECT 119.825 104.745 119.995 104.915 ;
        RECT 120.285 104.745 120.455 104.915 ;
        RECT 120.745 104.745 120.915 104.915 ;
        RECT 121.205 104.745 121.375 104.915 ;
        RECT 121.665 104.745 121.835 104.915 ;
        RECT 122.125 104.745 122.295 104.915 ;
        RECT 122.585 104.745 122.755 104.915 ;
        RECT 123.045 104.745 123.215 104.915 ;
        RECT 123.505 104.745 123.675 104.915 ;
        RECT 123.965 104.745 124.135 104.915 ;
        RECT 124.425 104.745 124.595 104.915 ;
        RECT 124.885 104.745 125.055 104.915 ;
        RECT 125.345 104.745 125.515 104.915 ;
        RECT 125.805 104.745 125.975 104.915 ;
        RECT 126.265 104.745 126.435 104.915 ;
        RECT 126.725 104.745 126.895 104.915 ;
        RECT 127.185 104.745 127.355 104.915 ;
        RECT 127.645 104.745 127.815 104.915 ;
        RECT 128.105 104.745 128.275 104.915 ;
        RECT 128.565 104.745 128.735 104.915 ;
        RECT 129.025 104.745 129.195 104.915 ;
        RECT 129.485 104.745 129.655 104.915 ;
        RECT 129.945 104.745 130.115 104.915 ;
        RECT 130.405 104.745 130.575 104.915 ;
        RECT 130.865 104.745 131.035 104.915 ;
        RECT 131.325 104.745 131.495 104.915 ;
        RECT 131.785 104.745 131.955 104.915 ;
        RECT 132.245 104.745 132.415 104.915 ;
        RECT 132.705 104.745 132.875 104.915 ;
        RECT 133.165 104.745 133.335 104.915 ;
        RECT 133.625 104.745 133.795 104.915 ;
        RECT 134.085 104.745 134.255 104.915 ;
        RECT 134.545 104.745 134.715 104.915 ;
        RECT 135.005 104.745 135.175 104.915 ;
        RECT 135.465 104.745 135.635 104.915 ;
        RECT 135.925 104.745 136.095 104.915 ;
        RECT 136.385 104.745 136.555 104.915 ;
        RECT 136.845 104.745 137.015 104.915 ;
        RECT 137.305 104.745 137.475 104.915 ;
        RECT 137.765 104.745 137.935 104.915 ;
        RECT 138.225 104.745 138.395 104.915 ;
        RECT 138.685 104.745 138.855 104.915 ;
        RECT 139.145 104.745 139.315 104.915 ;
        RECT 139.605 104.745 139.775 104.915 ;
        RECT 140.065 104.745 140.235 104.915 ;
        RECT 140.525 104.745 140.695 104.915 ;
        RECT 140.985 104.745 141.155 104.915 ;
        RECT 141.445 104.745 141.615 104.915 ;
        RECT 141.905 104.745 142.075 104.915 ;
        RECT 142.365 104.745 142.535 104.915 ;
        RECT 142.825 104.745 142.995 104.915 ;
        RECT 143.285 104.745 143.455 104.915 ;
        RECT 143.745 104.745 143.915 104.915 ;
        RECT 144.205 104.745 144.375 104.915 ;
        RECT 144.665 104.745 144.835 104.915 ;
        RECT 145.125 104.745 145.295 104.915 ;
        RECT 145.585 104.745 145.755 104.915 ;
        RECT 146.045 104.745 146.215 104.915 ;
        RECT 146.505 104.745 146.675 104.915 ;
        RECT 146.965 104.745 147.135 104.915 ;
        RECT 147.425 104.745 147.595 104.915 ;
        RECT 147.885 104.745 148.055 104.915 ;
        RECT 148.345 104.745 148.515 104.915 ;
        RECT 148.805 104.745 148.975 104.915 ;
        RECT 149.265 104.745 149.435 104.915 ;
        RECT 149.725 104.745 149.895 104.915 ;
        RECT 150.185 104.745 150.355 104.915 ;
        RECT 11.265 102.025 11.435 102.195 ;
        RECT 11.725 102.025 11.895 102.195 ;
        RECT 12.185 102.025 12.355 102.195 ;
        RECT 12.645 102.025 12.815 102.195 ;
        RECT 13.105 102.025 13.275 102.195 ;
        RECT 13.565 102.025 13.735 102.195 ;
        RECT 14.025 102.025 14.195 102.195 ;
        RECT 14.485 102.025 14.655 102.195 ;
        RECT 14.945 102.025 15.115 102.195 ;
        RECT 15.405 102.025 15.575 102.195 ;
        RECT 15.865 102.025 16.035 102.195 ;
        RECT 16.325 102.025 16.495 102.195 ;
        RECT 16.785 102.025 16.955 102.195 ;
        RECT 17.245 102.025 17.415 102.195 ;
        RECT 17.705 102.025 17.875 102.195 ;
        RECT 18.165 102.025 18.335 102.195 ;
        RECT 18.625 102.025 18.795 102.195 ;
        RECT 19.085 102.025 19.255 102.195 ;
        RECT 19.545 102.025 19.715 102.195 ;
        RECT 20.005 102.025 20.175 102.195 ;
        RECT 20.465 102.025 20.635 102.195 ;
        RECT 20.925 102.025 21.095 102.195 ;
        RECT 21.385 102.025 21.555 102.195 ;
        RECT 21.845 102.025 22.015 102.195 ;
        RECT 22.305 102.025 22.475 102.195 ;
        RECT 22.765 102.025 22.935 102.195 ;
        RECT 23.225 102.025 23.395 102.195 ;
        RECT 23.685 102.025 23.855 102.195 ;
        RECT 24.145 102.025 24.315 102.195 ;
        RECT 24.605 102.025 24.775 102.195 ;
        RECT 25.065 102.025 25.235 102.195 ;
        RECT 25.525 102.025 25.695 102.195 ;
        RECT 25.985 102.025 26.155 102.195 ;
        RECT 26.445 102.025 26.615 102.195 ;
        RECT 26.905 102.025 27.075 102.195 ;
        RECT 27.365 102.025 27.535 102.195 ;
        RECT 27.825 102.025 27.995 102.195 ;
        RECT 28.285 102.025 28.455 102.195 ;
        RECT 28.745 102.025 28.915 102.195 ;
        RECT 29.205 102.025 29.375 102.195 ;
        RECT 29.665 102.025 29.835 102.195 ;
        RECT 30.125 102.025 30.295 102.195 ;
        RECT 30.585 102.025 30.755 102.195 ;
        RECT 31.045 102.025 31.215 102.195 ;
        RECT 31.505 102.025 31.675 102.195 ;
        RECT 31.965 102.025 32.135 102.195 ;
        RECT 32.425 102.025 32.595 102.195 ;
        RECT 32.885 102.025 33.055 102.195 ;
        RECT 33.345 102.025 33.515 102.195 ;
        RECT 33.805 102.025 33.975 102.195 ;
        RECT 34.265 102.025 34.435 102.195 ;
        RECT 34.725 102.025 34.895 102.195 ;
        RECT 35.185 102.025 35.355 102.195 ;
        RECT 35.645 102.025 35.815 102.195 ;
        RECT 36.105 102.025 36.275 102.195 ;
        RECT 36.565 102.025 36.735 102.195 ;
        RECT 37.025 102.025 37.195 102.195 ;
        RECT 37.485 102.025 37.655 102.195 ;
        RECT 37.945 102.025 38.115 102.195 ;
        RECT 38.405 102.025 38.575 102.195 ;
        RECT 38.865 102.025 39.035 102.195 ;
        RECT 39.325 102.025 39.495 102.195 ;
        RECT 39.785 102.025 39.955 102.195 ;
        RECT 40.245 102.025 40.415 102.195 ;
        RECT 40.705 102.025 40.875 102.195 ;
        RECT 41.165 102.025 41.335 102.195 ;
        RECT 41.625 102.025 41.795 102.195 ;
        RECT 42.085 102.025 42.255 102.195 ;
        RECT 42.545 102.025 42.715 102.195 ;
        RECT 43.005 102.025 43.175 102.195 ;
        RECT 43.465 102.025 43.635 102.195 ;
        RECT 43.925 102.025 44.095 102.195 ;
        RECT 44.385 102.025 44.555 102.195 ;
        RECT 44.845 102.025 45.015 102.195 ;
        RECT 45.305 102.025 45.475 102.195 ;
        RECT 45.765 102.025 45.935 102.195 ;
        RECT 46.225 102.025 46.395 102.195 ;
        RECT 46.685 102.025 46.855 102.195 ;
        RECT 47.145 102.025 47.315 102.195 ;
        RECT 47.605 102.025 47.775 102.195 ;
        RECT 48.065 102.025 48.235 102.195 ;
        RECT 48.525 102.025 48.695 102.195 ;
        RECT 48.985 102.025 49.155 102.195 ;
        RECT 49.445 102.025 49.615 102.195 ;
        RECT 49.905 102.025 50.075 102.195 ;
        RECT 50.365 102.025 50.535 102.195 ;
        RECT 50.825 102.025 50.995 102.195 ;
        RECT 51.285 102.025 51.455 102.195 ;
        RECT 51.745 102.025 51.915 102.195 ;
        RECT 52.205 102.025 52.375 102.195 ;
        RECT 52.665 102.025 52.835 102.195 ;
        RECT 53.125 102.025 53.295 102.195 ;
        RECT 53.585 102.025 53.755 102.195 ;
        RECT 54.045 102.025 54.215 102.195 ;
        RECT 54.505 102.025 54.675 102.195 ;
        RECT 54.965 102.025 55.135 102.195 ;
        RECT 55.425 102.025 55.595 102.195 ;
        RECT 55.885 102.025 56.055 102.195 ;
        RECT 56.345 102.025 56.515 102.195 ;
        RECT 56.805 102.025 56.975 102.195 ;
        RECT 57.265 102.025 57.435 102.195 ;
        RECT 57.725 102.025 57.895 102.195 ;
        RECT 58.185 102.025 58.355 102.195 ;
        RECT 58.645 102.025 58.815 102.195 ;
        RECT 59.105 102.025 59.275 102.195 ;
        RECT 59.565 102.025 59.735 102.195 ;
        RECT 60.025 102.025 60.195 102.195 ;
        RECT 60.485 102.025 60.655 102.195 ;
        RECT 60.945 102.025 61.115 102.195 ;
        RECT 61.405 102.025 61.575 102.195 ;
        RECT 61.865 102.025 62.035 102.195 ;
        RECT 62.325 102.025 62.495 102.195 ;
        RECT 62.785 102.025 62.955 102.195 ;
        RECT 63.245 102.025 63.415 102.195 ;
        RECT 63.705 102.025 63.875 102.195 ;
        RECT 64.165 102.025 64.335 102.195 ;
        RECT 64.625 102.025 64.795 102.195 ;
        RECT 65.085 102.025 65.255 102.195 ;
        RECT 65.545 102.025 65.715 102.195 ;
        RECT 66.005 102.025 66.175 102.195 ;
        RECT 66.465 102.025 66.635 102.195 ;
        RECT 66.925 102.025 67.095 102.195 ;
        RECT 67.385 102.025 67.555 102.195 ;
        RECT 67.845 102.025 68.015 102.195 ;
        RECT 68.305 102.025 68.475 102.195 ;
        RECT 68.765 102.025 68.935 102.195 ;
        RECT 69.225 102.025 69.395 102.195 ;
        RECT 69.685 102.025 69.855 102.195 ;
        RECT 70.145 102.025 70.315 102.195 ;
        RECT 70.605 102.025 70.775 102.195 ;
        RECT 71.065 102.025 71.235 102.195 ;
        RECT 71.525 102.025 71.695 102.195 ;
        RECT 71.985 102.025 72.155 102.195 ;
        RECT 72.445 102.025 72.615 102.195 ;
        RECT 72.905 102.025 73.075 102.195 ;
        RECT 73.365 102.025 73.535 102.195 ;
        RECT 73.825 102.025 73.995 102.195 ;
        RECT 74.285 102.025 74.455 102.195 ;
        RECT 74.745 102.025 74.915 102.195 ;
        RECT 75.205 102.025 75.375 102.195 ;
        RECT 75.665 102.025 75.835 102.195 ;
        RECT 76.125 102.025 76.295 102.195 ;
        RECT 76.585 102.025 76.755 102.195 ;
        RECT 77.045 102.025 77.215 102.195 ;
        RECT 77.505 102.025 77.675 102.195 ;
        RECT 77.965 102.025 78.135 102.195 ;
        RECT 78.425 102.025 78.595 102.195 ;
        RECT 78.885 102.025 79.055 102.195 ;
        RECT 79.345 102.025 79.515 102.195 ;
        RECT 79.805 102.025 79.975 102.195 ;
        RECT 80.265 102.025 80.435 102.195 ;
        RECT 80.725 102.025 80.895 102.195 ;
        RECT 81.185 102.025 81.355 102.195 ;
        RECT 81.645 102.025 81.815 102.195 ;
        RECT 82.105 102.025 82.275 102.195 ;
        RECT 82.565 102.025 82.735 102.195 ;
        RECT 83.025 102.025 83.195 102.195 ;
        RECT 83.485 102.025 83.655 102.195 ;
        RECT 83.945 102.025 84.115 102.195 ;
        RECT 84.405 102.025 84.575 102.195 ;
        RECT 84.865 102.025 85.035 102.195 ;
        RECT 85.325 102.025 85.495 102.195 ;
        RECT 85.785 102.025 85.955 102.195 ;
        RECT 86.245 102.025 86.415 102.195 ;
        RECT 86.705 102.025 86.875 102.195 ;
        RECT 87.165 102.025 87.335 102.195 ;
        RECT 87.625 102.025 87.795 102.195 ;
        RECT 88.085 102.025 88.255 102.195 ;
        RECT 88.545 102.025 88.715 102.195 ;
        RECT 89.005 102.025 89.175 102.195 ;
        RECT 89.465 102.025 89.635 102.195 ;
        RECT 89.925 102.025 90.095 102.195 ;
        RECT 90.385 102.025 90.555 102.195 ;
        RECT 90.845 102.025 91.015 102.195 ;
        RECT 91.305 102.025 91.475 102.195 ;
        RECT 91.765 102.025 91.935 102.195 ;
        RECT 92.225 102.025 92.395 102.195 ;
        RECT 92.685 102.025 92.855 102.195 ;
        RECT 93.145 102.025 93.315 102.195 ;
        RECT 93.605 102.025 93.775 102.195 ;
        RECT 94.065 102.025 94.235 102.195 ;
        RECT 94.525 102.025 94.695 102.195 ;
        RECT 94.985 102.025 95.155 102.195 ;
        RECT 95.445 102.025 95.615 102.195 ;
        RECT 95.905 102.025 96.075 102.195 ;
        RECT 96.365 102.025 96.535 102.195 ;
        RECT 96.825 102.025 96.995 102.195 ;
        RECT 97.285 102.025 97.455 102.195 ;
        RECT 97.745 102.025 97.915 102.195 ;
        RECT 98.205 102.025 98.375 102.195 ;
        RECT 98.665 102.025 98.835 102.195 ;
        RECT 99.125 102.025 99.295 102.195 ;
        RECT 99.585 102.025 99.755 102.195 ;
        RECT 100.045 102.025 100.215 102.195 ;
        RECT 100.505 102.025 100.675 102.195 ;
        RECT 100.965 102.025 101.135 102.195 ;
        RECT 101.425 102.025 101.595 102.195 ;
        RECT 101.885 102.025 102.055 102.195 ;
        RECT 102.345 102.025 102.515 102.195 ;
        RECT 102.805 102.025 102.975 102.195 ;
        RECT 103.265 102.025 103.435 102.195 ;
        RECT 103.725 102.025 103.895 102.195 ;
        RECT 104.185 102.025 104.355 102.195 ;
        RECT 104.645 102.025 104.815 102.195 ;
        RECT 105.105 102.025 105.275 102.195 ;
        RECT 105.565 102.025 105.735 102.195 ;
        RECT 106.025 102.025 106.195 102.195 ;
        RECT 106.485 102.025 106.655 102.195 ;
        RECT 106.945 102.025 107.115 102.195 ;
        RECT 107.405 102.025 107.575 102.195 ;
        RECT 107.865 102.025 108.035 102.195 ;
        RECT 108.325 102.025 108.495 102.195 ;
        RECT 108.785 102.025 108.955 102.195 ;
        RECT 109.245 102.025 109.415 102.195 ;
        RECT 109.705 102.025 109.875 102.195 ;
        RECT 110.165 102.025 110.335 102.195 ;
        RECT 110.625 102.025 110.795 102.195 ;
        RECT 111.085 102.025 111.255 102.195 ;
        RECT 111.545 102.025 111.715 102.195 ;
        RECT 112.005 102.025 112.175 102.195 ;
        RECT 112.465 102.025 112.635 102.195 ;
        RECT 112.925 102.025 113.095 102.195 ;
        RECT 113.385 102.025 113.555 102.195 ;
        RECT 113.845 102.025 114.015 102.195 ;
        RECT 114.305 102.025 114.475 102.195 ;
        RECT 114.765 102.025 114.935 102.195 ;
        RECT 115.225 102.025 115.395 102.195 ;
        RECT 115.685 102.025 115.855 102.195 ;
        RECT 116.145 102.025 116.315 102.195 ;
        RECT 116.605 102.025 116.775 102.195 ;
        RECT 117.065 102.025 117.235 102.195 ;
        RECT 117.525 102.025 117.695 102.195 ;
        RECT 117.985 102.025 118.155 102.195 ;
        RECT 118.445 102.025 118.615 102.195 ;
        RECT 118.905 102.025 119.075 102.195 ;
        RECT 119.365 102.025 119.535 102.195 ;
        RECT 119.825 102.025 119.995 102.195 ;
        RECT 120.285 102.025 120.455 102.195 ;
        RECT 120.745 102.025 120.915 102.195 ;
        RECT 121.205 102.025 121.375 102.195 ;
        RECT 121.665 102.025 121.835 102.195 ;
        RECT 122.125 102.025 122.295 102.195 ;
        RECT 122.585 102.025 122.755 102.195 ;
        RECT 123.045 102.025 123.215 102.195 ;
        RECT 123.505 102.025 123.675 102.195 ;
        RECT 123.965 102.025 124.135 102.195 ;
        RECT 124.425 102.025 124.595 102.195 ;
        RECT 124.885 102.025 125.055 102.195 ;
        RECT 125.345 102.025 125.515 102.195 ;
        RECT 125.805 102.025 125.975 102.195 ;
        RECT 126.265 102.025 126.435 102.195 ;
        RECT 126.725 102.025 126.895 102.195 ;
        RECT 127.185 102.025 127.355 102.195 ;
        RECT 127.645 102.025 127.815 102.195 ;
        RECT 128.105 102.025 128.275 102.195 ;
        RECT 128.565 102.025 128.735 102.195 ;
        RECT 129.025 102.025 129.195 102.195 ;
        RECT 129.485 102.025 129.655 102.195 ;
        RECT 129.945 102.025 130.115 102.195 ;
        RECT 130.405 102.025 130.575 102.195 ;
        RECT 130.865 102.025 131.035 102.195 ;
        RECT 131.325 102.025 131.495 102.195 ;
        RECT 131.785 102.025 131.955 102.195 ;
        RECT 132.245 102.025 132.415 102.195 ;
        RECT 132.705 102.025 132.875 102.195 ;
        RECT 133.165 102.025 133.335 102.195 ;
        RECT 133.625 102.025 133.795 102.195 ;
        RECT 134.085 102.025 134.255 102.195 ;
        RECT 134.545 102.025 134.715 102.195 ;
        RECT 135.005 102.025 135.175 102.195 ;
        RECT 135.465 102.025 135.635 102.195 ;
        RECT 135.925 102.025 136.095 102.195 ;
        RECT 136.385 102.025 136.555 102.195 ;
        RECT 136.845 102.025 137.015 102.195 ;
        RECT 137.305 102.025 137.475 102.195 ;
        RECT 137.765 102.025 137.935 102.195 ;
        RECT 138.225 102.025 138.395 102.195 ;
        RECT 138.685 102.025 138.855 102.195 ;
        RECT 139.145 102.025 139.315 102.195 ;
        RECT 139.605 102.025 139.775 102.195 ;
        RECT 140.065 102.025 140.235 102.195 ;
        RECT 140.525 102.025 140.695 102.195 ;
        RECT 140.985 102.025 141.155 102.195 ;
        RECT 141.445 102.025 141.615 102.195 ;
        RECT 141.905 102.025 142.075 102.195 ;
        RECT 142.365 102.025 142.535 102.195 ;
        RECT 142.825 102.025 142.995 102.195 ;
        RECT 143.285 102.025 143.455 102.195 ;
        RECT 143.745 102.025 143.915 102.195 ;
        RECT 144.205 102.025 144.375 102.195 ;
        RECT 144.665 102.025 144.835 102.195 ;
        RECT 145.125 102.025 145.295 102.195 ;
        RECT 145.585 102.025 145.755 102.195 ;
        RECT 146.045 102.025 146.215 102.195 ;
        RECT 146.505 102.025 146.675 102.195 ;
        RECT 146.965 102.025 147.135 102.195 ;
        RECT 147.425 102.025 147.595 102.195 ;
        RECT 147.885 102.025 148.055 102.195 ;
        RECT 148.345 102.025 148.515 102.195 ;
        RECT 148.805 102.025 148.975 102.195 ;
        RECT 149.265 102.025 149.435 102.195 ;
        RECT 149.725 102.025 149.895 102.195 ;
        RECT 150.185 102.025 150.355 102.195 ;
        RECT 11.265 99.305 11.435 99.475 ;
        RECT 11.725 99.305 11.895 99.475 ;
        RECT 12.185 99.305 12.355 99.475 ;
        RECT 12.645 99.305 12.815 99.475 ;
        RECT 13.105 99.305 13.275 99.475 ;
        RECT 13.565 99.305 13.735 99.475 ;
        RECT 14.025 99.305 14.195 99.475 ;
        RECT 14.485 99.305 14.655 99.475 ;
        RECT 14.945 99.305 15.115 99.475 ;
        RECT 15.405 99.305 15.575 99.475 ;
        RECT 15.865 99.305 16.035 99.475 ;
        RECT 16.325 99.305 16.495 99.475 ;
        RECT 16.785 99.305 16.955 99.475 ;
        RECT 17.245 99.305 17.415 99.475 ;
        RECT 17.705 99.305 17.875 99.475 ;
        RECT 18.165 99.305 18.335 99.475 ;
        RECT 18.625 99.305 18.795 99.475 ;
        RECT 19.085 99.305 19.255 99.475 ;
        RECT 19.545 99.305 19.715 99.475 ;
        RECT 20.005 99.305 20.175 99.475 ;
        RECT 20.465 99.305 20.635 99.475 ;
        RECT 20.925 99.305 21.095 99.475 ;
        RECT 21.385 99.305 21.555 99.475 ;
        RECT 21.845 99.305 22.015 99.475 ;
        RECT 22.305 99.305 22.475 99.475 ;
        RECT 22.765 99.305 22.935 99.475 ;
        RECT 23.225 99.305 23.395 99.475 ;
        RECT 23.685 99.305 23.855 99.475 ;
        RECT 24.145 99.305 24.315 99.475 ;
        RECT 24.605 99.305 24.775 99.475 ;
        RECT 25.065 99.305 25.235 99.475 ;
        RECT 25.525 99.305 25.695 99.475 ;
        RECT 25.985 99.305 26.155 99.475 ;
        RECT 26.445 99.305 26.615 99.475 ;
        RECT 26.905 99.305 27.075 99.475 ;
        RECT 27.365 99.305 27.535 99.475 ;
        RECT 27.825 99.305 27.995 99.475 ;
        RECT 28.285 99.305 28.455 99.475 ;
        RECT 28.745 99.305 28.915 99.475 ;
        RECT 29.205 99.305 29.375 99.475 ;
        RECT 29.665 99.305 29.835 99.475 ;
        RECT 30.125 99.305 30.295 99.475 ;
        RECT 30.585 99.305 30.755 99.475 ;
        RECT 31.045 99.305 31.215 99.475 ;
        RECT 31.505 99.305 31.675 99.475 ;
        RECT 31.965 99.305 32.135 99.475 ;
        RECT 32.425 99.305 32.595 99.475 ;
        RECT 32.885 99.305 33.055 99.475 ;
        RECT 33.345 99.305 33.515 99.475 ;
        RECT 33.805 99.305 33.975 99.475 ;
        RECT 34.265 99.305 34.435 99.475 ;
        RECT 34.725 99.305 34.895 99.475 ;
        RECT 35.185 99.305 35.355 99.475 ;
        RECT 35.645 99.305 35.815 99.475 ;
        RECT 36.105 99.305 36.275 99.475 ;
        RECT 36.565 99.305 36.735 99.475 ;
        RECT 37.025 99.305 37.195 99.475 ;
        RECT 37.485 99.305 37.655 99.475 ;
        RECT 37.945 99.305 38.115 99.475 ;
        RECT 38.405 99.305 38.575 99.475 ;
        RECT 38.865 99.305 39.035 99.475 ;
        RECT 39.325 99.305 39.495 99.475 ;
        RECT 39.785 99.305 39.955 99.475 ;
        RECT 40.245 99.305 40.415 99.475 ;
        RECT 40.705 99.305 40.875 99.475 ;
        RECT 41.165 99.305 41.335 99.475 ;
        RECT 41.625 99.305 41.795 99.475 ;
        RECT 42.085 99.305 42.255 99.475 ;
        RECT 42.545 99.305 42.715 99.475 ;
        RECT 43.005 99.305 43.175 99.475 ;
        RECT 43.465 99.305 43.635 99.475 ;
        RECT 43.925 99.305 44.095 99.475 ;
        RECT 44.385 99.305 44.555 99.475 ;
        RECT 44.845 99.305 45.015 99.475 ;
        RECT 45.305 99.305 45.475 99.475 ;
        RECT 45.765 99.305 45.935 99.475 ;
        RECT 46.225 99.305 46.395 99.475 ;
        RECT 46.685 99.305 46.855 99.475 ;
        RECT 47.145 99.305 47.315 99.475 ;
        RECT 47.605 99.305 47.775 99.475 ;
        RECT 48.065 99.305 48.235 99.475 ;
        RECT 48.525 99.305 48.695 99.475 ;
        RECT 48.985 99.305 49.155 99.475 ;
        RECT 49.445 99.305 49.615 99.475 ;
        RECT 49.905 99.305 50.075 99.475 ;
        RECT 50.365 99.305 50.535 99.475 ;
        RECT 50.825 99.305 50.995 99.475 ;
        RECT 51.285 99.305 51.455 99.475 ;
        RECT 51.745 99.305 51.915 99.475 ;
        RECT 52.205 99.305 52.375 99.475 ;
        RECT 52.665 99.305 52.835 99.475 ;
        RECT 53.125 99.305 53.295 99.475 ;
        RECT 53.585 99.305 53.755 99.475 ;
        RECT 54.045 99.305 54.215 99.475 ;
        RECT 54.505 99.305 54.675 99.475 ;
        RECT 54.965 99.305 55.135 99.475 ;
        RECT 55.425 99.305 55.595 99.475 ;
        RECT 55.885 99.305 56.055 99.475 ;
        RECT 56.345 99.305 56.515 99.475 ;
        RECT 56.805 99.305 56.975 99.475 ;
        RECT 57.265 99.305 57.435 99.475 ;
        RECT 57.725 99.305 57.895 99.475 ;
        RECT 58.185 99.305 58.355 99.475 ;
        RECT 58.645 99.305 58.815 99.475 ;
        RECT 59.105 99.305 59.275 99.475 ;
        RECT 59.565 99.305 59.735 99.475 ;
        RECT 60.025 99.305 60.195 99.475 ;
        RECT 60.485 99.305 60.655 99.475 ;
        RECT 60.945 99.305 61.115 99.475 ;
        RECT 61.405 99.305 61.575 99.475 ;
        RECT 61.865 99.305 62.035 99.475 ;
        RECT 62.325 99.305 62.495 99.475 ;
        RECT 62.785 99.305 62.955 99.475 ;
        RECT 63.245 99.305 63.415 99.475 ;
        RECT 63.705 99.305 63.875 99.475 ;
        RECT 64.165 99.305 64.335 99.475 ;
        RECT 64.625 99.305 64.795 99.475 ;
        RECT 65.085 99.305 65.255 99.475 ;
        RECT 65.545 99.305 65.715 99.475 ;
        RECT 66.005 99.305 66.175 99.475 ;
        RECT 66.465 99.305 66.635 99.475 ;
        RECT 66.925 99.305 67.095 99.475 ;
        RECT 67.385 99.305 67.555 99.475 ;
        RECT 67.845 99.305 68.015 99.475 ;
        RECT 68.305 99.305 68.475 99.475 ;
        RECT 68.765 99.305 68.935 99.475 ;
        RECT 69.225 99.305 69.395 99.475 ;
        RECT 69.685 99.305 69.855 99.475 ;
        RECT 70.145 99.305 70.315 99.475 ;
        RECT 70.605 99.305 70.775 99.475 ;
        RECT 71.065 99.305 71.235 99.475 ;
        RECT 71.525 99.305 71.695 99.475 ;
        RECT 71.985 99.305 72.155 99.475 ;
        RECT 72.445 99.305 72.615 99.475 ;
        RECT 72.905 99.305 73.075 99.475 ;
        RECT 73.365 99.305 73.535 99.475 ;
        RECT 73.825 99.305 73.995 99.475 ;
        RECT 74.285 99.305 74.455 99.475 ;
        RECT 74.745 99.305 74.915 99.475 ;
        RECT 75.205 99.305 75.375 99.475 ;
        RECT 75.665 99.305 75.835 99.475 ;
        RECT 76.125 99.305 76.295 99.475 ;
        RECT 76.585 99.305 76.755 99.475 ;
        RECT 77.045 99.305 77.215 99.475 ;
        RECT 77.505 99.305 77.675 99.475 ;
        RECT 77.965 99.305 78.135 99.475 ;
        RECT 78.425 99.305 78.595 99.475 ;
        RECT 78.885 99.305 79.055 99.475 ;
        RECT 79.345 99.305 79.515 99.475 ;
        RECT 79.805 99.305 79.975 99.475 ;
        RECT 80.265 99.305 80.435 99.475 ;
        RECT 80.725 99.305 80.895 99.475 ;
        RECT 81.185 99.305 81.355 99.475 ;
        RECT 81.645 99.305 81.815 99.475 ;
        RECT 82.105 99.305 82.275 99.475 ;
        RECT 82.565 99.305 82.735 99.475 ;
        RECT 83.025 99.305 83.195 99.475 ;
        RECT 83.485 99.305 83.655 99.475 ;
        RECT 83.945 99.305 84.115 99.475 ;
        RECT 84.405 99.305 84.575 99.475 ;
        RECT 84.865 99.305 85.035 99.475 ;
        RECT 85.325 99.305 85.495 99.475 ;
        RECT 85.785 99.305 85.955 99.475 ;
        RECT 86.245 99.305 86.415 99.475 ;
        RECT 86.705 99.305 86.875 99.475 ;
        RECT 87.165 99.305 87.335 99.475 ;
        RECT 87.625 99.305 87.795 99.475 ;
        RECT 88.085 99.305 88.255 99.475 ;
        RECT 88.545 99.305 88.715 99.475 ;
        RECT 89.005 99.305 89.175 99.475 ;
        RECT 89.465 99.305 89.635 99.475 ;
        RECT 89.925 99.305 90.095 99.475 ;
        RECT 90.385 99.305 90.555 99.475 ;
        RECT 90.845 99.305 91.015 99.475 ;
        RECT 91.305 99.305 91.475 99.475 ;
        RECT 91.765 99.305 91.935 99.475 ;
        RECT 92.225 99.305 92.395 99.475 ;
        RECT 92.685 99.305 92.855 99.475 ;
        RECT 93.145 99.305 93.315 99.475 ;
        RECT 93.605 99.305 93.775 99.475 ;
        RECT 94.065 99.305 94.235 99.475 ;
        RECT 94.525 99.305 94.695 99.475 ;
        RECT 94.985 99.305 95.155 99.475 ;
        RECT 95.445 99.305 95.615 99.475 ;
        RECT 95.905 99.305 96.075 99.475 ;
        RECT 96.365 99.305 96.535 99.475 ;
        RECT 96.825 99.305 96.995 99.475 ;
        RECT 97.285 99.305 97.455 99.475 ;
        RECT 97.745 99.305 97.915 99.475 ;
        RECT 98.205 99.305 98.375 99.475 ;
        RECT 98.665 99.305 98.835 99.475 ;
        RECT 99.125 99.305 99.295 99.475 ;
        RECT 99.585 99.305 99.755 99.475 ;
        RECT 100.045 99.305 100.215 99.475 ;
        RECT 100.505 99.305 100.675 99.475 ;
        RECT 100.965 99.305 101.135 99.475 ;
        RECT 101.425 99.305 101.595 99.475 ;
        RECT 101.885 99.305 102.055 99.475 ;
        RECT 102.345 99.305 102.515 99.475 ;
        RECT 102.805 99.305 102.975 99.475 ;
        RECT 103.265 99.305 103.435 99.475 ;
        RECT 103.725 99.305 103.895 99.475 ;
        RECT 104.185 99.305 104.355 99.475 ;
        RECT 104.645 99.305 104.815 99.475 ;
        RECT 105.105 99.305 105.275 99.475 ;
        RECT 105.565 99.305 105.735 99.475 ;
        RECT 106.025 99.305 106.195 99.475 ;
        RECT 106.485 99.305 106.655 99.475 ;
        RECT 106.945 99.305 107.115 99.475 ;
        RECT 107.405 99.305 107.575 99.475 ;
        RECT 107.865 99.305 108.035 99.475 ;
        RECT 108.325 99.305 108.495 99.475 ;
        RECT 108.785 99.305 108.955 99.475 ;
        RECT 109.245 99.305 109.415 99.475 ;
        RECT 109.705 99.305 109.875 99.475 ;
        RECT 110.165 99.305 110.335 99.475 ;
        RECT 110.625 99.305 110.795 99.475 ;
        RECT 111.085 99.305 111.255 99.475 ;
        RECT 111.545 99.305 111.715 99.475 ;
        RECT 112.005 99.305 112.175 99.475 ;
        RECT 112.465 99.305 112.635 99.475 ;
        RECT 112.925 99.305 113.095 99.475 ;
        RECT 113.385 99.305 113.555 99.475 ;
        RECT 113.845 99.305 114.015 99.475 ;
        RECT 114.305 99.305 114.475 99.475 ;
        RECT 114.765 99.305 114.935 99.475 ;
        RECT 115.225 99.305 115.395 99.475 ;
        RECT 115.685 99.305 115.855 99.475 ;
        RECT 116.145 99.305 116.315 99.475 ;
        RECT 116.605 99.305 116.775 99.475 ;
        RECT 117.065 99.305 117.235 99.475 ;
        RECT 117.525 99.305 117.695 99.475 ;
        RECT 117.985 99.305 118.155 99.475 ;
        RECT 118.445 99.305 118.615 99.475 ;
        RECT 118.905 99.305 119.075 99.475 ;
        RECT 119.365 99.305 119.535 99.475 ;
        RECT 119.825 99.305 119.995 99.475 ;
        RECT 120.285 99.305 120.455 99.475 ;
        RECT 120.745 99.305 120.915 99.475 ;
        RECT 121.205 99.305 121.375 99.475 ;
        RECT 121.665 99.305 121.835 99.475 ;
        RECT 122.125 99.305 122.295 99.475 ;
        RECT 122.585 99.305 122.755 99.475 ;
        RECT 123.045 99.305 123.215 99.475 ;
        RECT 123.505 99.305 123.675 99.475 ;
        RECT 123.965 99.305 124.135 99.475 ;
        RECT 124.425 99.305 124.595 99.475 ;
        RECT 124.885 99.305 125.055 99.475 ;
        RECT 125.345 99.305 125.515 99.475 ;
        RECT 125.805 99.305 125.975 99.475 ;
        RECT 126.265 99.305 126.435 99.475 ;
        RECT 126.725 99.305 126.895 99.475 ;
        RECT 127.185 99.305 127.355 99.475 ;
        RECT 127.645 99.305 127.815 99.475 ;
        RECT 128.105 99.305 128.275 99.475 ;
        RECT 128.565 99.305 128.735 99.475 ;
        RECT 129.025 99.305 129.195 99.475 ;
        RECT 129.485 99.305 129.655 99.475 ;
        RECT 129.945 99.305 130.115 99.475 ;
        RECT 130.405 99.305 130.575 99.475 ;
        RECT 130.865 99.305 131.035 99.475 ;
        RECT 131.325 99.305 131.495 99.475 ;
        RECT 131.785 99.305 131.955 99.475 ;
        RECT 132.245 99.305 132.415 99.475 ;
        RECT 132.705 99.305 132.875 99.475 ;
        RECT 133.165 99.305 133.335 99.475 ;
        RECT 133.625 99.305 133.795 99.475 ;
        RECT 134.085 99.305 134.255 99.475 ;
        RECT 134.545 99.305 134.715 99.475 ;
        RECT 135.005 99.305 135.175 99.475 ;
        RECT 135.465 99.305 135.635 99.475 ;
        RECT 135.925 99.305 136.095 99.475 ;
        RECT 136.385 99.305 136.555 99.475 ;
        RECT 136.845 99.305 137.015 99.475 ;
        RECT 137.305 99.305 137.475 99.475 ;
        RECT 137.765 99.305 137.935 99.475 ;
        RECT 138.225 99.305 138.395 99.475 ;
        RECT 138.685 99.305 138.855 99.475 ;
        RECT 139.145 99.305 139.315 99.475 ;
        RECT 139.605 99.305 139.775 99.475 ;
        RECT 140.065 99.305 140.235 99.475 ;
        RECT 140.525 99.305 140.695 99.475 ;
        RECT 140.985 99.305 141.155 99.475 ;
        RECT 141.445 99.305 141.615 99.475 ;
        RECT 141.905 99.305 142.075 99.475 ;
        RECT 142.365 99.305 142.535 99.475 ;
        RECT 142.825 99.305 142.995 99.475 ;
        RECT 143.285 99.305 143.455 99.475 ;
        RECT 143.745 99.305 143.915 99.475 ;
        RECT 144.205 99.305 144.375 99.475 ;
        RECT 144.665 99.305 144.835 99.475 ;
        RECT 145.125 99.305 145.295 99.475 ;
        RECT 145.585 99.305 145.755 99.475 ;
        RECT 146.045 99.305 146.215 99.475 ;
        RECT 146.505 99.305 146.675 99.475 ;
        RECT 146.965 99.305 147.135 99.475 ;
        RECT 147.425 99.305 147.595 99.475 ;
        RECT 147.885 99.305 148.055 99.475 ;
        RECT 148.345 99.305 148.515 99.475 ;
        RECT 148.805 99.305 148.975 99.475 ;
        RECT 149.265 99.305 149.435 99.475 ;
        RECT 149.725 99.305 149.895 99.475 ;
        RECT 150.185 99.305 150.355 99.475 ;
        RECT 11.265 96.585 11.435 96.755 ;
        RECT 11.725 96.585 11.895 96.755 ;
        RECT 12.185 96.585 12.355 96.755 ;
        RECT 12.645 96.585 12.815 96.755 ;
        RECT 13.105 96.585 13.275 96.755 ;
        RECT 13.565 96.585 13.735 96.755 ;
        RECT 14.025 96.585 14.195 96.755 ;
        RECT 14.485 96.585 14.655 96.755 ;
        RECT 14.945 96.585 15.115 96.755 ;
        RECT 15.405 96.585 15.575 96.755 ;
        RECT 15.865 96.585 16.035 96.755 ;
        RECT 16.325 96.585 16.495 96.755 ;
        RECT 16.785 96.585 16.955 96.755 ;
        RECT 17.245 96.585 17.415 96.755 ;
        RECT 17.705 96.585 17.875 96.755 ;
        RECT 18.165 96.585 18.335 96.755 ;
        RECT 18.625 96.585 18.795 96.755 ;
        RECT 19.085 96.585 19.255 96.755 ;
        RECT 19.545 96.585 19.715 96.755 ;
        RECT 20.005 96.585 20.175 96.755 ;
        RECT 20.465 96.585 20.635 96.755 ;
        RECT 20.925 96.585 21.095 96.755 ;
        RECT 21.385 96.585 21.555 96.755 ;
        RECT 21.845 96.585 22.015 96.755 ;
        RECT 22.305 96.585 22.475 96.755 ;
        RECT 22.765 96.585 22.935 96.755 ;
        RECT 23.225 96.585 23.395 96.755 ;
        RECT 23.685 96.585 23.855 96.755 ;
        RECT 24.145 96.585 24.315 96.755 ;
        RECT 24.605 96.585 24.775 96.755 ;
        RECT 25.065 96.585 25.235 96.755 ;
        RECT 25.525 96.585 25.695 96.755 ;
        RECT 25.985 96.585 26.155 96.755 ;
        RECT 26.445 96.585 26.615 96.755 ;
        RECT 26.905 96.585 27.075 96.755 ;
        RECT 27.365 96.585 27.535 96.755 ;
        RECT 27.825 96.585 27.995 96.755 ;
        RECT 28.285 96.585 28.455 96.755 ;
        RECT 28.745 96.585 28.915 96.755 ;
        RECT 29.205 96.585 29.375 96.755 ;
        RECT 29.665 96.585 29.835 96.755 ;
        RECT 30.125 96.585 30.295 96.755 ;
        RECT 30.585 96.585 30.755 96.755 ;
        RECT 31.045 96.585 31.215 96.755 ;
        RECT 31.505 96.585 31.675 96.755 ;
        RECT 31.965 96.585 32.135 96.755 ;
        RECT 32.425 96.585 32.595 96.755 ;
        RECT 32.885 96.585 33.055 96.755 ;
        RECT 33.345 96.585 33.515 96.755 ;
        RECT 33.805 96.585 33.975 96.755 ;
        RECT 34.265 96.585 34.435 96.755 ;
        RECT 34.725 96.585 34.895 96.755 ;
        RECT 35.185 96.585 35.355 96.755 ;
        RECT 35.645 96.585 35.815 96.755 ;
        RECT 36.105 96.585 36.275 96.755 ;
        RECT 36.565 96.585 36.735 96.755 ;
        RECT 37.025 96.585 37.195 96.755 ;
        RECT 37.485 96.585 37.655 96.755 ;
        RECT 37.945 96.585 38.115 96.755 ;
        RECT 38.405 96.585 38.575 96.755 ;
        RECT 38.865 96.585 39.035 96.755 ;
        RECT 39.325 96.585 39.495 96.755 ;
        RECT 39.785 96.585 39.955 96.755 ;
        RECT 40.245 96.585 40.415 96.755 ;
        RECT 40.705 96.585 40.875 96.755 ;
        RECT 41.165 96.585 41.335 96.755 ;
        RECT 41.625 96.585 41.795 96.755 ;
        RECT 42.085 96.585 42.255 96.755 ;
        RECT 42.545 96.585 42.715 96.755 ;
        RECT 43.005 96.585 43.175 96.755 ;
        RECT 43.465 96.585 43.635 96.755 ;
        RECT 43.925 96.585 44.095 96.755 ;
        RECT 44.385 96.585 44.555 96.755 ;
        RECT 44.845 96.585 45.015 96.755 ;
        RECT 45.305 96.585 45.475 96.755 ;
        RECT 45.765 96.585 45.935 96.755 ;
        RECT 46.225 96.585 46.395 96.755 ;
        RECT 46.685 96.585 46.855 96.755 ;
        RECT 47.145 96.585 47.315 96.755 ;
        RECT 47.605 96.585 47.775 96.755 ;
        RECT 48.065 96.585 48.235 96.755 ;
        RECT 48.525 96.585 48.695 96.755 ;
        RECT 48.985 96.585 49.155 96.755 ;
        RECT 49.445 96.585 49.615 96.755 ;
        RECT 49.905 96.585 50.075 96.755 ;
        RECT 50.365 96.585 50.535 96.755 ;
        RECT 50.825 96.585 50.995 96.755 ;
        RECT 51.285 96.585 51.455 96.755 ;
        RECT 51.745 96.585 51.915 96.755 ;
        RECT 52.205 96.585 52.375 96.755 ;
        RECT 52.665 96.585 52.835 96.755 ;
        RECT 53.125 96.585 53.295 96.755 ;
        RECT 53.585 96.585 53.755 96.755 ;
        RECT 54.045 96.585 54.215 96.755 ;
        RECT 54.505 96.585 54.675 96.755 ;
        RECT 54.965 96.585 55.135 96.755 ;
        RECT 55.425 96.585 55.595 96.755 ;
        RECT 55.885 96.585 56.055 96.755 ;
        RECT 56.345 96.585 56.515 96.755 ;
        RECT 56.805 96.585 56.975 96.755 ;
        RECT 57.265 96.585 57.435 96.755 ;
        RECT 57.725 96.585 57.895 96.755 ;
        RECT 58.185 96.585 58.355 96.755 ;
        RECT 58.645 96.585 58.815 96.755 ;
        RECT 59.105 96.585 59.275 96.755 ;
        RECT 59.565 96.585 59.735 96.755 ;
        RECT 60.025 96.585 60.195 96.755 ;
        RECT 60.485 96.585 60.655 96.755 ;
        RECT 60.945 96.585 61.115 96.755 ;
        RECT 61.405 96.585 61.575 96.755 ;
        RECT 61.865 96.585 62.035 96.755 ;
        RECT 62.325 96.585 62.495 96.755 ;
        RECT 62.785 96.585 62.955 96.755 ;
        RECT 63.245 96.585 63.415 96.755 ;
        RECT 63.705 96.585 63.875 96.755 ;
        RECT 64.165 96.585 64.335 96.755 ;
        RECT 64.625 96.585 64.795 96.755 ;
        RECT 65.085 96.585 65.255 96.755 ;
        RECT 65.545 96.585 65.715 96.755 ;
        RECT 66.005 96.585 66.175 96.755 ;
        RECT 66.465 96.585 66.635 96.755 ;
        RECT 66.925 96.585 67.095 96.755 ;
        RECT 67.385 96.585 67.555 96.755 ;
        RECT 67.845 96.585 68.015 96.755 ;
        RECT 68.305 96.585 68.475 96.755 ;
        RECT 68.765 96.585 68.935 96.755 ;
        RECT 69.225 96.585 69.395 96.755 ;
        RECT 69.685 96.585 69.855 96.755 ;
        RECT 70.145 96.585 70.315 96.755 ;
        RECT 70.605 96.585 70.775 96.755 ;
        RECT 71.065 96.585 71.235 96.755 ;
        RECT 71.525 96.585 71.695 96.755 ;
        RECT 71.985 96.585 72.155 96.755 ;
        RECT 72.445 96.585 72.615 96.755 ;
        RECT 72.905 96.585 73.075 96.755 ;
        RECT 73.365 96.585 73.535 96.755 ;
        RECT 73.825 96.585 73.995 96.755 ;
        RECT 74.285 96.585 74.455 96.755 ;
        RECT 74.745 96.585 74.915 96.755 ;
        RECT 75.205 96.585 75.375 96.755 ;
        RECT 75.665 96.585 75.835 96.755 ;
        RECT 76.125 96.585 76.295 96.755 ;
        RECT 76.585 96.585 76.755 96.755 ;
        RECT 77.045 96.585 77.215 96.755 ;
        RECT 77.505 96.585 77.675 96.755 ;
        RECT 77.965 96.585 78.135 96.755 ;
        RECT 78.425 96.585 78.595 96.755 ;
        RECT 78.885 96.585 79.055 96.755 ;
        RECT 79.345 96.585 79.515 96.755 ;
        RECT 79.805 96.585 79.975 96.755 ;
        RECT 80.265 96.585 80.435 96.755 ;
        RECT 80.725 96.585 80.895 96.755 ;
        RECT 81.185 96.585 81.355 96.755 ;
        RECT 81.645 96.585 81.815 96.755 ;
        RECT 82.105 96.585 82.275 96.755 ;
        RECT 82.565 96.585 82.735 96.755 ;
        RECT 83.025 96.585 83.195 96.755 ;
        RECT 83.485 96.585 83.655 96.755 ;
        RECT 83.945 96.585 84.115 96.755 ;
        RECT 84.405 96.585 84.575 96.755 ;
        RECT 84.865 96.585 85.035 96.755 ;
        RECT 85.325 96.585 85.495 96.755 ;
        RECT 85.785 96.585 85.955 96.755 ;
        RECT 86.245 96.585 86.415 96.755 ;
        RECT 86.705 96.585 86.875 96.755 ;
        RECT 87.165 96.585 87.335 96.755 ;
        RECT 87.625 96.585 87.795 96.755 ;
        RECT 88.085 96.585 88.255 96.755 ;
        RECT 88.545 96.585 88.715 96.755 ;
        RECT 89.005 96.585 89.175 96.755 ;
        RECT 89.465 96.585 89.635 96.755 ;
        RECT 89.925 96.585 90.095 96.755 ;
        RECT 90.385 96.585 90.555 96.755 ;
        RECT 90.845 96.585 91.015 96.755 ;
        RECT 91.305 96.585 91.475 96.755 ;
        RECT 91.765 96.585 91.935 96.755 ;
        RECT 92.225 96.585 92.395 96.755 ;
        RECT 92.685 96.585 92.855 96.755 ;
        RECT 93.145 96.585 93.315 96.755 ;
        RECT 93.605 96.585 93.775 96.755 ;
        RECT 94.065 96.585 94.235 96.755 ;
        RECT 94.525 96.585 94.695 96.755 ;
        RECT 94.985 96.585 95.155 96.755 ;
        RECT 95.445 96.585 95.615 96.755 ;
        RECT 95.905 96.585 96.075 96.755 ;
        RECT 96.365 96.585 96.535 96.755 ;
        RECT 96.825 96.585 96.995 96.755 ;
        RECT 97.285 96.585 97.455 96.755 ;
        RECT 97.745 96.585 97.915 96.755 ;
        RECT 98.205 96.585 98.375 96.755 ;
        RECT 98.665 96.585 98.835 96.755 ;
        RECT 99.125 96.585 99.295 96.755 ;
        RECT 99.585 96.585 99.755 96.755 ;
        RECT 100.045 96.585 100.215 96.755 ;
        RECT 100.505 96.585 100.675 96.755 ;
        RECT 100.965 96.585 101.135 96.755 ;
        RECT 101.425 96.585 101.595 96.755 ;
        RECT 101.885 96.585 102.055 96.755 ;
        RECT 102.345 96.585 102.515 96.755 ;
        RECT 102.805 96.585 102.975 96.755 ;
        RECT 103.265 96.585 103.435 96.755 ;
        RECT 103.725 96.585 103.895 96.755 ;
        RECT 104.185 96.585 104.355 96.755 ;
        RECT 104.645 96.585 104.815 96.755 ;
        RECT 105.105 96.585 105.275 96.755 ;
        RECT 105.565 96.585 105.735 96.755 ;
        RECT 106.025 96.585 106.195 96.755 ;
        RECT 106.485 96.585 106.655 96.755 ;
        RECT 106.945 96.585 107.115 96.755 ;
        RECT 107.405 96.585 107.575 96.755 ;
        RECT 107.865 96.585 108.035 96.755 ;
        RECT 108.325 96.585 108.495 96.755 ;
        RECT 108.785 96.585 108.955 96.755 ;
        RECT 109.245 96.585 109.415 96.755 ;
        RECT 109.705 96.585 109.875 96.755 ;
        RECT 110.165 96.585 110.335 96.755 ;
        RECT 110.625 96.585 110.795 96.755 ;
        RECT 111.085 96.585 111.255 96.755 ;
        RECT 111.545 96.585 111.715 96.755 ;
        RECT 112.005 96.585 112.175 96.755 ;
        RECT 112.465 96.585 112.635 96.755 ;
        RECT 112.925 96.585 113.095 96.755 ;
        RECT 113.385 96.585 113.555 96.755 ;
        RECT 113.845 96.585 114.015 96.755 ;
        RECT 114.305 96.585 114.475 96.755 ;
        RECT 114.765 96.585 114.935 96.755 ;
        RECT 115.225 96.585 115.395 96.755 ;
        RECT 115.685 96.585 115.855 96.755 ;
        RECT 116.145 96.585 116.315 96.755 ;
        RECT 116.605 96.585 116.775 96.755 ;
        RECT 117.065 96.585 117.235 96.755 ;
        RECT 117.525 96.585 117.695 96.755 ;
        RECT 117.985 96.585 118.155 96.755 ;
        RECT 118.445 96.585 118.615 96.755 ;
        RECT 118.905 96.585 119.075 96.755 ;
        RECT 119.365 96.585 119.535 96.755 ;
        RECT 119.825 96.585 119.995 96.755 ;
        RECT 120.285 96.585 120.455 96.755 ;
        RECT 120.745 96.585 120.915 96.755 ;
        RECT 121.205 96.585 121.375 96.755 ;
        RECT 121.665 96.585 121.835 96.755 ;
        RECT 122.125 96.585 122.295 96.755 ;
        RECT 122.585 96.585 122.755 96.755 ;
        RECT 123.045 96.585 123.215 96.755 ;
        RECT 123.505 96.585 123.675 96.755 ;
        RECT 123.965 96.585 124.135 96.755 ;
        RECT 124.425 96.585 124.595 96.755 ;
        RECT 124.885 96.585 125.055 96.755 ;
        RECT 125.345 96.585 125.515 96.755 ;
        RECT 125.805 96.585 125.975 96.755 ;
        RECT 126.265 96.585 126.435 96.755 ;
        RECT 126.725 96.585 126.895 96.755 ;
        RECT 127.185 96.585 127.355 96.755 ;
        RECT 127.645 96.585 127.815 96.755 ;
        RECT 128.105 96.585 128.275 96.755 ;
        RECT 128.565 96.585 128.735 96.755 ;
        RECT 129.025 96.585 129.195 96.755 ;
        RECT 129.485 96.585 129.655 96.755 ;
        RECT 129.945 96.585 130.115 96.755 ;
        RECT 130.405 96.585 130.575 96.755 ;
        RECT 130.865 96.585 131.035 96.755 ;
        RECT 131.325 96.585 131.495 96.755 ;
        RECT 131.785 96.585 131.955 96.755 ;
        RECT 132.245 96.585 132.415 96.755 ;
        RECT 132.705 96.585 132.875 96.755 ;
        RECT 133.165 96.585 133.335 96.755 ;
        RECT 133.625 96.585 133.795 96.755 ;
        RECT 134.085 96.585 134.255 96.755 ;
        RECT 134.545 96.585 134.715 96.755 ;
        RECT 135.005 96.585 135.175 96.755 ;
        RECT 135.465 96.585 135.635 96.755 ;
        RECT 135.925 96.585 136.095 96.755 ;
        RECT 136.385 96.585 136.555 96.755 ;
        RECT 136.845 96.585 137.015 96.755 ;
        RECT 137.305 96.585 137.475 96.755 ;
        RECT 137.765 96.585 137.935 96.755 ;
        RECT 138.225 96.585 138.395 96.755 ;
        RECT 138.685 96.585 138.855 96.755 ;
        RECT 139.145 96.585 139.315 96.755 ;
        RECT 139.605 96.585 139.775 96.755 ;
        RECT 140.065 96.585 140.235 96.755 ;
        RECT 140.525 96.585 140.695 96.755 ;
        RECT 140.985 96.585 141.155 96.755 ;
        RECT 141.445 96.585 141.615 96.755 ;
        RECT 141.905 96.585 142.075 96.755 ;
        RECT 142.365 96.585 142.535 96.755 ;
        RECT 142.825 96.585 142.995 96.755 ;
        RECT 143.285 96.585 143.455 96.755 ;
        RECT 143.745 96.585 143.915 96.755 ;
        RECT 144.205 96.585 144.375 96.755 ;
        RECT 144.665 96.585 144.835 96.755 ;
        RECT 145.125 96.585 145.295 96.755 ;
        RECT 145.585 96.585 145.755 96.755 ;
        RECT 146.045 96.585 146.215 96.755 ;
        RECT 146.505 96.585 146.675 96.755 ;
        RECT 146.965 96.585 147.135 96.755 ;
        RECT 147.425 96.585 147.595 96.755 ;
        RECT 147.885 96.585 148.055 96.755 ;
        RECT 148.345 96.585 148.515 96.755 ;
        RECT 148.805 96.585 148.975 96.755 ;
        RECT 149.265 96.585 149.435 96.755 ;
        RECT 149.725 96.585 149.895 96.755 ;
        RECT 150.185 96.585 150.355 96.755 ;
        RECT 11.265 93.865 11.435 94.035 ;
        RECT 11.725 93.865 11.895 94.035 ;
        RECT 12.185 93.865 12.355 94.035 ;
        RECT 12.645 93.865 12.815 94.035 ;
        RECT 13.105 93.865 13.275 94.035 ;
        RECT 13.565 93.865 13.735 94.035 ;
        RECT 14.025 93.865 14.195 94.035 ;
        RECT 14.485 93.865 14.655 94.035 ;
        RECT 14.945 93.865 15.115 94.035 ;
        RECT 15.405 93.865 15.575 94.035 ;
        RECT 15.865 93.865 16.035 94.035 ;
        RECT 16.325 93.865 16.495 94.035 ;
        RECT 16.785 93.865 16.955 94.035 ;
        RECT 17.245 93.865 17.415 94.035 ;
        RECT 17.705 93.865 17.875 94.035 ;
        RECT 18.165 93.865 18.335 94.035 ;
        RECT 18.625 93.865 18.795 94.035 ;
        RECT 19.085 93.865 19.255 94.035 ;
        RECT 19.545 93.865 19.715 94.035 ;
        RECT 20.005 93.865 20.175 94.035 ;
        RECT 20.465 93.865 20.635 94.035 ;
        RECT 20.925 93.865 21.095 94.035 ;
        RECT 21.385 93.865 21.555 94.035 ;
        RECT 21.845 93.865 22.015 94.035 ;
        RECT 22.305 93.865 22.475 94.035 ;
        RECT 22.765 93.865 22.935 94.035 ;
        RECT 23.225 93.865 23.395 94.035 ;
        RECT 23.685 93.865 23.855 94.035 ;
        RECT 24.145 93.865 24.315 94.035 ;
        RECT 24.605 93.865 24.775 94.035 ;
        RECT 25.065 93.865 25.235 94.035 ;
        RECT 25.525 93.865 25.695 94.035 ;
        RECT 25.985 93.865 26.155 94.035 ;
        RECT 26.445 93.865 26.615 94.035 ;
        RECT 26.905 93.865 27.075 94.035 ;
        RECT 27.365 93.865 27.535 94.035 ;
        RECT 27.825 93.865 27.995 94.035 ;
        RECT 28.285 93.865 28.455 94.035 ;
        RECT 28.745 93.865 28.915 94.035 ;
        RECT 29.205 93.865 29.375 94.035 ;
        RECT 29.665 93.865 29.835 94.035 ;
        RECT 30.125 93.865 30.295 94.035 ;
        RECT 30.585 93.865 30.755 94.035 ;
        RECT 31.045 93.865 31.215 94.035 ;
        RECT 31.505 93.865 31.675 94.035 ;
        RECT 31.965 93.865 32.135 94.035 ;
        RECT 32.425 93.865 32.595 94.035 ;
        RECT 32.885 93.865 33.055 94.035 ;
        RECT 33.345 93.865 33.515 94.035 ;
        RECT 33.805 93.865 33.975 94.035 ;
        RECT 34.265 93.865 34.435 94.035 ;
        RECT 34.725 93.865 34.895 94.035 ;
        RECT 35.185 93.865 35.355 94.035 ;
        RECT 35.645 93.865 35.815 94.035 ;
        RECT 36.105 93.865 36.275 94.035 ;
        RECT 36.565 93.865 36.735 94.035 ;
        RECT 37.025 93.865 37.195 94.035 ;
        RECT 37.485 93.865 37.655 94.035 ;
        RECT 37.945 93.865 38.115 94.035 ;
        RECT 38.405 93.865 38.575 94.035 ;
        RECT 38.865 93.865 39.035 94.035 ;
        RECT 39.325 93.865 39.495 94.035 ;
        RECT 39.785 93.865 39.955 94.035 ;
        RECT 40.245 93.865 40.415 94.035 ;
        RECT 40.705 93.865 40.875 94.035 ;
        RECT 41.165 93.865 41.335 94.035 ;
        RECT 41.625 93.865 41.795 94.035 ;
        RECT 42.085 93.865 42.255 94.035 ;
        RECT 42.545 93.865 42.715 94.035 ;
        RECT 43.005 93.865 43.175 94.035 ;
        RECT 43.465 93.865 43.635 94.035 ;
        RECT 43.925 93.865 44.095 94.035 ;
        RECT 44.385 93.865 44.555 94.035 ;
        RECT 44.845 93.865 45.015 94.035 ;
        RECT 45.305 93.865 45.475 94.035 ;
        RECT 45.765 93.865 45.935 94.035 ;
        RECT 46.225 93.865 46.395 94.035 ;
        RECT 46.685 93.865 46.855 94.035 ;
        RECT 47.145 93.865 47.315 94.035 ;
        RECT 47.605 93.865 47.775 94.035 ;
        RECT 48.065 93.865 48.235 94.035 ;
        RECT 48.525 93.865 48.695 94.035 ;
        RECT 48.985 93.865 49.155 94.035 ;
        RECT 49.445 93.865 49.615 94.035 ;
        RECT 49.905 93.865 50.075 94.035 ;
        RECT 50.365 93.865 50.535 94.035 ;
        RECT 50.825 93.865 50.995 94.035 ;
        RECT 51.285 93.865 51.455 94.035 ;
        RECT 51.745 93.865 51.915 94.035 ;
        RECT 52.205 93.865 52.375 94.035 ;
        RECT 52.665 93.865 52.835 94.035 ;
        RECT 53.125 93.865 53.295 94.035 ;
        RECT 53.585 93.865 53.755 94.035 ;
        RECT 54.045 93.865 54.215 94.035 ;
        RECT 54.505 93.865 54.675 94.035 ;
        RECT 54.965 93.865 55.135 94.035 ;
        RECT 55.425 93.865 55.595 94.035 ;
        RECT 55.885 93.865 56.055 94.035 ;
        RECT 56.345 93.865 56.515 94.035 ;
        RECT 56.805 93.865 56.975 94.035 ;
        RECT 57.265 93.865 57.435 94.035 ;
        RECT 57.725 93.865 57.895 94.035 ;
        RECT 58.185 93.865 58.355 94.035 ;
        RECT 58.645 93.865 58.815 94.035 ;
        RECT 59.105 93.865 59.275 94.035 ;
        RECT 59.565 93.865 59.735 94.035 ;
        RECT 60.025 93.865 60.195 94.035 ;
        RECT 60.485 93.865 60.655 94.035 ;
        RECT 60.945 93.865 61.115 94.035 ;
        RECT 61.405 93.865 61.575 94.035 ;
        RECT 61.865 93.865 62.035 94.035 ;
        RECT 62.325 93.865 62.495 94.035 ;
        RECT 62.785 93.865 62.955 94.035 ;
        RECT 63.245 93.865 63.415 94.035 ;
        RECT 63.705 93.865 63.875 94.035 ;
        RECT 64.165 93.865 64.335 94.035 ;
        RECT 64.625 93.865 64.795 94.035 ;
        RECT 65.085 93.865 65.255 94.035 ;
        RECT 65.545 93.865 65.715 94.035 ;
        RECT 66.005 93.865 66.175 94.035 ;
        RECT 66.465 93.865 66.635 94.035 ;
        RECT 66.925 93.865 67.095 94.035 ;
        RECT 67.385 93.865 67.555 94.035 ;
        RECT 67.845 93.865 68.015 94.035 ;
        RECT 68.305 93.865 68.475 94.035 ;
        RECT 68.765 93.865 68.935 94.035 ;
        RECT 69.225 93.865 69.395 94.035 ;
        RECT 69.685 93.865 69.855 94.035 ;
        RECT 70.145 93.865 70.315 94.035 ;
        RECT 70.605 93.865 70.775 94.035 ;
        RECT 71.065 93.865 71.235 94.035 ;
        RECT 71.525 93.865 71.695 94.035 ;
        RECT 71.985 93.865 72.155 94.035 ;
        RECT 72.445 93.865 72.615 94.035 ;
        RECT 72.905 93.865 73.075 94.035 ;
        RECT 73.365 93.865 73.535 94.035 ;
        RECT 73.825 93.865 73.995 94.035 ;
        RECT 74.285 93.865 74.455 94.035 ;
        RECT 74.745 93.865 74.915 94.035 ;
        RECT 75.205 93.865 75.375 94.035 ;
        RECT 75.665 93.865 75.835 94.035 ;
        RECT 76.125 93.865 76.295 94.035 ;
        RECT 76.585 93.865 76.755 94.035 ;
        RECT 77.045 93.865 77.215 94.035 ;
        RECT 77.505 93.865 77.675 94.035 ;
        RECT 77.965 93.865 78.135 94.035 ;
        RECT 78.425 93.865 78.595 94.035 ;
        RECT 78.885 93.865 79.055 94.035 ;
        RECT 79.345 93.865 79.515 94.035 ;
        RECT 79.805 93.865 79.975 94.035 ;
        RECT 80.265 93.865 80.435 94.035 ;
        RECT 80.725 93.865 80.895 94.035 ;
        RECT 81.185 93.865 81.355 94.035 ;
        RECT 81.645 93.865 81.815 94.035 ;
        RECT 82.105 93.865 82.275 94.035 ;
        RECT 82.565 93.865 82.735 94.035 ;
        RECT 83.025 93.865 83.195 94.035 ;
        RECT 83.485 93.865 83.655 94.035 ;
        RECT 83.945 93.865 84.115 94.035 ;
        RECT 84.405 93.865 84.575 94.035 ;
        RECT 84.865 93.865 85.035 94.035 ;
        RECT 85.325 93.865 85.495 94.035 ;
        RECT 85.785 93.865 85.955 94.035 ;
        RECT 86.245 93.865 86.415 94.035 ;
        RECT 86.705 93.865 86.875 94.035 ;
        RECT 87.165 93.865 87.335 94.035 ;
        RECT 87.625 93.865 87.795 94.035 ;
        RECT 88.085 93.865 88.255 94.035 ;
        RECT 88.545 93.865 88.715 94.035 ;
        RECT 89.005 93.865 89.175 94.035 ;
        RECT 89.465 93.865 89.635 94.035 ;
        RECT 89.925 93.865 90.095 94.035 ;
        RECT 90.385 93.865 90.555 94.035 ;
        RECT 90.845 93.865 91.015 94.035 ;
        RECT 91.305 93.865 91.475 94.035 ;
        RECT 91.765 93.865 91.935 94.035 ;
        RECT 92.225 93.865 92.395 94.035 ;
        RECT 92.685 93.865 92.855 94.035 ;
        RECT 93.145 93.865 93.315 94.035 ;
        RECT 93.605 93.865 93.775 94.035 ;
        RECT 94.065 93.865 94.235 94.035 ;
        RECT 94.525 93.865 94.695 94.035 ;
        RECT 94.985 93.865 95.155 94.035 ;
        RECT 95.445 93.865 95.615 94.035 ;
        RECT 95.905 93.865 96.075 94.035 ;
        RECT 96.365 93.865 96.535 94.035 ;
        RECT 96.825 93.865 96.995 94.035 ;
        RECT 97.285 93.865 97.455 94.035 ;
        RECT 97.745 93.865 97.915 94.035 ;
        RECT 98.205 93.865 98.375 94.035 ;
        RECT 98.665 93.865 98.835 94.035 ;
        RECT 99.125 93.865 99.295 94.035 ;
        RECT 99.585 93.865 99.755 94.035 ;
        RECT 100.045 93.865 100.215 94.035 ;
        RECT 100.505 93.865 100.675 94.035 ;
        RECT 100.965 93.865 101.135 94.035 ;
        RECT 101.425 93.865 101.595 94.035 ;
        RECT 101.885 93.865 102.055 94.035 ;
        RECT 102.345 93.865 102.515 94.035 ;
        RECT 102.805 93.865 102.975 94.035 ;
        RECT 103.265 93.865 103.435 94.035 ;
        RECT 103.725 93.865 103.895 94.035 ;
        RECT 104.185 93.865 104.355 94.035 ;
        RECT 104.645 93.865 104.815 94.035 ;
        RECT 105.105 93.865 105.275 94.035 ;
        RECT 105.565 93.865 105.735 94.035 ;
        RECT 106.025 93.865 106.195 94.035 ;
        RECT 106.485 93.865 106.655 94.035 ;
        RECT 106.945 93.865 107.115 94.035 ;
        RECT 107.405 93.865 107.575 94.035 ;
        RECT 107.865 93.865 108.035 94.035 ;
        RECT 108.325 93.865 108.495 94.035 ;
        RECT 108.785 93.865 108.955 94.035 ;
        RECT 109.245 93.865 109.415 94.035 ;
        RECT 109.705 93.865 109.875 94.035 ;
        RECT 110.165 93.865 110.335 94.035 ;
        RECT 110.625 93.865 110.795 94.035 ;
        RECT 111.085 93.865 111.255 94.035 ;
        RECT 111.545 93.865 111.715 94.035 ;
        RECT 112.005 93.865 112.175 94.035 ;
        RECT 112.465 93.865 112.635 94.035 ;
        RECT 112.925 93.865 113.095 94.035 ;
        RECT 113.385 93.865 113.555 94.035 ;
        RECT 113.845 93.865 114.015 94.035 ;
        RECT 114.305 93.865 114.475 94.035 ;
        RECT 114.765 93.865 114.935 94.035 ;
        RECT 115.225 93.865 115.395 94.035 ;
        RECT 115.685 93.865 115.855 94.035 ;
        RECT 116.145 93.865 116.315 94.035 ;
        RECT 116.605 93.865 116.775 94.035 ;
        RECT 117.065 93.865 117.235 94.035 ;
        RECT 117.525 93.865 117.695 94.035 ;
        RECT 117.985 93.865 118.155 94.035 ;
        RECT 118.445 93.865 118.615 94.035 ;
        RECT 118.905 93.865 119.075 94.035 ;
        RECT 119.365 93.865 119.535 94.035 ;
        RECT 119.825 93.865 119.995 94.035 ;
        RECT 120.285 93.865 120.455 94.035 ;
        RECT 120.745 93.865 120.915 94.035 ;
        RECT 121.205 93.865 121.375 94.035 ;
        RECT 121.665 93.865 121.835 94.035 ;
        RECT 122.125 93.865 122.295 94.035 ;
        RECT 122.585 93.865 122.755 94.035 ;
        RECT 123.045 93.865 123.215 94.035 ;
        RECT 123.505 93.865 123.675 94.035 ;
        RECT 123.965 93.865 124.135 94.035 ;
        RECT 124.425 93.865 124.595 94.035 ;
        RECT 124.885 93.865 125.055 94.035 ;
        RECT 125.345 93.865 125.515 94.035 ;
        RECT 125.805 93.865 125.975 94.035 ;
        RECT 126.265 93.865 126.435 94.035 ;
        RECT 126.725 93.865 126.895 94.035 ;
        RECT 127.185 93.865 127.355 94.035 ;
        RECT 127.645 93.865 127.815 94.035 ;
        RECT 128.105 93.865 128.275 94.035 ;
        RECT 128.565 93.865 128.735 94.035 ;
        RECT 129.025 93.865 129.195 94.035 ;
        RECT 129.485 93.865 129.655 94.035 ;
        RECT 129.945 93.865 130.115 94.035 ;
        RECT 130.405 93.865 130.575 94.035 ;
        RECT 130.865 93.865 131.035 94.035 ;
        RECT 131.325 93.865 131.495 94.035 ;
        RECT 131.785 93.865 131.955 94.035 ;
        RECT 132.245 93.865 132.415 94.035 ;
        RECT 132.705 93.865 132.875 94.035 ;
        RECT 133.165 93.865 133.335 94.035 ;
        RECT 133.625 93.865 133.795 94.035 ;
        RECT 134.085 93.865 134.255 94.035 ;
        RECT 134.545 93.865 134.715 94.035 ;
        RECT 135.005 93.865 135.175 94.035 ;
        RECT 135.465 93.865 135.635 94.035 ;
        RECT 135.925 93.865 136.095 94.035 ;
        RECT 136.385 93.865 136.555 94.035 ;
        RECT 136.845 93.865 137.015 94.035 ;
        RECT 137.305 93.865 137.475 94.035 ;
        RECT 137.765 93.865 137.935 94.035 ;
        RECT 138.225 93.865 138.395 94.035 ;
        RECT 138.685 93.865 138.855 94.035 ;
        RECT 139.145 93.865 139.315 94.035 ;
        RECT 139.605 93.865 139.775 94.035 ;
        RECT 140.065 93.865 140.235 94.035 ;
        RECT 140.525 93.865 140.695 94.035 ;
        RECT 140.985 93.865 141.155 94.035 ;
        RECT 141.445 93.865 141.615 94.035 ;
        RECT 141.905 93.865 142.075 94.035 ;
        RECT 142.365 93.865 142.535 94.035 ;
        RECT 142.825 93.865 142.995 94.035 ;
        RECT 143.285 93.865 143.455 94.035 ;
        RECT 143.745 93.865 143.915 94.035 ;
        RECT 144.205 93.865 144.375 94.035 ;
        RECT 144.665 93.865 144.835 94.035 ;
        RECT 145.125 93.865 145.295 94.035 ;
        RECT 145.585 93.865 145.755 94.035 ;
        RECT 146.045 93.865 146.215 94.035 ;
        RECT 146.505 93.865 146.675 94.035 ;
        RECT 146.965 93.865 147.135 94.035 ;
        RECT 147.425 93.865 147.595 94.035 ;
        RECT 147.885 93.865 148.055 94.035 ;
        RECT 148.345 93.865 148.515 94.035 ;
        RECT 148.805 93.865 148.975 94.035 ;
        RECT 149.265 93.865 149.435 94.035 ;
        RECT 149.725 93.865 149.895 94.035 ;
        RECT 150.185 93.865 150.355 94.035 ;
        RECT 11.265 91.145 11.435 91.315 ;
        RECT 11.725 91.145 11.895 91.315 ;
        RECT 12.185 91.145 12.355 91.315 ;
        RECT 12.645 91.145 12.815 91.315 ;
        RECT 13.105 91.145 13.275 91.315 ;
        RECT 13.565 91.145 13.735 91.315 ;
        RECT 14.025 91.145 14.195 91.315 ;
        RECT 14.485 91.145 14.655 91.315 ;
        RECT 14.945 91.145 15.115 91.315 ;
        RECT 15.405 91.145 15.575 91.315 ;
        RECT 15.865 91.145 16.035 91.315 ;
        RECT 16.325 91.145 16.495 91.315 ;
        RECT 16.785 91.145 16.955 91.315 ;
        RECT 17.245 91.145 17.415 91.315 ;
        RECT 17.705 91.145 17.875 91.315 ;
        RECT 18.165 91.145 18.335 91.315 ;
        RECT 18.625 91.145 18.795 91.315 ;
        RECT 19.085 91.145 19.255 91.315 ;
        RECT 19.545 91.145 19.715 91.315 ;
        RECT 20.005 91.145 20.175 91.315 ;
        RECT 20.465 91.145 20.635 91.315 ;
        RECT 20.925 91.145 21.095 91.315 ;
        RECT 21.385 91.145 21.555 91.315 ;
        RECT 21.845 91.145 22.015 91.315 ;
        RECT 22.305 91.145 22.475 91.315 ;
        RECT 22.765 91.145 22.935 91.315 ;
        RECT 23.225 91.145 23.395 91.315 ;
        RECT 23.685 91.145 23.855 91.315 ;
        RECT 24.145 91.145 24.315 91.315 ;
        RECT 24.605 91.145 24.775 91.315 ;
        RECT 25.065 91.145 25.235 91.315 ;
        RECT 25.525 91.145 25.695 91.315 ;
        RECT 25.985 91.145 26.155 91.315 ;
        RECT 26.445 91.145 26.615 91.315 ;
        RECT 26.905 91.145 27.075 91.315 ;
        RECT 27.365 91.145 27.535 91.315 ;
        RECT 27.825 91.145 27.995 91.315 ;
        RECT 28.285 91.145 28.455 91.315 ;
        RECT 28.745 91.145 28.915 91.315 ;
        RECT 29.205 91.145 29.375 91.315 ;
        RECT 29.665 91.145 29.835 91.315 ;
        RECT 30.125 91.145 30.295 91.315 ;
        RECT 30.585 91.145 30.755 91.315 ;
        RECT 31.045 91.145 31.215 91.315 ;
        RECT 31.505 91.145 31.675 91.315 ;
        RECT 31.965 91.145 32.135 91.315 ;
        RECT 32.425 91.145 32.595 91.315 ;
        RECT 32.885 91.145 33.055 91.315 ;
        RECT 33.345 91.145 33.515 91.315 ;
        RECT 33.805 91.145 33.975 91.315 ;
        RECT 34.265 91.145 34.435 91.315 ;
        RECT 34.725 91.145 34.895 91.315 ;
        RECT 35.185 91.145 35.355 91.315 ;
        RECT 35.645 91.145 35.815 91.315 ;
        RECT 36.105 91.145 36.275 91.315 ;
        RECT 36.565 91.145 36.735 91.315 ;
        RECT 37.025 91.145 37.195 91.315 ;
        RECT 37.485 91.145 37.655 91.315 ;
        RECT 37.945 91.145 38.115 91.315 ;
        RECT 38.405 91.145 38.575 91.315 ;
        RECT 38.865 91.145 39.035 91.315 ;
        RECT 39.325 91.145 39.495 91.315 ;
        RECT 39.785 91.145 39.955 91.315 ;
        RECT 40.245 91.145 40.415 91.315 ;
        RECT 40.705 91.145 40.875 91.315 ;
        RECT 41.165 91.145 41.335 91.315 ;
        RECT 41.625 91.145 41.795 91.315 ;
        RECT 42.085 91.145 42.255 91.315 ;
        RECT 42.545 91.145 42.715 91.315 ;
        RECT 43.005 91.145 43.175 91.315 ;
        RECT 43.465 91.145 43.635 91.315 ;
        RECT 43.925 91.145 44.095 91.315 ;
        RECT 44.385 91.145 44.555 91.315 ;
        RECT 44.845 91.145 45.015 91.315 ;
        RECT 45.305 91.145 45.475 91.315 ;
        RECT 45.765 91.145 45.935 91.315 ;
        RECT 46.225 91.145 46.395 91.315 ;
        RECT 46.685 91.145 46.855 91.315 ;
        RECT 47.145 91.145 47.315 91.315 ;
        RECT 47.605 91.145 47.775 91.315 ;
        RECT 48.065 91.145 48.235 91.315 ;
        RECT 48.525 91.145 48.695 91.315 ;
        RECT 48.985 91.145 49.155 91.315 ;
        RECT 49.445 91.145 49.615 91.315 ;
        RECT 49.905 91.145 50.075 91.315 ;
        RECT 50.365 91.145 50.535 91.315 ;
        RECT 50.825 91.145 50.995 91.315 ;
        RECT 51.285 91.145 51.455 91.315 ;
        RECT 51.745 91.145 51.915 91.315 ;
        RECT 52.205 91.145 52.375 91.315 ;
        RECT 52.665 91.145 52.835 91.315 ;
        RECT 53.125 91.145 53.295 91.315 ;
        RECT 53.585 91.145 53.755 91.315 ;
        RECT 54.045 91.145 54.215 91.315 ;
        RECT 54.505 91.145 54.675 91.315 ;
        RECT 54.965 91.145 55.135 91.315 ;
        RECT 55.425 91.145 55.595 91.315 ;
        RECT 55.885 91.145 56.055 91.315 ;
        RECT 56.345 91.145 56.515 91.315 ;
        RECT 56.805 91.145 56.975 91.315 ;
        RECT 57.265 91.145 57.435 91.315 ;
        RECT 57.725 91.145 57.895 91.315 ;
        RECT 58.185 91.145 58.355 91.315 ;
        RECT 58.645 91.145 58.815 91.315 ;
        RECT 59.105 91.145 59.275 91.315 ;
        RECT 59.565 91.145 59.735 91.315 ;
        RECT 60.025 91.145 60.195 91.315 ;
        RECT 60.485 91.145 60.655 91.315 ;
        RECT 60.945 91.145 61.115 91.315 ;
        RECT 61.405 91.145 61.575 91.315 ;
        RECT 61.865 91.145 62.035 91.315 ;
        RECT 62.325 91.145 62.495 91.315 ;
        RECT 62.785 91.145 62.955 91.315 ;
        RECT 63.245 91.145 63.415 91.315 ;
        RECT 63.705 91.145 63.875 91.315 ;
        RECT 64.165 91.145 64.335 91.315 ;
        RECT 64.625 91.145 64.795 91.315 ;
        RECT 65.085 91.145 65.255 91.315 ;
        RECT 65.545 91.145 65.715 91.315 ;
        RECT 66.005 91.145 66.175 91.315 ;
        RECT 66.465 91.145 66.635 91.315 ;
        RECT 66.925 91.145 67.095 91.315 ;
        RECT 67.385 91.145 67.555 91.315 ;
        RECT 67.845 91.145 68.015 91.315 ;
        RECT 68.305 91.145 68.475 91.315 ;
        RECT 68.765 91.145 68.935 91.315 ;
        RECT 69.225 91.145 69.395 91.315 ;
        RECT 69.685 91.145 69.855 91.315 ;
        RECT 70.145 91.145 70.315 91.315 ;
        RECT 70.605 91.145 70.775 91.315 ;
        RECT 71.065 91.145 71.235 91.315 ;
        RECT 71.525 91.145 71.695 91.315 ;
        RECT 71.985 91.145 72.155 91.315 ;
        RECT 72.445 91.145 72.615 91.315 ;
        RECT 72.905 91.145 73.075 91.315 ;
        RECT 73.365 91.145 73.535 91.315 ;
        RECT 73.825 91.145 73.995 91.315 ;
        RECT 74.285 91.145 74.455 91.315 ;
        RECT 74.745 91.145 74.915 91.315 ;
        RECT 75.205 91.145 75.375 91.315 ;
        RECT 75.665 91.145 75.835 91.315 ;
        RECT 76.125 91.145 76.295 91.315 ;
        RECT 76.585 91.145 76.755 91.315 ;
        RECT 77.045 91.145 77.215 91.315 ;
        RECT 77.505 91.145 77.675 91.315 ;
        RECT 77.965 91.145 78.135 91.315 ;
        RECT 78.425 91.145 78.595 91.315 ;
        RECT 78.885 91.145 79.055 91.315 ;
        RECT 79.345 91.145 79.515 91.315 ;
        RECT 79.805 91.145 79.975 91.315 ;
        RECT 80.265 91.145 80.435 91.315 ;
        RECT 80.725 91.145 80.895 91.315 ;
        RECT 81.185 91.145 81.355 91.315 ;
        RECT 81.645 91.145 81.815 91.315 ;
        RECT 82.105 91.145 82.275 91.315 ;
        RECT 82.565 91.145 82.735 91.315 ;
        RECT 83.025 91.145 83.195 91.315 ;
        RECT 83.485 91.145 83.655 91.315 ;
        RECT 83.945 91.145 84.115 91.315 ;
        RECT 84.405 91.145 84.575 91.315 ;
        RECT 84.865 91.145 85.035 91.315 ;
        RECT 85.325 91.145 85.495 91.315 ;
        RECT 85.785 91.145 85.955 91.315 ;
        RECT 86.245 91.145 86.415 91.315 ;
        RECT 86.705 91.145 86.875 91.315 ;
        RECT 87.165 91.145 87.335 91.315 ;
        RECT 87.625 91.145 87.795 91.315 ;
        RECT 88.085 91.145 88.255 91.315 ;
        RECT 88.545 91.145 88.715 91.315 ;
        RECT 89.005 91.145 89.175 91.315 ;
        RECT 89.465 91.145 89.635 91.315 ;
        RECT 89.925 91.145 90.095 91.315 ;
        RECT 90.385 91.145 90.555 91.315 ;
        RECT 90.845 91.145 91.015 91.315 ;
        RECT 91.305 91.145 91.475 91.315 ;
        RECT 91.765 91.145 91.935 91.315 ;
        RECT 92.225 91.145 92.395 91.315 ;
        RECT 92.685 91.145 92.855 91.315 ;
        RECT 93.145 91.145 93.315 91.315 ;
        RECT 93.605 91.145 93.775 91.315 ;
        RECT 94.065 91.145 94.235 91.315 ;
        RECT 94.525 91.145 94.695 91.315 ;
        RECT 94.985 91.145 95.155 91.315 ;
        RECT 95.445 91.145 95.615 91.315 ;
        RECT 95.905 91.145 96.075 91.315 ;
        RECT 96.365 91.145 96.535 91.315 ;
        RECT 96.825 91.145 96.995 91.315 ;
        RECT 97.285 91.145 97.455 91.315 ;
        RECT 97.745 91.145 97.915 91.315 ;
        RECT 98.205 91.145 98.375 91.315 ;
        RECT 98.665 91.145 98.835 91.315 ;
        RECT 99.125 91.145 99.295 91.315 ;
        RECT 99.585 91.145 99.755 91.315 ;
        RECT 100.045 91.145 100.215 91.315 ;
        RECT 100.505 91.145 100.675 91.315 ;
        RECT 100.965 91.145 101.135 91.315 ;
        RECT 101.425 91.145 101.595 91.315 ;
        RECT 101.885 91.145 102.055 91.315 ;
        RECT 102.345 91.145 102.515 91.315 ;
        RECT 102.805 91.145 102.975 91.315 ;
        RECT 103.265 91.145 103.435 91.315 ;
        RECT 103.725 91.145 103.895 91.315 ;
        RECT 104.185 91.145 104.355 91.315 ;
        RECT 104.645 91.145 104.815 91.315 ;
        RECT 105.105 91.145 105.275 91.315 ;
        RECT 105.565 91.145 105.735 91.315 ;
        RECT 106.025 91.145 106.195 91.315 ;
        RECT 106.485 91.145 106.655 91.315 ;
        RECT 106.945 91.145 107.115 91.315 ;
        RECT 107.405 91.145 107.575 91.315 ;
        RECT 107.865 91.145 108.035 91.315 ;
        RECT 108.325 91.145 108.495 91.315 ;
        RECT 108.785 91.145 108.955 91.315 ;
        RECT 109.245 91.145 109.415 91.315 ;
        RECT 109.705 91.145 109.875 91.315 ;
        RECT 110.165 91.145 110.335 91.315 ;
        RECT 110.625 91.145 110.795 91.315 ;
        RECT 111.085 91.145 111.255 91.315 ;
        RECT 111.545 91.145 111.715 91.315 ;
        RECT 112.005 91.145 112.175 91.315 ;
        RECT 112.465 91.145 112.635 91.315 ;
        RECT 112.925 91.145 113.095 91.315 ;
        RECT 113.385 91.145 113.555 91.315 ;
        RECT 113.845 91.145 114.015 91.315 ;
        RECT 114.305 91.145 114.475 91.315 ;
        RECT 114.765 91.145 114.935 91.315 ;
        RECT 115.225 91.145 115.395 91.315 ;
        RECT 115.685 91.145 115.855 91.315 ;
        RECT 116.145 91.145 116.315 91.315 ;
        RECT 116.605 91.145 116.775 91.315 ;
        RECT 117.065 91.145 117.235 91.315 ;
        RECT 117.525 91.145 117.695 91.315 ;
        RECT 117.985 91.145 118.155 91.315 ;
        RECT 118.445 91.145 118.615 91.315 ;
        RECT 118.905 91.145 119.075 91.315 ;
        RECT 119.365 91.145 119.535 91.315 ;
        RECT 119.825 91.145 119.995 91.315 ;
        RECT 120.285 91.145 120.455 91.315 ;
        RECT 120.745 91.145 120.915 91.315 ;
        RECT 121.205 91.145 121.375 91.315 ;
        RECT 121.665 91.145 121.835 91.315 ;
        RECT 122.125 91.145 122.295 91.315 ;
        RECT 122.585 91.145 122.755 91.315 ;
        RECT 123.045 91.145 123.215 91.315 ;
        RECT 123.505 91.145 123.675 91.315 ;
        RECT 123.965 91.145 124.135 91.315 ;
        RECT 124.425 91.145 124.595 91.315 ;
        RECT 124.885 91.145 125.055 91.315 ;
        RECT 125.345 91.145 125.515 91.315 ;
        RECT 125.805 91.145 125.975 91.315 ;
        RECT 126.265 91.145 126.435 91.315 ;
        RECT 126.725 91.145 126.895 91.315 ;
        RECT 127.185 91.145 127.355 91.315 ;
        RECT 127.645 91.145 127.815 91.315 ;
        RECT 128.105 91.145 128.275 91.315 ;
        RECT 128.565 91.145 128.735 91.315 ;
        RECT 129.025 91.145 129.195 91.315 ;
        RECT 129.485 91.145 129.655 91.315 ;
        RECT 129.945 91.145 130.115 91.315 ;
        RECT 130.405 91.145 130.575 91.315 ;
        RECT 130.865 91.145 131.035 91.315 ;
        RECT 131.325 91.145 131.495 91.315 ;
        RECT 131.785 91.145 131.955 91.315 ;
        RECT 132.245 91.145 132.415 91.315 ;
        RECT 132.705 91.145 132.875 91.315 ;
        RECT 133.165 91.145 133.335 91.315 ;
        RECT 133.625 91.145 133.795 91.315 ;
        RECT 134.085 91.145 134.255 91.315 ;
        RECT 134.545 91.145 134.715 91.315 ;
        RECT 135.005 91.145 135.175 91.315 ;
        RECT 135.465 91.145 135.635 91.315 ;
        RECT 135.925 91.145 136.095 91.315 ;
        RECT 136.385 91.145 136.555 91.315 ;
        RECT 136.845 91.145 137.015 91.315 ;
        RECT 137.305 91.145 137.475 91.315 ;
        RECT 137.765 91.145 137.935 91.315 ;
        RECT 138.225 91.145 138.395 91.315 ;
        RECT 138.685 91.145 138.855 91.315 ;
        RECT 139.145 91.145 139.315 91.315 ;
        RECT 139.605 91.145 139.775 91.315 ;
        RECT 140.065 91.145 140.235 91.315 ;
        RECT 140.525 91.145 140.695 91.315 ;
        RECT 140.985 91.145 141.155 91.315 ;
        RECT 141.445 91.145 141.615 91.315 ;
        RECT 141.905 91.145 142.075 91.315 ;
        RECT 142.365 91.145 142.535 91.315 ;
        RECT 142.825 91.145 142.995 91.315 ;
        RECT 143.285 91.145 143.455 91.315 ;
        RECT 143.745 91.145 143.915 91.315 ;
        RECT 144.205 91.145 144.375 91.315 ;
        RECT 144.665 91.145 144.835 91.315 ;
        RECT 145.125 91.145 145.295 91.315 ;
        RECT 145.585 91.145 145.755 91.315 ;
        RECT 146.045 91.145 146.215 91.315 ;
        RECT 146.505 91.145 146.675 91.315 ;
        RECT 146.965 91.145 147.135 91.315 ;
        RECT 147.425 91.145 147.595 91.315 ;
        RECT 147.885 91.145 148.055 91.315 ;
        RECT 148.345 91.145 148.515 91.315 ;
        RECT 148.805 91.145 148.975 91.315 ;
        RECT 149.265 91.145 149.435 91.315 ;
        RECT 149.725 91.145 149.895 91.315 ;
        RECT 150.185 91.145 150.355 91.315 ;
        RECT 11.265 88.425 11.435 88.595 ;
        RECT 11.725 88.425 11.895 88.595 ;
        RECT 12.185 88.425 12.355 88.595 ;
        RECT 12.645 88.425 12.815 88.595 ;
        RECT 13.105 88.425 13.275 88.595 ;
        RECT 13.565 88.425 13.735 88.595 ;
        RECT 14.025 88.425 14.195 88.595 ;
        RECT 14.485 88.425 14.655 88.595 ;
        RECT 14.945 88.425 15.115 88.595 ;
        RECT 15.405 88.425 15.575 88.595 ;
        RECT 15.865 88.425 16.035 88.595 ;
        RECT 16.325 88.425 16.495 88.595 ;
        RECT 16.785 88.425 16.955 88.595 ;
        RECT 17.245 88.425 17.415 88.595 ;
        RECT 17.705 88.425 17.875 88.595 ;
        RECT 18.165 88.425 18.335 88.595 ;
        RECT 18.625 88.425 18.795 88.595 ;
        RECT 19.085 88.425 19.255 88.595 ;
        RECT 19.545 88.425 19.715 88.595 ;
        RECT 20.005 88.425 20.175 88.595 ;
        RECT 20.465 88.425 20.635 88.595 ;
        RECT 20.925 88.425 21.095 88.595 ;
        RECT 21.385 88.425 21.555 88.595 ;
        RECT 21.845 88.425 22.015 88.595 ;
        RECT 22.305 88.425 22.475 88.595 ;
        RECT 22.765 88.425 22.935 88.595 ;
        RECT 23.225 88.425 23.395 88.595 ;
        RECT 23.685 88.425 23.855 88.595 ;
        RECT 24.145 88.425 24.315 88.595 ;
        RECT 24.605 88.425 24.775 88.595 ;
        RECT 25.065 88.425 25.235 88.595 ;
        RECT 25.525 88.425 25.695 88.595 ;
        RECT 25.985 88.425 26.155 88.595 ;
        RECT 26.445 88.425 26.615 88.595 ;
        RECT 26.905 88.425 27.075 88.595 ;
        RECT 27.365 88.425 27.535 88.595 ;
        RECT 27.825 88.425 27.995 88.595 ;
        RECT 28.285 88.425 28.455 88.595 ;
        RECT 28.745 88.425 28.915 88.595 ;
        RECT 29.205 88.425 29.375 88.595 ;
        RECT 29.665 88.425 29.835 88.595 ;
        RECT 30.125 88.425 30.295 88.595 ;
        RECT 30.585 88.425 30.755 88.595 ;
        RECT 31.045 88.425 31.215 88.595 ;
        RECT 31.505 88.425 31.675 88.595 ;
        RECT 31.965 88.425 32.135 88.595 ;
        RECT 32.425 88.425 32.595 88.595 ;
        RECT 32.885 88.425 33.055 88.595 ;
        RECT 33.345 88.425 33.515 88.595 ;
        RECT 33.805 88.425 33.975 88.595 ;
        RECT 34.265 88.425 34.435 88.595 ;
        RECT 34.725 88.425 34.895 88.595 ;
        RECT 35.185 88.425 35.355 88.595 ;
        RECT 35.645 88.425 35.815 88.595 ;
        RECT 36.105 88.425 36.275 88.595 ;
        RECT 36.565 88.425 36.735 88.595 ;
        RECT 37.025 88.425 37.195 88.595 ;
        RECT 37.485 88.425 37.655 88.595 ;
        RECT 37.945 88.425 38.115 88.595 ;
        RECT 38.405 88.425 38.575 88.595 ;
        RECT 38.865 88.425 39.035 88.595 ;
        RECT 39.325 88.425 39.495 88.595 ;
        RECT 39.785 88.425 39.955 88.595 ;
        RECT 40.245 88.425 40.415 88.595 ;
        RECT 40.705 88.425 40.875 88.595 ;
        RECT 41.165 88.425 41.335 88.595 ;
        RECT 41.625 88.425 41.795 88.595 ;
        RECT 42.085 88.425 42.255 88.595 ;
        RECT 42.545 88.425 42.715 88.595 ;
        RECT 43.005 88.425 43.175 88.595 ;
        RECT 43.465 88.425 43.635 88.595 ;
        RECT 43.925 88.425 44.095 88.595 ;
        RECT 44.385 88.425 44.555 88.595 ;
        RECT 44.845 88.425 45.015 88.595 ;
        RECT 45.305 88.425 45.475 88.595 ;
        RECT 45.765 88.425 45.935 88.595 ;
        RECT 46.225 88.425 46.395 88.595 ;
        RECT 46.685 88.425 46.855 88.595 ;
        RECT 47.145 88.425 47.315 88.595 ;
        RECT 47.605 88.425 47.775 88.595 ;
        RECT 48.065 88.425 48.235 88.595 ;
        RECT 48.525 88.425 48.695 88.595 ;
        RECT 48.985 88.425 49.155 88.595 ;
        RECT 49.445 88.425 49.615 88.595 ;
        RECT 49.905 88.425 50.075 88.595 ;
        RECT 50.365 88.425 50.535 88.595 ;
        RECT 50.825 88.425 50.995 88.595 ;
        RECT 51.285 88.425 51.455 88.595 ;
        RECT 51.745 88.425 51.915 88.595 ;
        RECT 52.205 88.425 52.375 88.595 ;
        RECT 52.665 88.425 52.835 88.595 ;
        RECT 53.125 88.425 53.295 88.595 ;
        RECT 53.585 88.425 53.755 88.595 ;
        RECT 54.045 88.425 54.215 88.595 ;
        RECT 54.505 88.425 54.675 88.595 ;
        RECT 54.965 88.425 55.135 88.595 ;
        RECT 55.425 88.425 55.595 88.595 ;
        RECT 55.885 88.425 56.055 88.595 ;
        RECT 56.345 88.425 56.515 88.595 ;
        RECT 56.805 88.425 56.975 88.595 ;
        RECT 57.265 88.425 57.435 88.595 ;
        RECT 57.725 88.425 57.895 88.595 ;
        RECT 58.185 88.425 58.355 88.595 ;
        RECT 58.645 88.425 58.815 88.595 ;
        RECT 59.105 88.425 59.275 88.595 ;
        RECT 59.565 88.425 59.735 88.595 ;
        RECT 60.025 88.425 60.195 88.595 ;
        RECT 60.485 88.425 60.655 88.595 ;
        RECT 60.945 88.425 61.115 88.595 ;
        RECT 61.405 88.425 61.575 88.595 ;
        RECT 61.865 88.425 62.035 88.595 ;
        RECT 62.325 88.425 62.495 88.595 ;
        RECT 62.785 88.425 62.955 88.595 ;
        RECT 63.245 88.425 63.415 88.595 ;
        RECT 63.705 88.425 63.875 88.595 ;
        RECT 64.165 88.425 64.335 88.595 ;
        RECT 64.625 88.425 64.795 88.595 ;
        RECT 65.085 88.425 65.255 88.595 ;
        RECT 65.545 88.425 65.715 88.595 ;
        RECT 66.005 88.425 66.175 88.595 ;
        RECT 66.465 88.425 66.635 88.595 ;
        RECT 66.925 88.425 67.095 88.595 ;
        RECT 67.385 88.425 67.555 88.595 ;
        RECT 67.845 88.425 68.015 88.595 ;
        RECT 68.305 88.425 68.475 88.595 ;
        RECT 68.765 88.425 68.935 88.595 ;
        RECT 69.225 88.425 69.395 88.595 ;
        RECT 69.685 88.425 69.855 88.595 ;
        RECT 70.145 88.425 70.315 88.595 ;
        RECT 70.605 88.425 70.775 88.595 ;
        RECT 71.065 88.425 71.235 88.595 ;
        RECT 71.525 88.425 71.695 88.595 ;
        RECT 71.985 88.425 72.155 88.595 ;
        RECT 72.445 88.425 72.615 88.595 ;
        RECT 72.905 88.425 73.075 88.595 ;
        RECT 73.365 88.425 73.535 88.595 ;
        RECT 73.825 88.425 73.995 88.595 ;
        RECT 74.285 88.425 74.455 88.595 ;
        RECT 74.745 88.425 74.915 88.595 ;
        RECT 75.205 88.425 75.375 88.595 ;
        RECT 75.665 88.425 75.835 88.595 ;
        RECT 76.125 88.425 76.295 88.595 ;
        RECT 76.585 88.425 76.755 88.595 ;
        RECT 77.045 88.425 77.215 88.595 ;
        RECT 77.505 88.425 77.675 88.595 ;
        RECT 77.965 88.425 78.135 88.595 ;
        RECT 78.425 88.425 78.595 88.595 ;
        RECT 78.885 88.425 79.055 88.595 ;
        RECT 79.345 88.425 79.515 88.595 ;
        RECT 79.805 88.425 79.975 88.595 ;
        RECT 80.265 88.425 80.435 88.595 ;
        RECT 80.725 88.425 80.895 88.595 ;
        RECT 81.185 88.425 81.355 88.595 ;
        RECT 81.645 88.425 81.815 88.595 ;
        RECT 82.105 88.425 82.275 88.595 ;
        RECT 82.565 88.425 82.735 88.595 ;
        RECT 83.025 88.425 83.195 88.595 ;
        RECT 83.485 88.425 83.655 88.595 ;
        RECT 83.945 88.425 84.115 88.595 ;
        RECT 84.405 88.425 84.575 88.595 ;
        RECT 84.865 88.425 85.035 88.595 ;
        RECT 85.325 88.425 85.495 88.595 ;
        RECT 85.785 88.425 85.955 88.595 ;
        RECT 86.245 88.425 86.415 88.595 ;
        RECT 86.705 88.425 86.875 88.595 ;
        RECT 87.165 88.425 87.335 88.595 ;
        RECT 87.625 88.425 87.795 88.595 ;
        RECT 88.085 88.425 88.255 88.595 ;
        RECT 88.545 88.425 88.715 88.595 ;
        RECT 89.005 88.425 89.175 88.595 ;
        RECT 89.465 88.425 89.635 88.595 ;
        RECT 89.925 88.425 90.095 88.595 ;
        RECT 90.385 88.425 90.555 88.595 ;
        RECT 90.845 88.425 91.015 88.595 ;
        RECT 91.305 88.425 91.475 88.595 ;
        RECT 91.765 88.425 91.935 88.595 ;
        RECT 92.225 88.425 92.395 88.595 ;
        RECT 92.685 88.425 92.855 88.595 ;
        RECT 93.145 88.425 93.315 88.595 ;
        RECT 93.605 88.425 93.775 88.595 ;
        RECT 94.065 88.425 94.235 88.595 ;
        RECT 94.525 88.425 94.695 88.595 ;
        RECT 94.985 88.425 95.155 88.595 ;
        RECT 95.445 88.425 95.615 88.595 ;
        RECT 95.905 88.425 96.075 88.595 ;
        RECT 96.365 88.425 96.535 88.595 ;
        RECT 96.825 88.425 96.995 88.595 ;
        RECT 97.285 88.425 97.455 88.595 ;
        RECT 97.745 88.425 97.915 88.595 ;
        RECT 98.205 88.425 98.375 88.595 ;
        RECT 98.665 88.425 98.835 88.595 ;
        RECT 99.125 88.425 99.295 88.595 ;
        RECT 99.585 88.425 99.755 88.595 ;
        RECT 100.045 88.425 100.215 88.595 ;
        RECT 100.505 88.425 100.675 88.595 ;
        RECT 100.965 88.425 101.135 88.595 ;
        RECT 101.425 88.425 101.595 88.595 ;
        RECT 101.885 88.425 102.055 88.595 ;
        RECT 102.345 88.425 102.515 88.595 ;
        RECT 102.805 88.425 102.975 88.595 ;
        RECT 103.265 88.425 103.435 88.595 ;
        RECT 103.725 88.425 103.895 88.595 ;
        RECT 104.185 88.425 104.355 88.595 ;
        RECT 104.645 88.425 104.815 88.595 ;
        RECT 105.105 88.425 105.275 88.595 ;
        RECT 105.565 88.425 105.735 88.595 ;
        RECT 106.025 88.425 106.195 88.595 ;
        RECT 106.485 88.425 106.655 88.595 ;
        RECT 106.945 88.425 107.115 88.595 ;
        RECT 107.405 88.425 107.575 88.595 ;
        RECT 107.865 88.425 108.035 88.595 ;
        RECT 108.325 88.425 108.495 88.595 ;
        RECT 108.785 88.425 108.955 88.595 ;
        RECT 109.245 88.425 109.415 88.595 ;
        RECT 109.705 88.425 109.875 88.595 ;
        RECT 110.165 88.425 110.335 88.595 ;
        RECT 110.625 88.425 110.795 88.595 ;
        RECT 111.085 88.425 111.255 88.595 ;
        RECT 111.545 88.425 111.715 88.595 ;
        RECT 112.005 88.425 112.175 88.595 ;
        RECT 112.465 88.425 112.635 88.595 ;
        RECT 112.925 88.425 113.095 88.595 ;
        RECT 113.385 88.425 113.555 88.595 ;
        RECT 113.845 88.425 114.015 88.595 ;
        RECT 114.305 88.425 114.475 88.595 ;
        RECT 114.765 88.425 114.935 88.595 ;
        RECT 115.225 88.425 115.395 88.595 ;
        RECT 115.685 88.425 115.855 88.595 ;
        RECT 116.145 88.425 116.315 88.595 ;
        RECT 116.605 88.425 116.775 88.595 ;
        RECT 117.065 88.425 117.235 88.595 ;
        RECT 117.525 88.425 117.695 88.595 ;
        RECT 117.985 88.425 118.155 88.595 ;
        RECT 118.445 88.425 118.615 88.595 ;
        RECT 118.905 88.425 119.075 88.595 ;
        RECT 119.365 88.425 119.535 88.595 ;
        RECT 119.825 88.425 119.995 88.595 ;
        RECT 120.285 88.425 120.455 88.595 ;
        RECT 120.745 88.425 120.915 88.595 ;
        RECT 121.205 88.425 121.375 88.595 ;
        RECT 121.665 88.425 121.835 88.595 ;
        RECT 122.125 88.425 122.295 88.595 ;
        RECT 122.585 88.425 122.755 88.595 ;
        RECT 123.045 88.425 123.215 88.595 ;
        RECT 123.505 88.425 123.675 88.595 ;
        RECT 123.965 88.425 124.135 88.595 ;
        RECT 124.425 88.425 124.595 88.595 ;
        RECT 124.885 88.425 125.055 88.595 ;
        RECT 125.345 88.425 125.515 88.595 ;
        RECT 125.805 88.425 125.975 88.595 ;
        RECT 126.265 88.425 126.435 88.595 ;
        RECT 126.725 88.425 126.895 88.595 ;
        RECT 127.185 88.425 127.355 88.595 ;
        RECT 127.645 88.425 127.815 88.595 ;
        RECT 128.105 88.425 128.275 88.595 ;
        RECT 128.565 88.425 128.735 88.595 ;
        RECT 129.025 88.425 129.195 88.595 ;
        RECT 129.485 88.425 129.655 88.595 ;
        RECT 129.945 88.425 130.115 88.595 ;
        RECT 130.405 88.425 130.575 88.595 ;
        RECT 130.865 88.425 131.035 88.595 ;
        RECT 131.325 88.425 131.495 88.595 ;
        RECT 131.785 88.425 131.955 88.595 ;
        RECT 132.245 88.425 132.415 88.595 ;
        RECT 132.705 88.425 132.875 88.595 ;
        RECT 133.165 88.425 133.335 88.595 ;
        RECT 133.625 88.425 133.795 88.595 ;
        RECT 134.085 88.425 134.255 88.595 ;
        RECT 134.545 88.425 134.715 88.595 ;
        RECT 135.005 88.425 135.175 88.595 ;
        RECT 135.465 88.425 135.635 88.595 ;
        RECT 135.925 88.425 136.095 88.595 ;
        RECT 136.385 88.425 136.555 88.595 ;
        RECT 136.845 88.425 137.015 88.595 ;
        RECT 137.305 88.425 137.475 88.595 ;
        RECT 137.765 88.425 137.935 88.595 ;
        RECT 138.225 88.425 138.395 88.595 ;
        RECT 138.685 88.425 138.855 88.595 ;
        RECT 139.145 88.425 139.315 88.595 ;
        RECT 139.605 88.425 139.775 88.595 ;
        RECT 140.065 88.425 140.235 88.595 ;
        RECT 140.525 88.425 140.695 88.595 ;
        RECT 140.985 88.425 141.155 88.595 ;
        RECT 141.445 88.425 141.615 88.595 ;
        RECT 141.905 88.425 142.075 88.595 ;
        RECT 142.365 88.425 142.535 88.595 ;
        RECT 142.825 88.425 142.995 88.595 ;
        RECT 143.285 88.425 143.455 88.595 ;
        RECT 143.745 88.425 143.915 88.595 ;
        RECT 144.205 88.425 144.375 88.595 ;
        RECT 144.665 88.425 144.835 88.595 ;
        RECT 145.125 88.425 145.295 88.595 ;
        RECT 145.585 88.425 145.755 88.595 ;
        RECT 146.045 88.425 146.215 88.595 ;
        RECT 146.505 88.425 146.675 88.595 ;
        RECT 146.965 88.425 147.135 88.595 ;
        RECT 147.425 88.425 147.595 88.595 ;
        RECT 147.885 88.425 148.055 88.595 ;
        RECT 148.345 88.425 148.515 88.595 ;
        RECT 148.805 88.425 148.975 88.595 ;
        RECT 149.265 88.425 149.435 88.595 ;
        RECT 149.725 88.425 149.895 88.595 ;
        RECT 150.185 88.425 150.355 88.595 ;
        RECT 11.265 85.705 11.435 85.875 ;
        RECT 11.725 85.705 11.895 85.875 ;
        RECT 12.185 85.705 12.355 85.875 ;
        RECT 12.645 85.705 12.815 85.875 ;
        RECT 13.105 85.705 13.275 85.875 ;
        RECT 13.565 85.705 13.735 85.875 ;
        RECT 14.025 85.705 14.195 85.875 ;
        RECT 14.485 85.705 14.655 85.875 ;
        RECT 14.945 85.705 15.115 85.875 ;
        RECT 15.405 85.705 15.575 85.875 ;
        RECT 15.865 85.705 16.035 85.875 ;
        RECT 16.325 85.705 16.495 85.875 ;
        RECT 16.785 85.705 16.955 85.875 ;
        RECT 17.245 85.705 17.415 85.875 ;
        RECT 17.705 85.705 17.875 85.875 ;
        RECT 18.165 85.705 18.335 85.875 ;
        RECT 18.625 85.705 18.795 85.875 ;
        RECT 19.085 85.705 19.255 85.875 ;
        RECT 19.545 85.705 19.715 85.875 ;
        RECT 20.005 85.705 20.175 85.875 ;
        RECT 20.465 85.705 20.635 85.875 ;
        RECT 20.925 85.705 21.095 85.875 ;
        RECT 21.385 85.705 21.555 85.875 ;
        RECT 21.845 85.705 22.015 85.875 ;
        RECT 22.305 85.705 22.475 85.875 ;
        RECT 22.765 85.705 22.935 85.875 ;
        RECT 23.225 85.705 23.395 85.875 ;
        RECT 23.685 85.705 23.855 85.875 ;
        RECT 24.145 85.705 24.315 85.875 ;
        RECT 24.605 85.705 24.775 85.875 ;
        RECT 25.065 85.705 25.235 85.875 ;
        RECT 25.525 85.705 25.695 85.875 ;
        RECT 25.985 85.705 26.155 85.875 ;
        RECT 26.445 85.705 26.615 85.875 ;
        RECT 26.905 85.705 27.075 85.875 ;
        RECT 27.365 85.705 27.535 85.875 ;
        RECT 27.825 85.705 27.995 85.875 ;
        RECT 28.285 85.705 28.455 85.875 ;
        RECT 28.745 85.705 28.915 85.875 ;
        RECT 29.205 85.705 29.375 85.875 ;
        RECT 29.665 85.705 29.835 85.875 ;
        RECT 30.125 85.705 30.295 85.875 ;
        RECT 30.585 85.705 30.755 85.875 ;
        RECT 31.045 85.705 31.215 85.875 ;
        RECT 31.505 85.705 31.675 85.875 ;
        RECT 31.965 85.705 32.135 85.875 ;
        RECT 32.425 85.705 32.595 85.875 ;
        RECT 32.885 85.705 33.055 85.875 ;
        RECT 33.345 85.705 33.515 85.875 ;
        RECT 33.805 85.705 33.975 85.875 ;
        RECT 34.265 85.705 34.435 85.875 ;
        RECT 34.725 85.705 34.895 85.875 ;
        RECT 35.185 85.705 35.355 85.875 ;
        RECT 35.645 85.705 35.815 85.875 ;
        RECT 36.105 85.705 36.275 85.875 ;
        RECT 36.565 85.705 36.735 85.875 ;
        RECT 37.025 85.705 37.195 85.875 ;
        RECT 37.485 85.705 37.655 85.875 ;
        RECT 37.945 85.705 38.115 85.875 ;
        RECT 38.405 85.705 38.575 85.875 ;
        RECT 38.865 85.705 39.035 85.875 ;
        RECT 39.325 85.705 39.495 85.875 ;
        RECT 39.785 85.705 39.955 85.875 ;
        RECT 40.245 85.705 40.415 85.875 ;
        RECT 40.705 85.705 40.875 85.875 ;
        RECT 41.165 85.705 41.335 85.875 ;
        RECT 41.625 85.705 41.795 85.875 ;
        RECT 42.085 85.705 42.255 85.875 ;
        RECT 42.545 85.705 42.715 85.875 ;
        RECT 43.005 85.705 43.175 85.875 ;
        RECT 43.465 85.705 43.635 85.875 ;
        RECT 43.925 85.705 44.095 85.875 ;
        RECT 44.385 85.705 44.555 85.875 ;
        RECT 44.845 85.705 45.015 85.875 ;
        RECT 45.305 85.705 45.475 85.875 ;
        RECT 45.765 85.705 45.935 85.875 ;
        RECT 46.225 85.705 46.395 85.875 ;
        RECT 46.685 85.705 46.855 85.875 ;
        RECT 47.145 85.705 47.315 85.875 ;
        RECT 47.605 85.705 47.775 85.875 ;
        RECT 48.065 85.705 48.235 85.875 ;
        RECT 48.525 85.705 48.695 85.875 ;
        RECT 48.985 85.705 49.155 85.875 ;
        RECT 49.445 85.705 49.615 85.875 ;
        RECT 49.905 85.705 50.075 85.875 ;
        RECT 50.365 85.705 50.535 85.875 ;
        RECT 50.825 85.705 50.995 85.875 ;
        RECT 51.285 85.705 51.455 85.875 ;
        RECT 51.745 85.705 51.915 85.875 ;
        RECT 52.205 85.705 52.375 85.875 ;
        RECT 52.665 85.705 52.835 85.875 ;
        RECT 53.125 85.705 53.295 85.875 ;
        RECT 53.585 85.705 53.755 85.875 ;
        RECT 54.045 85.705 54.215 85.875 ;
        RECT 54.505 85.705 54.675 85.875 ;
        RECT 54.965 85.705 55.135 85.875 ;
        RECT 55.425 85.705 55.595 85.875 ;
        RECT 55.885 85.705 56.055 85.875 ;
        RECT 56.345 85.705 56.515 85.875 ;
        RECT 56.805 85.705 56.975 85.875 ;
        RECT 57.265 85.705 57.435 85.875 ;
        RECT 57.725 85.705 57.895 85.875 ;
        RECT 58.185 85.705 58.355 85.875 ;
        RECT 58.645 85.705 58.815 85.875 ;
        RECT 59.105 85.705 59.275 85.875 ;
        RECT 59.565 85.705 59.735 85.875 ;
        RECT 60.025 85.705 60.195 85.875 ;
        RECT 60.485 85.705 60.655 85.875 ;
        RECT 60.945 85.705 61.115 85.875 ;
        RECT 61.405 85.705 61.575 85.875 ;
        RECT 61.865 85.705 62.035 85.875 ;
        RECT 62.325 85.705 62.495 85.875 ;
        RECT 62.785 85.705 62.955 85.875 ;
        RECT 63.245 85.705 63.415 85.875 ;
        RECT 63.705 85.705 63.875 85.875 ;
        RECT 64.165 85.705 64.335 85.875 ;
        RECT 64.625 85.705 64.795 85.875 ;
        RECT 65.085 85.705 65.255 85.875 ;
        RECT 65.545 85.705 65.715 85.875 ;
        RECT 66.005 85.705 66.175 85.875 ;
        RECT 66.465 85.705 66.635 85.875 ;
        RECT 66.925 85.705 67.095 85.875 ;
        RECT 67.385 85.705 67.555 85.875 ;
        RECT 67.845 85.705 68.015 85.875 ;
        RECT 68.305 85.705 68.475 85.875 ;
        RECT 68.765 85.705 68.935 85.875 ;
        RECT 69.225 85.705 69.395 85.875 ;
        RECT 69.685 85.705 69.855 85.875 ;
        RECT 70.145 85.705 70.315 85.875 ;
        RECT 70.605 85.705 70.775 85.875 ;
        RECT 71.065 85.705 71.235 85.875 ;
        RECT 71.525 85.705 71.695 85.875 ;
        RECT 71.985 85.705 72.155 85.875 ;
        RECT 72.445 85.705 72.615 85.875 ;
        RECT 72.905 85.705 73.075 85.875 ;
        RECT 73.365 85.705 73.535 85.875 ;
        RECT 73.825 85.705 73.995 85.875 ;
        RECT 74.285 85.705 74.455 85.875 ;
        RECT 74.745 85.705 74.915 85.875 ;
        RECT 75.205 85.705 75.375 85.875 ;
        RECT 75.665 85.705 75.835 85.875 ;
        RECT 76.125 85.705 76.295 85.875 ;
        RECT 76.585 85.705 76.755 85.875 ;
        RECT 77.045 85.705 77.215 85.875 ;
        RECT 77.505 85.705 77.675 85.875 ;
        RECT 77.965 85.705 78.135 85.875 ;
        RECT 78.425 85.705 78.595 85.875 ;
        RECT 78.885 85.705 79.055 85.875 ;
        RECT 79.345 85.705 79.515 85.875 ;
        RECT 79.805 85.705 79.975 85.875 ;
        RECT 80.265 85.705 80.435 85.875 ;
        RECT 80.725 85.705 80.895 85.875 ;
        RECT 81.185 85.705 81.355 85.875 ;
        RECT 81.645 85.705 81.815 85.875 ;
        RECT 82.105 85.705 82.275 85.875 ;
        RECT 82.565 85.705 82.735 85.875 ;
        RECT 83.025 85.705 83.195 85.875 ;
        RECT 83.485 85.705 83.655 85.875 ;
        RECT 83.945 85.705 84.115 85.875 ;
        RECT 84.405 85.705 84.575 85.875 ;
        RECT 84.865 85.705 85.035 85.875 ;
        RECT 85.325 85.705 85.495 85.875 ;
        RECT 85.785 85.705 85.955 85.875 ;
        RECT 86.245 85.705 86.415 85.875 ;
        RECT 86.705 85.705 86.875 85.875 ;
        RECT 87.165 85.705 87.335 85.875 ;
        RECT 87.625 85.705 87.795 85.875 ;
        RECT 88.085 85.705 88.255 85.875 ;
        RECT 88.545 85.705 88.715 85.875 ;
        RECT 89.005 85.705 89.175 85.875 ;
        RECT 89.465 85.705 89.635 85.875 ;
        RECT 89.925 85.705 90.095 85.875 ;
        RECT 90.385 85.705 90.555 85.875 ;
        RECT 90.845 85.705 91.015 85.875 ;
        RECT 91.305 85.705 91.475 85.875 ;
        RECT 91.765 85.705 91.935 85.875 ;
        RECT 92.225 85.705 92.395 85.875 ;
        RECT 92.685 85.705 92.855 85.875 ;
        RECT 93.145 85.705 93.315 85.875 ;
        RECT 93.605 85.705 93.775 85.875 ;
        RECT 94.065 85.705 94.235 85.875 ;
        RECT 94.525 85.705 94.695 85.875 ;
        RECT 94.985 85.705 95.155 85.875 ;
        RECT 95.445 85.705 95.615 85.875 ;
        RECT 95.905 85.705 96.075 85.875 ;
        RECT 96.365 85.705 96.535 85.875 ;
        RECT 96.825 85.705 96.995 85.875 ;
        RECT 97.285 85.705 97.455 85.875 ;
        RECT 97.745 85.705 97.915 85.875 ;
        RECT 98.205 85.705 98.375 85.875 ;
        RECT 98.665 85.705 98.835 85.875 ;
        RECT 99.125 85.705 99.295 85.875 ;
        RECT 99.585 85.705 99.755 85.875 ;
        RECT 100.045 85.705 100.215 85.875 ;
        RECT 100.505 85.705 100.675 85.875 ;
        RECT 100.965 85.705 101.135 85.875 ;
        RECT 101.425 85.705 101.595 85.875 ;
        RECT 101.885 85.705 102.055 85.875 ;
        RECT 102.345 85.705 102.515 85.875 ;
        RECT 102.805 85.705 102.975 85.875 ;
        RECT 103.265 85.705 103.435 85.875 ;
        RECT 103.725 85.705 103.895 85.875 ;
        RECT 104.185 85.705 104.355 85.875 ;
        RECT 104.645 85.705 104.815 85.875 ;
        RECT 105.105 85.705 105.275 85.875 ;
        RECT 105.565 85.705 105.735 85.875 ;
        RECT 106.025 85.705 106.195 85.875 ;
        RECT 106.485 85.705 106.655 85.875 ;
        RECT 106.945 85.705 107.115 85.875 ;
        RECT 107.405 85.705 107.575 85.875 ;
        RECT 107.865 85.705 108.035 85.875 ;
        RECT 108.325 85.705 108.495 85.875 ;
        RECT 108.785 85.705 108.955 85.875 ;
        RECT 109.245 85.705 109.415 85.875 ;
        RECT 109.705 85.705 109.875 85.875 ;
        RECT 110.165 85.705 110.335 85.875 ;
        RECT 110.625 85.705 110.795 85.875 ;
        RECT 111.085 85.705 111.255 85.875 ;
        RECT 111.545 85.705 111.715 85.875 ;
        RECT 112.005 85.705 112.175 85.875 ;
        RECT 112.465 85.705 112.635 85.875 ;
        RECT 112.925 85.705 113.095 85.875 ;
        RECT 113.385 85.705 113.555 85.875 ;
        RECT 113.845 85.705 114.015 85.875 ;
        RECT 114.305 85.705 114.475 85.875 ;
        RECT 114.765 85.705 114.935 85.875 ;
        RECT 115.225 85.705 115.395 85.875 ;
        RECT 115.685 85.705 115.855 85.875 ;
        RECT 116.145 85.705 116.315 85.875 ;
        RECT 116.605 85.705 116.775 85.875 ;
        RECT 117.065 85.705 117.235 85.875 ;
        RECT 117.525 85.705 117.695 85.875 ;
        RECT 117.985 85.705 118.155 85.875 ;
        RECT 118.445 85.705 118.615 85.875 ;
        RECT 118.905 85.705 119.075 85.875 ;
        RECT 119.365 85.705 119.535 85.875 ;
        RECT 119.825 85.705 119.995 85.875 ;
        RECT 120.285 85.705 120.455 85.875 ;
        RECT 120.745 85.705 120.915 85.875 ;
        RECT 121.205 85.705 121.375 85.875 ;
        RECT 121.665 85.705 121.835 85.875 ;
        RECT 122.125 85.705 122.295 85.875 ;
        RECT 122.585 85.705 122.755 85.875 ;
        RECT 123.045 85.705 123.215 85.875 ;
        RECT 123.505 85.705 123.675 85.875 ;
        RECT 123.965 85.705 124.135 85.875 ;
        RECT 124.425 85.705 124.595 85.875 ;
        RECT 124.885 85.705 125.055 85.875 ;
        RECT 125.345 85.705 125.515 85.875 ;
        RECT 125.805 85.705 125.975 85.875 ;
        RECT 126.265 85.705 126.435 85.875 ;
        RECT 126.725 85.705 126.895 85.875 ;
        RECT 127.185 85.705 127.355 85.875 ;
        RECT 127.645 85.705 127.815 85.875 ;
        RECT 128.105 85.705 128.275 85.875 ;
        RECT 128.565 85.705 128.735 85.875 ;
        RECT 129.025 85.705 129.195 85.875 ;
        RECT 129.485 85.705 129.655 85.875 ;
        RECT 129.945 85.705 130.115 85.875 ;
        RECT 130.405 85.705 130.575 85.875 ;
        RECT 130.865 85.705 131.035 85.875 ;
        RECT 131.325 85.705 131.495 85.875 ;
        RECT 131.785 85.705 131.955 85.875 ;
        RECT 132.245 85.705 132.415 85.875 ;
        RECT 132.705 85.705 132.875 85.875 ;
        RECT 133.165 85.705 133.335 85.875 ;
        RECT 133.625 85.705 133.795 85.875 ;
        RECT 134.085 85.705 134.255 85.875 ;
        RECT 134.545 85.705 134.715 85.875 ;
        RECT 135.005 85.705 135.175 85.875 ;
        RECT 135.465 85.705 135.635 85.875 ;
        RECT 135.925 85.705 136.095 85.875 ;
        RECT 136.385 85.705 136.555 85.875 ;
        RECT 136.845 85.705 137.015 85.875 ;
        RECT 137.305 85.705 137.475 85.875 ;
        RECT 137.765 85.705 137.935 85.875 ;
        RECT 138.225 85.705 138.395 85.875 ;
        RECT 138.685 85.705 138.855 85.875 ;
        RECT 139.145 85.705 139.315 85.875 ;
        RECT 139.605 85.705 139.775 85.875 ;
        RECT 140.065 85.705 140.235 85.875 ;
        RECT 140.525 85.705 140.695 85.875 ;
        RECT 140.985 85.705 141.155 85.875 ;
        RECT 141.445 85.705 141.615 85.875 ;
        RECT 141.905 85.705 142.075 85.875 ;
        RECT 142.365 85.705 142.535 85.875 ;
        RECT 142.825 85.705 142.995 85.875 ;
        RECT 143.285 85.705 143.455 85.875 ;
        RECT 143.745 85.705 143.915 85.875 ;
        RECT 144.205 85.705 144.375 85.875 ;
        RECT 144.665 85.705 144.835 85.875 ;
        RECT 145.125 85.705 145.295 85.875 ;
        RECT 145.585 85.705 145.755 85.875 ;
        RECT 146.045 85.705 146.215 85.875 ;
        RECT 146.505 85.705 146.675 85.875 ;
        RECT 146.965 85.705 147.135 85.875 ;
        RECT 147.425 85.705 147.595 85.875 ;
        RECT 147.885 85.705 148.055 85.875 ;
        RECT 148.345 85.705 148.515 85.875 ;
        RECT 148.805 85.705 148.975 85.875 ;
        RECT 149.265 85.705 149.435 85.875 ;
        RECT 149.725 85.705 149.895 85.875 ;
        RECT 150.185 85.705 150.355 85.875 ;
        RECT 11.265 82.985 11.435 83.155 ;
        RECT 11.725 82.985 11.895 83.155 ;
        RECT 12.185 82.985 12.355 83.155 ;
        RECT 12.645 82.985 12.815 83.155 ;
        RECT 13.105 82.985 13.275 83.155 ;
        RECT 13.565 82.985 13.735 83.155 ;
        RECT 14.025 82.985 14.195 83.155 ;
        RECT 14.485 82.985 14.655 83.155 ;
        RECT 14.945 82.985 15.115 83.155 ;
        RECT 15.405 82.985 15.575 83.155 ;
        RECT 15.865 82.985 16.035 83.155 ;
        RECT 16.325 82.985 16.495 83.155 ;
        RECT 16.785 82.985 16.955 83.155 ;
        RECT 17.245 82.985 17.415 83.155 ;
        RECT 17.705 82.985 17.875 83.155 ;
        RECT 18.165 82.985 18.335 83.155 ;
        RECT 18.625 82.985 18.795 83.155 ;
        RECT 19.085 82.985 19.255 83.155 ;
        RECT 19.545 82.985 19.715 83.155 ;
        RECT 20.005 82.985 20.175 83.155 ;
        RECT 20.465 82.985 20.635 83.155 ;
        RECT 20.925 82.985 21.095 83.155 ;
        RECT 21.385 82.985 21.555 83.155 ;
        RECT 21.845 82.985 22.015 83.155 ;
        RECT 22.305 82.985 22.475 83.155 ;
        RECT 22.765 82.985 22.935 83.155 ;
        RECT 23.225 82.985 23.395 83.155 ;
        RECT 23.685 82.985 23.855 83.155 ;
        RECT 24.145 82.985 24.315 83.155 ;
        RECT 24.605 82.985 24.775 83.155 ;
        RECT 25.065 82.985 25.235 83.155 ;
        RECT 25.525 82.985 25.695 83.155 ;
        RECT 25.985 82.985 26.155 83.155 ;
        RECT 26.445 82.985 26.615 83.155 ;
        RECT 26.905 82.985 27.075 83.155 ;
        RECT 27.365 82.985 27.535 83.155 ;
        RECT 27.825 82.985 27.995 83.155 ;
        RECT 28.285 82.985 28.455 83.155 ;
        RECT 28.745 82.985 28.915 83.155 ;
        RECT 29.205 82.985 29.375 83.155 ;
        RECT 29.665 82.985 29.835 83.155 ;
        RECT 30.125 82.985 30.295 83.155 ;
        RECT 30.585 82.985 30.755 83.155 ;
        RECT 31.045 82.985 31.215 83.155 ;
        RECT 31.505 82.985 31.675 83.155 ;
        RECT 31.965 82.985 32.135 83.155 ;
        RECT 32.425 82.985 32.595 83.155 ;
        RECT 32.885 82.985 33.055 83.155 ;
        RECT 33.345 82.985 33.515 83.155 ;
        RECT 33.805 82.985 33.975 83.155 ;
        RECT 34.265 82.985 34.435 83.155 ;
        RECT 34.725 82.985 34.895 83.155 ;
        RECT 35.185 82.985 35.355 83.155 ;
        RECT 35.645 82.985 35.815 83.155 ;
        RECT 36.105 82.985 36.275 83.155 ;
        RECT 36.565 82.985 36.735 83.155 ;
        RECT 37.025 82.985 37.195 83.155 ;
        RECT 37.485 82.985 37.655 83.155 ;
        RECT 37.945 82.985 38.115 83.155 ;
        RECT 38.405 82.985 38.575 83.155 ;
        RECT 38.865 82.985 39.035 83.155 ;
        RECT 39.325 82.985 39.495 83.155 ;
        RECT 39.785 82.985 39.955 83.155 ;
        RECT 40.245 82.985 40.415 83.155 ;
        RECT 40.705 82.985 40.875 83.155 ;
        RECT 41.165 82.985 41.335 83.155 ;
        RECT 41.625 82.985 41.795 83.155 ;
        RECT 42.085 82.985 42.255 83.155 ;
        RECT 42.545 82.985 42.715 83.155 ;
        RECT 43.005 82.985 43.175 83.155 ;
        RECT 43.465 82.985 43.635 83.155 ;
        RECT 43.925 82.985 44.095 83.155 ;
        RECT 44.385 82.985 44.555 83.155 ;
        RECT 44.845 82.985 45.015 83.155 ;
        RECT 45.305 82.985 45.475 83.155 ;
        RECT 45.765 82.985 45.935 83.155 ;
        RECT 46.225 82.985 46.395 83.155 ;
        RECT 46.685 82.985 46.855 83.155 ;
        RECT 47.145 82.985 47.315 83.155 ;
        RECT 47.605 82.985 47.775 83.155 ;
        RECT 48.065 82.985 48.235 83.155 ;
        RECT 48.525 82.985 48.695 83.155 ;
        RECT 48.985 82.985 49.155 83.155 ;
        RECT 49.445 82.985 49.615 83.155 ;
        RECT 49.905 82.985 50.075 83.155 ;
        RECT 50.365 82.985 50.535 83.155 ;
        RECT 50.825 82.985 50.995 83.155 ;
        RECT 51.285 82.985 51.455 83.155 ;
        RECT 51.745 82.985 51.915 83.155 ;
        RECT 52.205 82.985 52.375 83.155 ;
        RECT 52.665 82.985 52.835 83.155 ;
        RECT 53.125 82.985 53.295 83.155 ;
        RECT 53.585 82.985 53.755 83.155 ;
        RECT 54.045 82.985 54.215 83.155 ;
        RECT 54.505 82.985 54.675 83.155 ;
        RECT 54.965 82.985 55.135 83.155 ;
        RECT 55.425 82.985 55.595 83.155 ;
        RECT 55.885 82.985 56.055 83.155 ;
        RECT 56.345 82.985 56.515 83.155 ;
        RECT 56.805 82.985 56.975 83.155 ;
        RECT 57.265 82.985 57.435 83.155 ;
        RECT 57.725 82.985 57.895 83.155 ;
        RECT 58.185 82.985 58.355 83.155 ;
        RECT 58.645 82.985 58.815 83.155 ;
        RECT 59.105 82.985 59.275 83.155 ;
        RECT 59.565 82.985 59.735 83.155 ;
        RECT 60.025 82.985 60.195 83.155 ;
        RECT 60.485 82.985 60.655 83.155 ;
        RECT 60.945 82.985 61.115 83.155 ;
        RECT 61.405 82.985 61.575 83.155 ;
        RECT 61.865 82.985 62.035 83.155 ;
        RECT 62.325 82.985 62.495 83.155 ;
        RECT 62.785 82.985 62.955 83.155 ;
        RECT 63.245 82.985 63.415 83.155 ;
        RECT 63.705 82.985 63.875 83.155 ;
        RECT 64.165 82.985 64.335 83.155 ;
        RECT 64.625 82.985 64.795 83.155 ;
        RECT 65.085 82.985 65.255 83.155 ;
        RECT 65.545 82.985 65.715 83.155 ;
        RECT 66.005 82.985 66.175 83.155 ;
        RECT 66.465 82.985 66.635 83.155 ;
        RECT 66.925 82.985 67.095 83.155 ;
        RECT 67.385 82.985 67.555 83.155 ;
        RECT 67.845 82.985 68.015 83.155 ;
        RECT 68.305 82.985 68.475 83.155 ;
        RECT 68.765 82.985 68.935 83.155 ;
        RECT 69.225 82.985 69.395 83.155 ;
        RECT 69.685 82.985 69.855 83.155 ;
        RECT 70.145 82.985 70.315 83.155 ;
        RECT 70.605 82.985 70.775 83.155 ;
        RECT 71.065 82.985 71.235 83.155 ;
        RECT 71.525 82.985 71.695 83.155 ;
        RECT 71.985 82.985 72.155 83.155 ;
        RECT 72.445 82.985 72.615 83.155 ;
        RECT 72.905 82.985 73.075 83.155 ;
        RECT 73.365 82.985 73.535 83.155 ;
        RECT 73.825 82.985 73.995 83.155 ;
        RECT 74.285 82.985 74.455 83.155 ;
        RECT 74.745 82.985 74.915 83.155 ;
        RECT 75.205 82.985 75.375 83.155 ;
        RECT 75.665 82.985 75.835 83.155 ;
        RECT 76.125 82.985 76.295 83.155 ;
        RECT 76.585 82.985 76.755 83.155 ;
        RECT 77.045 82.985 77.215 83.155 ;
        RECT 77.505 82.985 77.675 83.155 ;
        RECT 77.965 82.985 78.135 83.155 ;
        RECT 78.425 82.985 78.595 83.155 ;
        RECT 78.885 82.985 79.055 83.155 ;
        RECT 79.345 82.985 79.515 83.155 ;
        RECT 79.805 82.985 79.975 83.155 ;
        RECT 80.265 82.985 80.435 83.155 ;
        RECT 80.725 82.985 80.895 83.155 ;
        RECT 81.185 82.985 81.355 83.155 ;
        RECT 81.645 82.985 81.815 83.155 ;
        RECT 82.105 82.985 82.275 83.155 ;
        RECT 82.565 82.985 82.735 83.155 ;
        RECT 83.025 82.985 83.195 83.155 ;
        RECT 83.485 82.985 83.655 83.155 ;
        RECT 83.945 82.985 84.115 83.155 ;
        RECT 84.405 82.985 84.575 83.155 ;
        RECT 84.865 82.985 85.035 83.155 ;
        RECT 85.325 82.985 85.495 83.155 ;
        RECT 85.785 82.985 85.955 83.155 ;
        RECT 86.245 82.985 86.415 83.155 ;
        RECT 86.705 82.985 86.875 83.155 ;
        RECT 87.165 82.985 87.335 83.155 ;
        RECT 87.625 82.985 87.795 83.155 ;
        RECT 88.085 82.985 88.255 83.155 ;
        RECT 88.545 82.985 88.715 83.155 ;
        RECT 89.005 82.985 89.175 83.155 ;
        RECT 89.465 82.985 89.635 83.155 ;
        RECT 89.925 82.985 90.095 83.155 ;
        RECT 90.385 82.985 90.555 83.155 ;
        RECT 90.845 82.985 91.015 83.155 ;
        RECT 91.305 82.985 91.475 83.155 ;
        RECT 91.765 82.985 91.935 83.155 ;
        RECT 92.225 82.985 92.395 83.155 ;
        RECT 92.685 82.985 92.855 83.155 ;
        RECT 93.145 82.985 93.315 83.155 ;
        RECT 93.605 82.985 93.775 83.155 ;
        RECT 94.065 82.985 94.235 83.155 ;
        RECT 94.525 82.985 94.695 83.155 ;
        RECT 94.985 82.985 95.155 83.155 ;
        RECT 95.445 82.985 95.615 83.155 ;
        RECT 95.905 82.985 96.075 83.155 ;
        RECT 96.365 82.985 96.535 83.155 ;
        RECT 96.825 82.985 96.995 83.155 ;
        RECT 97.285 82.985 97.455 83.155 ;
        RECT 97.745 82.985 97.915 83.155 ;
        RECT 98.205 82.985 98.375 83.155 ;
        RECT 98.665 82.985 98.835 83.155 ;
        RECT 99.125 82.985 99.295 83.155 ;
        RECT 99.585 82.985 99.755 83.155 ;
        RECT 100.045 82.985 100.215 83.155 ;
        RECT 100.505 82.985 100.675 83.155 ;
        RECT 100.965 82.985 101.135 83.155 ;
        RECT 101.425 82.985 101.595 83.155 ;
        RECT 101.885 82.985 102.055 83.155 ;
        RECT 102.345 82.985 102.515 83.155 ;
        RECT 102.805 82.985 102.975 83.155 ;
        RECT 103.265 82.985 103.435 83.155 ;
        RECT 103.725 82.985 103.895 83.155 ;
        RECT 104.185 82.985 104.355 83.155 ;
        RECT 104.645 82.985 104.815 83.155 ;
        RECT 105.105 82.985 105.275 83.155 ;
        RECT 105.565 82.985 105.735 83.155 ;
        RECT 106.025 82.985 106.195 83.155 ;
        RECT 106.485 82.985 106.655 83.155 ;
        RECT 106.945 82.985 107.115 83.155 ;
        RECT 107.405 82.985 107.575 83.155 ;
        RECT 107.865 82.985 108.035 83.155 ;
        RECT 108.325 82.985 108.495 83.155 ;
        RECT 108.785 82.985 108.955 83.155 ;
        RECT 109.245 82.985 109.415 83.155 ;
        RECT 109.705 82.985 109.875 83.155 ;
        RECT 110.165 82.985 110.335 83.155 ;
        RECT 110.625 82.985 110.795 83.155 ;
        RECT 111.085 82.985 111.255 83.155 ;
        RECT 111.545 82.985 111.715 83.155 ;
        RECT 112.005 82.985 112.175 83.155 ;
        RECT 112.465 82.985 112.635 83.155 ;
        RECT 112.925 82.985 113.095 83.155 ;
        RECT 113.385 82.985 113.555 83.155 ;
        RECT 113.845 82.985 114.015 83.155 ;
        RECT 114.305 82.985 114.475 83.155 ;
        RECT 114.765 82.985 114.935 83.155 ;
        RECT 115.225 82.985 115.395 83.155 ;
        RECT 115.685 82.985 115.855 83.155 ;
        RECT 116.145 82.985 116.315 83.155 ;
        RECT 116.605 82.985 116.775 83.155 ;
        RECT 117.065 82.985 117.235 83.155 ;
        RECT 117.525 82.985 117.695 83.155 ;
        RECT 117.985 82.985 118.155 83.155 ;
        RECT 118.445 82.985 118.615 83.155 ;
        RECT 118.905 82.985 119.075 83.155 ;
        RECT 119.365 82.985 119.535 83.155 ;
        RECT 119.825 82.985 119.995 83.155 ;
        RECT 120.285 82.985 120.455 83.155 ;
        RECT 120.745 82.985 120.915 83.155 ;
        RECT 121.205 82.985 121.375 83.155 ;
        RECT 121.665 82.985 121.835 83.155 ;
        RECT 122.125 82.985 122.295 83.155 ;
        RECT 122.585 82.985 122.755 83.155 ;
        RECT 123.045 82.985 123.215 83.155 ;
        RECT 123.505 82.985 123.675 83.155 ;
        RECT 123.965 82.985 124.135 83.155 ;
        RECT 124.425 82.985 124.595 83.155 ;
        RECT 124.885 82.985 125.055 83.155 ;
        RECT 125.345 82.985 125.515 83.155 ;
        RECT 125.805 82.985 125.975 83.155 ;
        RECT 126.265 82.985 126.435 83.155 ;
        RECT 126.725 82.985 126.895 83.155 ;
        RECT 127.185 82.985 127.355 83.155 ;
        RECT 127.645 82.985 127.815 83.155 ;
        RECT 128.105 82.985 128.275 83.155 ;
        RECT 128.565 82.985 128.735 83.155 ;
        RECT 129.025 82.985 129.195 83.155 ;
        RECT 129.485 82.985 129.655 83.155 ;
        RECT 129.945 82.985 130.115 83.155 ;
        RECT 130.405 82.985 130.575 83.155 ;
        RECT 130.865 82.985 131.035 83.155 ;
        RECT 131.325 82.985 131.495 83.155 ;
        RECT 131.785 82.985 131.955 83.155 ;
        RECT 132.245 82.985 132.415 83.155 ;
        RECT 132.705 82.985 132.875 83.155 ;
        RECT 133.165 82.985 133.335 83.155 ;
        RECT 133.625 82.985 133.795 83.155 ;
        RECT 134.085 82.985 134.255 83.155 ;
        RECT 134.545 82.985 134.715 83.155 ;
        RECT 135.005 82.985 135.175 83.155 ;
        RECT 135.465 82.985 135.635 83.155 ;
        RECT 135.925 82.985 136.095 83.155 ;
        RECT 136.385 82.985 136.555 83.155 ;
        RECT 136.845 82.985 137.015 83.155 ;
        RECT 137.305 82.985 137.475 83.155 ;
        RECT 137.765 82.985 137.935 83.155 ;
        RECT 138.225 82.985 138.395 83.155 ;
        RECT 138.685 82.985 138.855 83.155 ;
        RECT 139.145 82.985 139.315 83.155 ;
        RECT 139.605 82.985 139.775 83.155 ;
        RECT 140.065 82.985 140.235 83.155 ;
        RECT 140.525 82.985 140.695 83.155 ;
        RECT 140.985 82.985 141.155 83.155 ;
        RECT 141.445 82.985 141.615 83.155 ;
        RECT 141.905 82.985 142.075 83.155 ;
        RECT 142.365 82.985 142.535 83.155 ;
        RECT 142.825 82.985 142.995 83.155 ;
        RECT 143.285 82.985 143.455 83.155 ;
        RECT 143.745 82.985 143.915 83.155 ;
        RECT 144.205 82.985 144.375 83.155 ;
        RECT 144.665 82.985 144.835 83.155 ;
        RECT 145.125 82.985 145.295 83.155 ;
        RECT 145.585 82.985 145.755 83.155 ;
        RECT 146.045 82.985 146.215 83.155 ;
        RECT 146.505 82.985 146.675 83.155 ;
        RECT 146.965 82.985 147.135 83.155 ;
        RECT 147.425 82.985 147.595 83.155 ;
        RECT 147.885 82.985 148.055 83.155 ;
        RECT 148.345 82.985 148.515 83.155 ;
        RECT 148.805 82.985 148.975 83.155 ;
        RECT 149.265 82.985 149.435 83.155 ;
        RECT 149.725 82.985 149.895 83.155 ;
        RECT 150.185 82.985 150.355 83.155 ;
        RECT 11.265 80.265 11.435 80.435 ;
        RECT 11.725 80.265 11.895 80.435 ;
        RECT 12.185 80.265 12.355 80.435 ;
        RECT 12.645 80.265 12.815 80.435 ;
        RECT 13.105 80.265 13.275 80.435 ;
        RECT 13.565 80.265 13.735 80.435 ;
        RECT 14.025 80.265 14.195 80.435 ;
        RECT 14.485 80.265 14.655 80.435 ;
        RECT 14.945 80.265 15.115 80.435 ;
        RECT 15.405 80.265 15.575 80.435 ;
        RECT 15.865 80.265 16.035 80.435 ;
        RECT 16.325 80.265 16.495 80.435 ;
        RECT 16.785 80.265 16.955 80.435 ;
        RECT 17.245 80.265 17.415 80.435 ;
        RECT 17.705 80.265 17.875 80.435 ;
        RECT 18.165 80.265 18.335 80.435 ;
        RECT 18.625 80.265 18.795 80.435 ;
        RECT 19.085 80.265 19.255 80.435 ;
        RECT 19.545 80.265 19.715 80.435 ;
        RECT 20.005 80.265 20.175 80.435 ;
        RECT 20.465 80.265 20.635 80.435 ;
        RECT 20.925 80.265 21.095 80.435 ;
        RECT 21.385 80.265 21.555 80.435 ;
        RECT 21.845 80.265 22.015 80.435 ;
        RECT 22.305 80.265 22.475 80.435 ;
        RECT 22.765 80.265 22.935 80.435 ;
        RECT 23.225 80.265 23.395 80.435 ;
        RECT 23.685 80.265 23.855 80.435 ;
        RECT 24.145 80.265 24.315 80.435 ;
        RECT 24.605 80.265 24.775 80.435 ;
        RECT 25.065 80.265 25.235 80.435 ;
        RECT 25.525 80.265 25.695 80.435 ;
        RECT 25.985 80.265 26.155 80.435 ;
        RECT 26.445 80.265 26.615 80.435 ;
        RECT 26.905 80.265 27.075 80.435 ;
        RECT 27.365 80.265 27.535 80.435 ;
        RECT 27.825 80.265 27.995 80.435 ;
        RECT 28.285 80.265 28.455 80.435 ;
        RECT 28.745 80.265 28.915 80.435 ;
        RECT 29.205 80.265 29.375 80.435 ;
        RECT 29.665 80.265 29.835 80.435 ;
        RECT 30.125 80.265 30.295 80.435 ;
        RECT 30.585 80.265 30.755 80.435 ;
        RECT 31.045 80.265 31.215 80.435 ;
        RECT 31.505 80.265 31.675 80.435 ;
        RECT 31.965 80.265 32.135 80.435 ;
        RECT 32.425 80.265 32.595 80.435 ;
        RECT 32.885 80.265 33.055 80.435 ;
        RECT 33.345 80.265 33.515 80.435 ;
        RECT 33.805 80.265 33.975 80.435 ;
        RECT 34.265 80.265 34.435 80.435 ;
        RECT 34.725 80.265 34.895 80.435 ;
        RECT 35.185 80.265 35.355 80.435 ;
        RECT 35.645 80.265 35.815 80.435 ;
        RECT 36.105 80.265 36.275 80.435 ;
        RECT 36.565 80.265 36.735 80.435 ;
        RECT 37.025 80.265 37.195 80.435 ;
        RECT 37.485 80.265 37.655 80.435 ;
        RECT 37.945 80.265 38.115 80.435 ;
        RECT 38.405 80.265 38.575 80.435 ;
        RECT 38.865 80.265 39.035 80.435 ;
        RECT 39.325 80.265 39.495 80.435 ;
        RECT 39.785 80.265 39.955 80.435 ;
        RECT 40.245 80.265 40.415 80.435 ;
        RECT 40.705 80.265 40.875 80.435 ;
        RECT 41.165 80.265 41.335 80.435 ;
        RECT 41.625 80.265 41.795 80.435 ;
        RECT 42.085 80.265 42.255 80.435 ;
        RECT 42.545 80.265 42.715 80.435 ;
        RECT 43.005 80.265 43.175 80.435 ;
        RECT 43.465 80.265 43.635 80.435 ;
        RECT 43.925 80.265 44.095 80.435 ;
        RECT 44.385 80.265 44.555 80.435 ;
        RECT 44.845 80.265 45.015 80.435 ;
        RECT 45.305 80.265 45.475 80.435 ;
        RECT 45.765 80.265 45.935 80.435 ;
        RECT 46.225 80.265 46.395 80.435 ;
        RECT 46.685 80.265 46.855 80.435 ;
        RECT 47.145 80.265 47.315 80.435 ;
        RECT 47.605 80.265 47.775 80.435 ;
        RECT 48.065 80.265 48.235 80.435 ;
        RECT 48.525 80.265 48.695 80.435 ;
        RECT 48.985 80.265 49.155 80.435 ;
        RECT 49.445 80.265 49.615 80.435 ;
        RECT 49.905 80.265 50.075 80.435 ;
        RECT 50.365 80.265 50.535 80.435 ;
        RECT 50.825 80.265 50.995 80.435 ;
        RECT 51.285 80.265 51.455 80.435 ;
        RECT 51.745 80.265 51.915 80.435 ;
        RECT 52.205 80.265 52.375 80.435 ;
        RECT 52.665 80.265 52.835 80.435 ;
        RECT 53.125 80.265 53.295 80.435 ;
        RECT 53.585 80.265 53.755 80.435 ;
        RECT 54.045 80.265 54.215 80.435 ;
        RECT 54.505 80.265 54.675 80.435 ;
        RECT 54.965 80.265 55.135 80.435 ;
        RECT 55.425 80.265 55.595 80.435 ;
        RECT 55.885 80.265 56.055 80.435 ;
        RECT 56.345 80.265 56.515 80.435 ;
        RECT 56.805 80.265 56.975 80.435 ;
        RECT 57.265 80.265 57.435 80.435 ;
        RECT 57.725 80.265 57.895 80.435 ;
        RECT 58.185 80.265 58.355 80.435 ;
        RECT 58.645 80.265 58.815 80.435 ;
        RECT 59.105 80.265 59.275 80.435 ;
        RECT 59.565 80.265 59.735 80.435 ;
        RECT 60.025 80.265 60.195 80.435 ;
        RECT 60.485 80.265 60.655 80.435 ;
        RECT 60.945 80.265 61.115 80.435 ;
        RECT 61.405 80.265 61.575 80.435 ;
        RECT 61.865 80.265 62.035 80.435 ;
        RECT 62.325 80.265 62.495 80.435 ;
        RECT 62.785 80.265 62.955 80.435 ;
        RECT 63.245 80.265 63.415 80.435 ;
        RECT 63.705 80.265 63.875 80.435 ;
        RECT 64.165 80.265 64.335 80.435 ;
        RECT 64.625 80.265 64.795 80.435 ;
        RECT 65.085 80.265 65.255 80.435 ;
        RECT 65.545 80.265 65.715 80.435 ;
        RECT 66.005 80.265 66.175 80.435 ;
        RECT 66.465 80.265 66.635 80.435 ;
        RECT 66.925 80.265 67.095 80.435 ;
        RECT 67.385 80.265 67.555 80.435 ;
        RECT 67.845 80.265 68.015 80.435 ;
        RECT 68.305 80.265 68.475 80.435 ;
        RECT 68.765 80.265 68.935 80.435 ;
        RECT 69.225 80.265 69.395 80.435 ;
        RECT 69.685 80.265 69.855 80.435 ;
        RECT 70.145 80.265 70.315 80.435 ;
        RECT 70.605 80.265 70.775 80.435 ;
        RECT 71.065 80.265 71.235 80.435 ;
        RECT 71.525 80.265 71.695 80.435 ;
        RECT 71.985 80.265 72.155 80.435 ;
        RECT 72.445 80.265 72.615 80.435 ;
        RECT 72.905 80.265 73.075 80.435 ;
        RECT 73.365 80.265 73.535 80.435 ;
        RECT 73.825 80.265 73.995 80.435 ;
        RECT 74.285 80.265 74.455 80.435 ;
        RECT 74.745 80.265 74.915 80.435 ;
        RECT 75.205 80.265 75.375 80.435 ;
        RECT 75.665 80.265 75.835 80.435 ;
        RECT 76.125 80.265 76.295 80.435 ;
        RECT 76.585 80.265 76.755 80.435 ;
        RECT 77.045 80.265 77.215 80.435 ;
        RECT 77.505 80.265 77.675 80.435 ;
        RECT 77.965 80.265 78.135 80.435 ;
        RECT 78.425 80.265 78.595 80.435 ;
        RECT 78.885 80.265 79.055 80.435 ;
        RECT 79.345 80.265 79.515 80.435 ;
        RECT 79.805 80.265 79.975 80.435 ;
        RECT 80.265 80.265 80.435 80.435 ;
        RECT 80.725 80.265 80.895 80.435 ;
        RECT 81.185 80.265 81.355 80.435 ;
        RECT 81.645 80.265 81.815 80.435 ;
        RECT 82.105 80.265 82.275 80.435 ;
        RECT 82.565 80.265 82.735 80.435 ;
        RECT 83.025 80.265 83.195 80.435 ;
        RECT 83.485 80.265 83.655 80.435 ;
        RECT 83.945 80.265 84.115 80.435 ;
        RECT 84.405 80.265 84.575 80.435 ;
        RECT 84.865 80.265 85.035 80.435 ;
        RECT 85.325 80.265 85.495 80.435 ;
        RECT 85.785 80.265 85.955 80.435 ;
        RECT 86.245 80.265 86.415 80.435 ;
        RECT 86.705 80.265 86.875 80.435 ;
        RECT 87.165 80.265 87.335 80.435 ;
        RECT 87.625 80.265 87.795 80.435 ;
        RECT 88.085 80.265 88.255 80.435 ;
        RECT 88.545 80.265 88.715 80.435 ;
        RECT 89.005 80.265 89.175 80.435 ;
        RECT 89.465 80.265 89.635 80.435 ;
        RECT 89.925 80.265 90.095 80.435 ;
        RECT 90.385 80.265 90.555 80.435 ;
        RECT 90.845 80.265 91.015 80.435 ;
        RECT 91.305 80.265 91.475 80.435 ;
        RECT 91.765 80.265 91.935 80.435 ;
        RECT 92.225 80.265 92.395 80.435 ;
        RECT 92.685 80.265 92.855 80.435 ;
        RECT 93.145 80.265 93.315 80.435 ;
        RECT 93.605 80.265 93.775 80.435 ;
        RECT 94.065 80.265 94.235 80.435 ;
        RECT 94.525 80.265 94.695 80.435 ;
        RECT 94.985 80.265 95.155 80.435 ;
        RECT 95.445 80.265 95.615 80.435 ;
        RECT 95.905 80.265 96.075 80.435 ;
        RECT 96.365 80.265 96.535 80.435 ;
        RECT 96.825 80.265 96.995 80.435 ;
        RECT 97.285 80.265 97.455 80.435 ;
        RECT 97.745 80.265 97.915 80.435 ;
        RECT 98.205 80.265 98.375 80.435 ;
        RECT 98.665 80.265 98.835 80.435 ;
        RECT 99.125 80.265 99.295 80.435 ;
        RECT 99.585 80.265 99.755 80.435 ;
        RECT 100.045 80.265 100.215 80.435 ;
        RECT 100.505 80.265 100.675 80.435 ;
        RECT 100.965 80.265 101.135 80.435 ;
        RECT 101.425 80.265 101.595 80.435 ;
        RECT 101.885 80.265 102.055 80.435 ;
        RECT 102.345 80.265 102.515 80.435 ;
        RECT 102.805 80.265 102.975 80.435 ;
        RECT 103.265 80.265 103.435 80.435 ;
        RECT 103.725 80.265 103.895 80.435 ;
        RECT 104.185 80.265 104.355 80.435 ;
        RECT 104.645 80.265 104.815 80.435 ;
        RECT 105.105 80.265 105.275 80.435 ;
        RECT 105.565 80.265 105.735 80.435 ;
        RECT 106.025 80.265 106.195 80.435 ;
        RECT 106.485 80.265 106.655 80.435 ;
        RECT 106.945 80.265 107.115 80.435 ;
        RECT 107.405 80.265 107.575 80.435 ;
        RECT 107.865 80.265 108.035 80.435 ;
        RECT 108.325 80.265 108.495 80.435 ;
        RECT 108.785 80.265 108.955 80.435 ;
        RECT 109.245 80.265 109.415 80.435 ;
        RECT 109.705 80.265 109.875 80.435 ;
        RECT 110.165 80.265 110.335 80.435 ;
        RECT 110.625 80.265 110.795 80.435 ;
        RECT 111.085 80.265 111.255 80.435 ;
        RECT 111.545 80.265 111.715 80.435 ;
        RECT 112.005 80.265 112.175 80.435 ;
        RECT 112.465 80.265 112.635 80.435 ;
        RECT 112.925 80.265 113.095 80.435 ;
        RECT 113.385 80.265 113.555 80.435 ;
        RECT 113.845 80.265 114.015 80.435 ;
        RECT 114.305 80.265 114.475 80.435 ;
        RECT 114.765 80.265 114.935 80.435 ;
        RECT 115.225 80.265 115.395 80.435 ;
        RECT 115.685 80.265 115.855 80.435 ;
        RECT 116.145 80.265 116.315 80.435 ;
        RECT 116.605 80.265 116.775 80.435 ;
        RECT 117.065 80.265 117.235 80.435 ;
        RECT 117.525 80.265 117.695 80.435 ;
        RECT 117.985 80.265 118.155 80.435 ;
        RECT 118.445 80.265 118.615 80.435 ;
        RECT 118.905 80.265 119.075 80.435 ;
        RECT 119.365 80.265 119.535 80.435 ;
        RECT 119.825 80.265 119.995 80.435 ;
        RECT 120.285 80.265 120.455 80.435 ;
        RECT 120.745 80.265 120.915 80.435 ;
        RECT 121.205 80.265 121.375 80.435 ;
        RECT 121.665 80.265 121.835 80.435 ;
        RECT 122.125 80.265 122.295 80.435 ;
        RECT 122.585 80.265 122.755 80.435 ;
        RECT 123.045 80.265 123.215 80.435 ;
        RECT 123.505 80.265 123.675 80.435 ;
        RECT 123.965 80.265 124.135 80.435 ;
        RECT 124.425 80.265 124.595 80.435 ;
        RECT 124.885 80.265 125.055 80.435 ;
        RECT 125.345 80.265 125.515 80.435 ;
        RECT 125.805 80.265 125.975 80.435 ;
        RECT 126.265 80.265 126.435 80.435 ;
        RECT 126.725 80.265 126.895 80.435 ;
        RECT 127.185 80.265 127.355 80.435 ;
        RECT 127.645 80.265 127.815 80.435 ;
        RECT 128.105 80.265 128.275 80.435 ;
        RECT 128.565 80.265 128.735 80.435 ;
        RECT 129.025 80.265 129.195 80.435 ;
        RECT 129.485 80.265 129.655 80.435 ;
        RECT 129.945 80.265 130.115 80.435 ;
        RECT 130.405 80.265 130.575 80.435 ;
        RECT 130.865 80.265 131.035 80.435 ;
        RECT 131.325 80.265 131.495 80.435 ;
        RECT 131.785 80.265 131.955 80.435 ;
        RECT 132.245 80.265 132.415 80.435 ;
        RECT 132.705 80.265 132.875 80.435 ;
        RECT 133.165 80.265 133.335 80.435 ;
        RECT 133.625 80.265 133.795 80.435 ;
        RECT 134.085 80.265 134.255 80.435 ;
        RECT 134.545 80.265 134.715 80.435 ;
        RECT 135.005 80.265 135.175 80.435 ;
        RECT 135.465 80.265 135.635 80.435 ;
        RECT 135.925 80.265 136.095 80.435 ;
        RECT 136.385 80.265 136.555 80.435 ;
        RECT 136.845 80.265 137.015 80.435 ;
        RECT 137.305 80.265 137.475 80.435 ;
        RECT 137.765 80.265 137.935 80.435 ;
        RECT 138.225 80.265 138.395 80.435 ;
        RECT 138.685 80.265 138.855 80.435 ;
        RECT 139.145 80.265 139.315 80.435 ;
        RECT 139.605 80.265 139.775 80.435 ;
        RECT 140.065 80.265 140.235 80.435 ;
        RECT 140.525 80.265 140.695 80.435 ;
        RECT 140.985 80.265 141.155 80.435 ;
        RECT 141.445 80.265 141.615 80.435 ;
        RECT 141.905 80.265 142.075 80.435 ;
        RECT 142.365 80.265 142.535 80.435 ;
        RECT 142.825 80.265 142.995 80.435 ;
        RECT 143.285 80.265 143.455 80.435 ;
        RECT 143.745 80.265 143.915 80.435 ;
        RECT 144.205 80.265 144.375 80.435 ;
        RECT 144.665 80.265 144.835 80.435 ;
        RECT 145.125 80.265 145.295 80.435 ;
        RECT 145.585 80.265 145.755 80.435 ;
        RECT 146.045 80.265 146.215 80.435 ;
        RECT 146.505 80.265 146.675 80.435 ;
        RECT 146.965 80.265 147.135 80.435 ;
        RECT 147.425 80.265 147.595 80.435 ;
        RECT 147.885 80.265 148.055 80.435 ;
        RECT 148.345 80.265 148.515 80.435 ;
        RECT 148.805 80.265 148.975 80.435 ;
        RECT 149.265 80.265 149.435 80.435 ;
        RECT 149.725 80.265 149.895 80.435 ;
        RECT 150.185 80.265 150.355 80.435 ;
        RECT 11.265 77.545 11.435 77.715 ;
        RECT 11.725 77.545 11.895 77.715 ;
        RECT 12.185 77.545 12.355 77.715 ;
        RECT 12.645 77.545 12.815 77.715 ;
        RECT 13.105 77.545 13.275 77.715 ;
        RECT 13.565 77.545 13.735 77.715 ;
        RECT 14.025 77.545 14.195 77.715 ;
        RECT 14.485 77.545 14.655 77.715 ;
        RECT 14.945 77.545 15.115 77.715 ;
        RECT 15.405 77.545 15.575 77.715 ;
        RECT 15.865 77.545 16.035 77.715 ;
        RECT 16.325 77.545 16.495 77.715 ;
        RECT 16.785 77.545 16.955 77.715 ;
        RECT 17.245 77.545 17.415 77.715 ;
        RECT 17.705 77.545 17.875 77.715 ;
        RECT 18.165 77.545 18.335 77.715 ;
        RECT 18.625 77.545 18.795 77.715 ;
        RECT 19.085 77.545 19.255 77.715 ;
        RECT 19.545 77.545 19.715 77.715 ;
        RECT 20.005 77.545 20.175 77.715 ;
        RECT 20.465 77.545 20.635 77.715 ;
        RECT 20.925 77.545 21.095 77.715 ;
        RECT 21.385 77.545 21.555 77.715 ;
        RECT 21.845 77.545 22.015 77.715 ;
        RECT 22.305 77.545 22.475 77.715 ;
        RECT 22.765 77.545 22.935 77.715 ;
        RECT 23.225 77.545 23.395 77.715 ;
        RECT 23.685 77.545 23.855 77.715 ;
        RECT 24.145 77.545 24.315 77.715 ;
        RECT 24.605 77.545 24.775 77.715 ;
        RECT 25.065 77.545 25.235 77.715 ;
        RECT 25.525 77.545 25.695 77.715 ;
        RECT 25.985 77.545 26.155 77.715 ;
        RECT 26.445 77.545 26.615 77.715 ;
        RECT 26.905 77.545 27.075 77.715 ;
        RECT 27.365 77.545 27.535 77.715 ;
        RECT 27.825 77.545 27.995 77.715 ;
        RECT 28.285 77.545 28.455 77.715 ;
        RECT 28.745 77.545 28.915 77.715 ;
        RECT 29.205 77.545 29.375 77.715 ;
        RECT 29.665 77.545 29.835 77.715 ;
        RECT 30.125 77.545 30.295 77.715 ;
        RECT 30.585 77.545 30.755 77.715 ;
        RECT 31.045 77.545 31.215 77.715 ;
        RECT 31.505 77.545 31.675 77.715 ;
        RECT 31.965 77.545 32.135 77.715 ;
        RECT 32.425 77.545 32.595 77.715 ;
        RECT 32.885 77.545 33.055 77.715 ;
        RECT 33.345 77.545 33.515 77.715 ;
        RECT 33.805 77.545 33.975 77.715 ;
        RECT 34.265 77.545 34.435 77.715 ;
        RECT 34.725 77.545 34.895 77.715 ;
        RECT 35.185 77.545 35.355 77.715 ;
        RECT 35.645 77.545 35.815 77.715 ;
        RECT 36.105 77.545 36.275 77.715 ;
        RECT 36.565 77.545 36.735 77.715 ;
        RECT 37.025 77.545 37.195 77.715 ;
        RECT 37.485 77.545 37.655 77.715 ;
        RECT 37.945 77.545 38.115 77.715 ;
        RECT 38.405 77.545 38.575 77.715 ;
        RECT 38.865 77.545 39.035 77.715 ;
        RECT 39.325 77.545 39.495 77.715 ;
        RECT 39.785 77.545 39.955 77.715 ;
        RECT 40.245 77.545 40.415 77.715 ;
        RECT 40.705 77.545 40.875 77.715 ;
        RECT 41.165 77.545 41.335 77.715 ;
        RECT 41.625 77.545 41.795 77.715 ;
        RECT 42.085 77.545 42.255 77.715 ;
        RECT 42.545 77.545 42.715 77.715 ;
        RECT 43.005 77.545 43.175 77.715 ;
        RECT 43.465 77.545 43.635 77.715 ;
        RECT 43.925 77.545 44.095 77.715 ;
        RECT 44.385 77.545 44.555 77.715 ;
        RECT 44.845 77.545 45.015 77.715 ;
        RECT 45.305 77.545 45.475 77.715 ;
        RECT 45.765 77.545 45.935 77.715 ;
        RECT 46.225 77.545 46.395 77.715 ;
        RECT 46.685 77.545 46.855 77.715 ;
        RECT 47.145 77.545 47.315 77.715 ;
        RECT 47.605 77.545 47.775 77.715 ;
        RECT 48.065 77.545 48.235 77.715 ;
        RECT 48.525 77.545 48.695 77.715 ;
        RECT 48.985 77.545 49.155 77.715 ;
        RECT 49.445 77.545 49.615 77.715 ;
        RECT 49.905 77.545 50.075 77.715 ;
        RECT 50.365 77.545 50.535 77.715 ;
        RECT 50.825 77.545 50.995 77.715 ;
        RECT 51.285 77.545 51.455 77.715 ;
        RECT 51.745 77.545 51.915 77.715 ;
        RECT 52.205 77.545 52.375 77.715 ;
        RECT 52.665 77.545 52.835 77.715 ;
        RECT 53.125 77.545 53.295 77.715 ;
        RECT 53.585 77.545 53.755 77.715 ;
        RECT 54.045 77.545 54.215 77.715 ;
        RECT 54.505 77.545 54.675 77.715 ;
        RECT 54.965 77.545 55.135 77.715 ;
        RECT 55.425 77.545 55.595 77.715 ;
        RECT 55.885 77.545 56.055 77.715 ;
        RECT 56.345 77.545 56.515 77.715 ;
        RECT 56.805 77.545 56.975 77.715 ;
        RECT 57.265 77.545 57.435 77.715 ;
        RECT 57.725 77.545 57.895 77.715 ;
        RECT 58.185 77.545 58.355 77.715 ;
        RECT 58.645 77.545 58.815 77.715 ;
        RECT 59.105 77.545 59.275 77.715 ;
        RECT 59.565 77.545 59.735 77.715 ;
        RECT 60.025 77.545 60.195 77.715 ;
        RECT 60.485 77.545 60.655 77.715 ;
        RECT 60.945 77.545 61.115 77.715 ;
        RECT 61.405 77.545 61.575 77.715 ;
        RECT 61.865 77.545 62.035 77.715 ;
        RECT 62.325 77.545 62.495 77.715 ;
        RECT 62.785 77.545 62.955 77.715 ;
        RECT 63.245 77.545 63.415 77.715 ;
        RECT 63.705 77.545 63.875 77.715 ;
        RECT 64.165 77.545 64.335 77.715 ;
        RECT 64.625 77.545 64.795 77.715 ;
        RECT 65.085 77.545 65.255 77.715 ;
        RECT 65.545 77.545 65.715 77.715 ;
        RECT 66.005 77.545 66.175 77.715 ;
        RECT 66.465 77.545 66.635 77.715 ;
        RECT 66.925 77.545 67.095 77.715 ;
        RECT 67.385 77.545 67.555 77.715 ;
        RECT 67.845 77.545 68.015 77.715 ;
        RECT 68.305 77.545 68.475 77.715 ;
        RECT 68.765 77.545 68.935 77.715 ;
        RECT 69.225 77.545 69.395 77.715 ;
        RECT 69.685 77.545 69.855 77.715 ;
        RECT 70.145 77.545 70.315 77.715 ;
        RECT 70.605 77.545 70.775 77.715 ;
        RECT 71.065 77.545 71.235 77.715 ;
        RECT 71.525 77.545 71.695 77.715 ;
        RECT 71.985 77.545 72.155 77.715 ;
        RECT 72.445 77.545 72.615 77.715 ;
        RECT 72.905 77.545 73.075 77.715 ;
        RECT 73.365 77.545 73.535 77.715 ;
        RECT 73.825 77.545 73.995 77.715 ;
        RECT 74.285 77.545 74.455 77.715 ;
        RECT 74.745 77.545 74.915 77.715 ;
        RECT 75.205 77.545 75.375 77.715 ;
        RECT 75.665 77.545 75.835 77.715 ;
        RECT 76.125 77.545 76.295 77.715 ;
        RECT 76.585 77.545 76.755 77.715 ;
        RECT 77.045 77.545 77.215 77.715 ;
        RECT 77.505 77.545 77.675 77.715 ;
        RECT 77.965 77.545 78.135 77.715 ;
        RECT 78.425 77.545 78.595 77.715 ;
        RECT 78.885 77.545 79.055 77.715 ;
        RECT 79.345 77.545 79.515 77.715 ;
        RECT 79.805 77.545 79.975 77.715 ;
        RECT 80.265 77.545 80.435 77.715 ;
        RECT 80.725 77.545 80.895 77.715 ;
        RECT 81.185 77.545 81.355 77.715 ;
        RECT 81.645 77.545 81.815 77.715 ;
        RECT 82.105 77.545 82.275 77.715 ;
        RECT 82.565 77.545 82.735 77.715 ;
        RECT 83.025 77.545 83.195 77.715 ;
        RECT 83.485 77.545 83.655 77.715 ;
        RECT 83.945 77.545 84.115 77.715 ;
        RECT 84.405 77.545 84.575 77.715 ;
        RECT 84.865 77.545 85.035 77.715 ;
        RECT 85.325 77.545 85.495 77.715 ;
        RECT 85.785 77.545 85.955 77.715 ;
        RECT 86.245 77.545 86.415 77.715 ;
        RECT 86.705 77.545 86.875 77.715 ;
        RECT 87.165 77.545 87.335 77.715 ;
        RECT 87.625 77.545 87.795 77.715 ;
        RECT 88.085 77.545 88.255 77.715 ;
        RECT 88.545 77.545 88.715 77.715 ;
        RECT 89.005 77.545 89.175 77.715 ;
        RECT 89.465 77.545 89.635 77.715 ;
        RECT 89.925 77.545 90.095 77.715 ;
        RECT 90.385 77.545 90.555 77.715 ;
        RECT 90.845 77.545 91.015 77.715 ;
        RECT 91.305 77.545 91.475 77.715 ;
        RECT 91.765 77.545 91.935 77.715 ;
        RECT 92.225 77.545 92.395 77.715 ;
        RECT 92.685 77.545 92.855 77.715 ;
        RECT 93.145 77.545 93.315 77.715 ;
        RECT 93.605 77.545 93.775 77.715 ;
        RECT 94.065 77.545 94.235 77.715 ;
        RECT 94.525 77.545 94.695 77.715 ;
        RECT 94.985 77.545 95.155 77.715 ;
        RECT 95.445 77.545 95.615 77.715 ;
        RECT 95.905 77.545 96.075 77.715 ;
        RECT 96.365 77.545 96.535 77.715 ;
        RECT 96.825 77.545 96.995 77.715 ;
        RECT 97.285 77.545 97.455 77.715 ;
        RECT 97.745 77.545 97.915 77.715 ;
        RECT 98.205 77.545 98.375 77.715 ;
        RECT 98.665 77.545 98.835 77.715 ;
        RECT 99.125 77.545 99.295 77.715 ;
        RECT 99.585 77.545 99.755 77.715 ;
        RECT 100.045 77.545 100.215 77.715 ;
        RECT 100.505 77.545 100.675 77.715 ;
        RECT 100.965 77.545 101.135 77.715 ;
        RECT 101.425 77.545 101.595 77.715 ;
        RECT 101.885 77.545 102.055 77.715 ;
        RECT 102.345 77.545 102.515 77.715 ;
        RECT 102.805 77.545 102.975 77.715 ;
        RECT 103.265 77.545 103.435 77.715 ;
        RECT 103.725 77.545 103.895 77.715 ;
        RECT 104.185 77.545 104.355 77.715 ;
        RECT 104.645 77.545 104.815 77.715 ;
        RECT 105.105 77.545 105.275 77.715 ;
        RECT 105.565 77.545 105.735 77.715 ;
        RECT 106.025 77.545 106.195 77.715 ;
        RECT 106.485 77.545 106.655 77.715 ;
        RECT 106.945 77.545 107.115 77.715 ;
        RECT 107.405 77.545 107.575 77.715 ;
        RECT 107.865 77.545 108.035 77.715 ;
        RECT 108.325 77.545 108.495 77.715 ;
        RECT 108.785 77.545 108.955 77.715 ;
        RECT 109.245 77.545 109.415 77.715 ;
        RECT 109.705 77.545 109.875 77.715 ;
        RECT 110.165 77.545 110.335 77.715 ;
        RECT 110.625 77.545 110.795 77.715 ;
        RECT 111.085 77.545 111.255 77.715 ;
        RECT 111.545 77.545 111.715 77.715 ;
        RECT 112.005 77.545 112.175 77.715 ;
        RECT 112.465 77.545 112.635 77.715 ;
        RECT 112.925 77.545 113.095 77.715 ;
        RECT 113.385 77.545 113.555 77.715 ;
        RECT 113.845 77.545 114.015 77.715 ;
        RECT 114.305 77.545 114.475 77.715 ;
        RECT 114.765 77.545 114.935 77.715 ;
        RECT 115.225 77.545 115.395 77.715 ;
        RECT 115.685 77.545 115.855 77.715 ;
        RECT 116.145 77.545 116.315 77.715 ;
        RECT 116.605 77.545 116.775 77.715 ;
        RECT 117.065 77.545 117.235 77.715 ;
        RECT 117.525 77.545 117.695 77.715 ;
        RECT 117.985 77.545 118.155 77.715 ;
        RECT 118.445 77.545 118.615 77.715 ;
        RECT 118.905 77.545 119.075 77.715 ;
        RECT 119.365 77.545 119.535 77.715 ;
        RECT 119.825 77.545 119.995 77.715 ;
        RECT 120.285 77.545 120.455 77.715 ;
        RECT 120.745 77.545 120.915 77.715 ;
        RECT 121.205 77.545 121.375 77.715 ;
        RECT 121.665 77.545 121.835 77.715 ;
        RECT 122.125 77.545 122.295 77.715 ;
        RECT 122.585 77.545 122.755 77.715 ;
        RECT 123.045 77.545 123.215 77.715 ;
        RECT 123.505 77.545 123.675 77.715 ;
        RECT 123.965 77.545 124.135 77.715 ;
        RECT 124.425 77.545 124.595 77.715 ;
        RECT 124.885 77.545 125.055 77.715 ;
        RECT 125.345 77.545 125.515 77.715 ;
        RECT 125.805 77.545 125.975 77.715 ;
        RECT 126.265 77.545 126.435 77.715 ;
        RECT 126.725 77.545 126.895 77.715 ;
        RECT 127.185 77.545 127.355 77.715 ;
        RECT 127.645 77.545 127.815 77.715 ;
        RECT 128.105 77.545 128.275 77.715 ;
        RECT 128.565 77.545 128.735 77.715 ;
        RECT 129.025 77.545 129.195 77.715 ;
        RECT 129.485 77.545 129.655 77.715 ;
        RECT 129.945 77.545 130.115 77.715 ;
        RECT 130.405 77.545 130.575 77.715 ;
        RECT 130.865 77.545 131.035 77.715 ;
        RECT 131.325 77.545 131.495 77.715 ;
        RECT 131.785 77.545 131.955 77.715 ;
        RECT 132.245 77.545 132.415 77.715 ;
        RECT 132.705 77.545 132.875 77.715 ;
        RECT 133.165 77.545 133.335 77.715 ;
        RECT 133.625 77.545 133.795 77.715 ;
        RECT 134.085 77.545 134.255 77.715 ;
        RECT 134.545 77.545 134.715 77.715 ;
        RECT 135.005 77.545 135.175 77.715 ;
        RECT 135.465 77.545 135.635 77.715 ;
        RECT 135.925 77.545 136.095 77.715 ;
        RECT 136.385 77.545 136.555 77.715 ;
        RECT 136.845 77.545 137.015 77.715 ;
        RECT 137.305 77.545 137.475 77.715 ;
        RECT 137.765 77.545 137.935 77.715 ;
        RECT 138.225 77.545 138.395 77.715 ;
        RECT 138.685 77.545 138.855 77.715 ;
        RECT 139.145 77.545 139.315 77.715 ;
        RECT 139.605 77.545 139.775 77.715 ;
        RECT 140.065 77.545 140.235 77.715 ;
        RECT 140.525 77.545 140.695 77.715 ;
        RECT 140.985 77.545 141.155 77.715 ;
        RECT 141.445 77.545 141.615 77.715 ;
        RECT 141.905 77.545 142.075 77.715 ;
        RECT 142.365 77.545 142.535 77.715 ;
        RECT 142.825 77.545 142.995 77.715 ;
        RECT 143.285 77.545 143.455 77.715 ;
        RECT 143.745 77.545 143.915 77.715 ;
        RECT 144.205 77.545 144.375 77.715 ;
        RECT 144.665 77.545 144.835 77.715 ;
        RECT 145.125 77.545 145.295 77.715 ;
        RECT 145.585 77.545 145.755 77.715 ;
        RECT 146.045 77.545 146.215 77.715 ;
        RECT 146.505 77.545 146.675 77.715 ;
        RECT 146.965 77.545 147.135 77.715 ;
        RECT 147.425 77.545 147.595 77.715 ;
        RECT 147.885 77.545 148.055 77.715 ;
        RECT 148.345 77.545 148.515 77.715 ;
        RECT 148.805 77.545 148.975 77.715 ;
        RECT 149.265 77.545 149.435 77.715 ;
        RECT 149.725 77.545 149.895 77.715 ;
        RECT 150.185 77.545 150.355 77.715 ;
        RECT 11.265 74.825 11.435 74.995 ;
        RECT 11.725 74.825 11.895 74.995 ;
        RECT 12.185 74.825 12.355 74.995 ;
        RECT 12.645 74.825 12.815 74.995 ;
        RECT 13.105 74.825 13.275 74.995 ;
        RECT 13.565 74.825 13.735 74.995 ;
        RECT 14.025 74.825 14.195 74.995 ;
        RECT 14.485 74.825 14.655 74.995 ;
        RECT 14.945 74.825 15.115 74.995 ;
        RECT 15.405 74.825 15.575 74.995 ;
        RECT 15.865 74.825 16.035 74.995 ;
        RECT 16.325 74.825 16.495 74.995 ;
        RECT 16.785 74.825 16.955 74.995 ;
        RECT 17.245 74.825 17.415 74.995 ;
        RECT 17.705 74.825 17.875 74.995 ;
        RECT 18.165 74.825 18.335 74.995 ;
        RECT 18.625 74.825 18.795 74.995 ;
        RECT 19.085 74.825 19.255 74.995 ;
        RECT 19.545 74.825 19.715 74.995 ;
        RECT 20.005 74.825 20.175 74.995 ;
        RECT 20.465 74.825 20.635 74.995 ;
        RECT 20.925 74.825 21.095 74.995 ;
        RECT 21.385 74.825 21.555 74.995 ;
        RECT 21.845 74.825 22.015 74.995 ;
        RECT 22.305 74.825 22.475 74.995 ;
        RECT 22.765 74.825 22.935 74.995 ;
        RECT 23.225 74.825 23.395 74.995 ;
        RECT 23.685 74.825 23.855 74.995 ;
        RECT 24.145 74.825 24.315 74.995 ;
        RECT 24.605 74.825 24.775 74.995 ;
        RECT 25.065 74.825 25.235 74.995 ;
        RECT 25.525 74.825 25.695 74.995 ;
        RECT 25.985 74.825 26.155 74.995 ;
        RECT 26.445 74.825 26.615 74.995 ;
        RECT 26.905 74.825 27.075 74.995 ;
        RECT 27.365 74.825 27.535 74.995 ;
        RECT 27.825 74.825 27.995 74.995 ;
        RECT 28.285 74.825 28.455 74.995 ;
        RECT 28.745 74.825 28.915 74.995 ;
        RECT 29.205 74.825 29.375 74.995 ;
        RECT 29.665 74.825 29.835 74.995 ;
        RECT 30.125 74.825 30.295 74.995 ;
        RECT 30.585 74.825 30.755 74.995 ;
        RECT 31.045 74.825 31.215 74.995 ;
        RECT 31.505 74.825 31.675 74.995 ;
        RECT 31.965 74.825 32.135 74.995 ;
        RECT 32.425 74.825 32.595 74.995 ;
        RECT 32.885 74.825 33.055 74.995 ;
        RECT 33.345 74.825 33.515 74.995 ;
        RECT 33.805 74.825 33.975 74.995 ;
        RECT 34.265 74.825 34.435 74.995 ;
        RECT 34.725 74.825 34.895 74.995 ;
        RECT 35.185 74.825 35.355 74.995 ;
        RECT 35.645 74.825 35.815 74.995 ;
        RECT 36.105 74.825 36.275 74.995 ;
        RECT 36.565 74.825 36.735 74.995 ;
        RECT 37.025 74.825 37.195 74.995 ;
        RECT 37.485 74.825 37.655 74.995 ;
        RECT 37.945 74.825 38.115 74.995 ;
        RECT 38.405 74.825 38.575 74.995 ;
        RECT 38.865 74.825 39.035 74.995 ;
        RECT 39.325 74.825 39.495 74.995 ;
        RECT 39.785 74.825 39.955 74.995 ;
        RECT 40.245 74.825 40.415 74.995 ;
        RECT 40.705 74.825 40.875 74.995 ;
        RECT 41.165 74.825 41.335 74.995 ;
        RECT 41.625 74.825 41.795 74.995 ;
        RECT 42.085 74.825 42.255 74.995 ;
        RECT 42.545 74.825 42.715 74.995 ;
        RECT 43.005 74.825 43.175 74.995 ;
        RECT 43.465 74.825 43.635 74.995 ;
        RECT 43.925 74.825 44.095 74.995 ;
        RECT 44.385 74.825 44.555 74.995 ;
        RECT 44.845 74.825 45.015 74.995 ;
        RECT 45.305 74.825 45.475 74.995 ;
        RECT 45.765 74.825 45.935 74.995 ;
        RECT 46.225 74.825 46.395 74.995 ;
        RECT 46.685 74.825 46.855 74.995 ;
        RECT 47.145 74.825 47.315 74.995 ;
        RECT 47.605 74.825 47.775 74.995 ;
        RECT 48.065 74.825 48.235 74.995 ;
        RECT 48.525 74.825 48.695 74.995 ;
        RECT 48.985 74.825 49.155 74.995 ;
        RECT 49.445 74.825 49.615 74.995 ;
        RECT 49.905 74.825 50.075 74.995 ;
        RECT 50.365 74.825 50.535 74.995 ;
        RECT 50.825 74.825 50.995 74.995 ;
        RECT 51.285 74.825 51.455 74.995 ;
        RECT 51.745 74.825 51.915 74.995 ;
        RECT 52.205 74.825 52.375 74.995 ;
        RECT 52.665 74.825 52.835 74.995 ;
        RECT 53.125 74.825 53.295 74.995 ;
        RECT 53.585 74.825 53.755 74.995 ;
        RECT 54.045 74.825 54.215 74.995 ;
        RECT 54.505 74.825 54.675 74.995 ;
        RECT 54.965 74.825 55.135 74.995 ;
        RECT 55.425 74.825 55.595 74.995 ;
        RECT 55.885 74.825 56.055 74.995 ;
        RECT 56.345 74.825 56.515 74.995 ;
        RECT 56.805 74.825 56.975 74.995 ;
        RECT 57.265 74.825 57.435 74.995 ;
        RECT 57.725 74.825 57.895 74.995 ;
        RECT 58.185 74.825 58.355 74.995 ;
        RECT 58.645 74.825 58.815 74.995 ;
        RECT 59.105 74.825 59.275 74.995 ;
        RECT 59.565 74.825 59.735 74.995 ;
        RECT 60.025 74.825 60.195 74.995 ;
        RECT 60.485 74.825 60.655 74.995 ;
        RECT 60.945 74.825 61.115 74.995 ;
        RECT 61.405 74.825 61.575 74.995 ;
        RECT 61.865 74.825 62.035 74.995 ;
        RECT 62.325 74.825 62.495 74.995 ;
        RECT 62.785 74.825 62.955 74.995 ;
        RECT 63.245 74.825 63.415 74.995 ;
        RECT 63.705 74.825 63.875 74.995 ;
        RECT 64.165 74.825 64.335 74.995 ;
        RECT 64.625 74.825 64.795 74.995 ;
        RECT 65.085 74.825 65.255 74.995 ;
        RECT 65.545 74.825 65.715 74.995 ;
        RECT 66.005 74.825 66.175 74.995 ;
        RECT 66.465 74.825 66.635 74.995 ;
        RECT 66.925 74.825 67.095 74.995 ;
        RECT 67.385 74.825 67.555 74.995 ;
        RECT 67.845 74.825 68.015 74.995 ;
        RECT 68.305 74.825 68.475 74.995 ;
        RECT 68.765 74.825 68.935 74.995 ;
        RECT 69.225 74.825 69.395 74.995 ;
        RECT 69.685 74.825 69.855 74.995 ;
        RECT 70.145 74.825 70.315 74.995 ;
        RECT 70.605 74.825 70.775 74.995 ;
        RECT 71.065 74.825 71.235 74.995 ;
        RECT 71.525 74.825 71.695 74.995 ;
        RECT 71.985 74.825 72.155 74.995 ;
        RECT 72.445 74.825 72.615 74.995 ;
        RECT 72.905 74.825 73.075 74.995 ;
        RECT 73.365 74.825 73.535 74.995 ;
        RECT 73.825 74.825 73.995 74.995 ;
        RECT 74.285 74.825 74.455 74.995 ;
        RECT 74.745 74.825 74.915 74.995 ;
        RECT 75.205 74.825 75.375 74.995 ;
        RECT 75.665 74.825 75.835 74.995 ;
        RECT 76.125 74.825 76.295 74.995 ;
        RECT 76.585 74.825 76.755 74.995 ;
        RECT 77.045 74.825 77.215 74.995 ;
        RECT 77.505 74.825 77.675 74.995 ;
        RECT 77.965 74.825 78.135 74.995 ;
        RECT 78.425 74.825 78.595 74.995 ;
        RECT 78.885 74.825 79.055 74.995 ;
        RECT 79.345 74.825 79.515 74.995 ;
        RECT 79.805 74.825 79.975 74.995 ;
        RECT 80.265 74.825 80.435 74.995 ;
        RECT 80.725 74.825 80.895 74.995 ;
        RECT 81.185 74.825 81.355 74.995 ;
        RECT 81.645 74.825 81.815 74.995 ;
        RECT 82.105 74.825 82.275 74.995 ;
        RECT 82.565 74.825 82.735 74.995 ;
        RECT 83.025 74.825 83.195 74.995 ;
        RECT 83.485 74.825 83.655 74.995 ;
        RECT 83.945 74.825 84.115 74.995 ;
        RECT 84.405 74.825 84.575 74.995 ;
        RECT 84.865 74.825 85.035 74.995 ;
        RECT 85.325 74.825 85.495 74.995 ;
        RECT 85.785 74.825 85.955 74.995 ;
        RECT 86.245 74.825 86.415 74.995 ;
        RECT 86.705 74.825 86.875 74.995 ;
        RECT 87.165 74.825 87.335 74.995 ;
        RECT 87.625 74.825 87.795 74.995 ;
        RECT 88.085 74.825 88.255 74.995 ;
        RECT 88.545 74.825 88.715 74.995 ;
        RECT 89.005 74.825 89.175 74.995 ;
        RECT 89.465 74.825 89.635 74.995 ;
        RECT 89.925 74.825 90.095 74.995 ;
        RECT 90.385 74.825 90.555 74.995 ;
        RECT 90.845 74.825 91.015 74.995 ;
        RECT 91.305 74.825 91.475 74.995 ;
        RECT 91.765 74.825 91.935 74.995 ;
        RECT 92.225 74.825 92.395 74.995 ;
        RECT 92.685 74.825 92.855 74.995 ;
        RECT 93.145 74.825 93.315 74.995 ;
        RECT 93.605 74.825 93.775 74.995 ;
        RECT 94.065 74.825 94.235 74.995 ;
        RECT 94.525 74.825 94.695 74.995 ;
        RECT 94.985 74.825 95.155 74.995 ;
        RECT 95.445 74.825 95.615 74.995 ;
        RECT 95.905 74.825 96.075 74.995 ;
        RECT 96.365 74.825 96.535 74.995 ;
        RECT 96.825 74.825 96.995 74.995 ;
        RECT 97.285 74.825 97.455 74.995 ;
        RECT 97.745 74.825 97.915 74.995 ;
        RECT 98.205 74.825 98.375 74.995 ;
        RECT 98.665 74.825 98.835 74.995 ;
        RECT 99.125 74.825 99.295 74.995 ;
        RECT 99.585 74.825 99.755 74.995 ;
        RECT 100.045 74.825 100.215 74.995 ;
        RECT 100.505 74.825 100.675 74.995 ;
        RECT 100.965 74.825 101.135 74.995 ;
        RECT 101.425 74.825 101.595 74.995 ;
        RECT 101.885 74.825 102.055 74.995 ;
        RECT 102.345 74.825 102.515 74.995 ;
        RECT 102.805 74.825 102.975 74.995 ;
        RECT 103.265 74.825 103.435 74.995 ;
        RECT 103.725 74.825 103.895 74.995 ;
        RECT 104.185 74.825 104.355 74.995 ;
        RECT 104.645 74.825 104.815 74.995 ;
        RECT 105.105 74.825 105.275 74.995 ;
        RECT 105.565 74.825 105.735 74.995 ;
        RECT 106.025 74.825 106.195 74.995 ;
        RECT 106.485 74.825 106.655 74.995 ;
        RECT 106.945 74.825 107.115 74.995 ;
        RECT 107.405 74.825 107.575 74.995 ;
        RECT 107.865 74.825 108.035 74.995 ;
        RECT 108.325 74.825 108.495 74.995 ;
        RECT 108.785 74.825 108.955 74.995 ;
        RECT 109.245 74.825 109.415 74.995 ;
        RECT 109.705 74.825 109.875 74.995 ;
        RECT 110.165 74.825 110.335 74.995 ;
        RECT 110.625 74.825 110.795 74.995 ;
        RECT 111.085 74.825 111.255 74.995 ;
        RECT 111.545 74.825 111.715 74.995 ;
        RECT 112.005 74.825 112.175 74.995 ;
        RECT 112.465 74.825 112.635 74.995 ;
        RECT 112.925 74.825 113.095 74.995 ;
        RECT 113.385 74.825 113.555 74.995 ;
        RECT 113.845 74.825 114.015 74.995 ;
        RECT 114.305 74.825 114.475 74.995 ;
        RECT 114.765 74.825 114.935 74.995 ;
        RECT 115.225 74.825 115.395 74.995 ;
        RECT 115.685 74.825 115.855 74.995 ;
        RECT 116.145 74.825 116.315 74.995 ;
        RECT 116.605 74.825 116.775 74.995 ;
        RECT 117.065 74.825 117.235 74.995 ;
        RECT 117.525 74.825 117.695 74.995 ;
        RECT 117.985 74.825 118.155 74.995 ;
        RECT 118.445 74.825 118.615 74.995 ;
        RECT 118.905 74.825 119.075 74.995 ;
        RECT 119.365 74.825 119.535 74.995 ;
        RECT 119.825 74.825 119.995 74.995 ;
        RECT 120.285 74.825 120.455 74.995 ;
        RECT 120.745 74.825 120.915 74.995 ;
        RECT 121.205 74.825 121.375 74.995 ;
        RECT 121.665 74.825 121.835 74.995 ;
        RECT 122.125 74.825 122.295 74.995 ;
        RECT 122.585 74.825 122.755 74.995 ;
        RECT 123.045 74.825 123.215 74.995 ;
        RECT 123.505 74.825 123.675 74.995 ;
        RECT 123.965 74.825 124.135 74.995 ;
        RECT 124.425 74.825 124.595 74.995 ;
        RECT 124.885 74.825 125.055 74.995 ;
        RECT 125.345 74.825 125.515 74.995 ;
        RECT 125.805 74.825 125.975 74.995 ;
        RECT 126.265 74.825 126.435 74.995 ;
        RECT 126.725 74.825 126.895 74.995 ;
        RECT 127.185 74.825 127.355 74.995 ;
        RECT 127.645 74.825 127.815 74.995 ;
        RECT 128.105 74.825 128.275 74.995 ;
        RECT 128.565 74.825 128.735 74.995 ;
        RECT 129.025 74.825 129.195 74.995 ;
        RECT 129.485 74.825 129.655 74.995 ;
        RECT 129.945 74.825 130.115 74.995 ;
        RECT 130.405 74.825 130.575 74.995 ;
        RECT 130.865 74.825 131.035 74.995 ;
        RECT 131.325 74.825 131.495 74.995 ;
        RECT 131.785 74.825 131.955 74.995 ;
        RECT 132.245 74.825 132.415 74.995 ;
        RECT 132.705 74.825 132.875 74.995 ;
        RECT 133.165 74.825 133.335 74.995 ;
        RECT 133.625 74.825 133.795 74.995 ;
        RECT 134.085 74.825 134.255 74.995 ;
        RECT 134.545 74.825 134.715 74.995 ;
        RECT 135.005 74.825 135.175 74.995 ;
        RECT 135.465 74.825 135.635 74.995 ;
        RECT 135.925 74.825 136.095 74.995 ;
        RECT 136.385 74.825 136.555 74.995 ;
        RECT 136.845 74.825 137.015 74.995 ;
        RECT 137.305 74.825 137.475 74.995 ;
        RECT 137.765 74.825 137.935 74.995 ;
        RECT 138.225 74.825 138.395 74.995 ;
        RECT 138.685 74.825 138.855 74.995 ;
        RECT 139.145 74.825 139.315 74.995 ;
        RECT 139.605 74.825 139.775 74.995 ;
        RECT 140.065 74.825 140.235 74.995 ;
        RECT 140.525 74.825 140.695 74.995 ;
        RECT 140.985 74.825 141.155 74.995 ;
        RECT 141.445 74.825 141.615 74.995 ;
        RECT 141.905 74.825 142.075 74.995 ;
        RECT 142.365 74.825 142.535 74.995 ;
        RECT 142.825 74.825 142.995 74.995 ;
        RECT 143.285 74.825 143.455 74.995 ;
        RECT 143.745 74.825 143.915 74.995 ;
        RECT 144.205 74.825 144.375 74.995 ;
        RECT 144.665 74.825 144.835 74.995 ;
        RECT 145.125 74.825 145.295 74.995 ;
        RECT 145.585 74.825 145.755 74.995 ;
        RECT 146.045 74.825 146.215 74.995 ;
        RECT 146.505 74.825 146.675 74.995 ;
        RECT 146.965 74.825 147.135 74.995 ;
        RECT 147.425 74.825 147.595 74.995 ;
        RECT 147.885 74.825 148.055 74.995 ;
        RECT 148.345 74.825 148.515 74.995 ;
        RECT 148.805 74.825 148.975 74.995 ;
        RECT 149.265 74.825 149.435 74.995 ;
        RECT 149.725 74.825 149.895 74.995 ;
        RECT 150.185 74.825 150.355 74.995 ;
        RECT 56.100 51.140 84.500 52.080 ;
        RECT 55.040 50.560 84.500 51.140 ;
        RECT 55.040 46.070 60.510 50.560 ;
        RECT 62.035 49.320 62.915 49.490 ;
        RECT 61.570 47.340 61.740 49.180 ;
        RECT 63.210 47.340 63.380 49.180 ;
        RECT 62.035 47.030 62.915 47.200 ;
        RECT 61.570 45.050 61.740 46.890 ;
        RECT 63.210 45.050 63.380 46.890 ;
        RECT 62.035 44.740 62.915 44.910 ;
        RECT 61.570 42.760 61.740 44.600 ;
        RECT 63.210 42.760 63.380 44.600 ;
        RECT 62.035 42.450 62.915 42.620 ;
        RECT 61.570 40.470 61.740 42.310 ;
        RECT 63.210 40.470 63.380 42.310 ;
        RECT 62.035 40.160 62.915 40.330 ;
        RECT 61.570 38.180 61.740 40.020 ;
        RECT 63.210 38.180 63.380 40.020 ;
        RECT 62.035 37.870 62.915 38.040 ;
        RECT 61.570 35.890 61.740 37.730 ;
        RECT 63.210 35.890 63.380 37.730 ;
        RECT 62.035 35.580 62.915 35.750 ;
        RECT 64.695 49.320 65.575 49.490 ;
        RECT 64.230 47.340 64.400 49.180 ;
        RECT 65.870 47.340 66.040 49.180 ;
        RECT 67.030 48.190 77.340 50.560 ;
        RECT 96.080 50.740 105.390 51.570 ;
        RECT 118.330 50.740 146.730 51.680 ;
        RECT 78.805 49.310 79.685 49.480 ;
        RECT 78.340 48.830 78.510 49.170 ;
        RECT 79.980 48.830 80.150 49.170 ;
        RECT 78.805 48.520 79.685 48.690 ;
        RECT 64.695 47.030 65.575 47.200 ;
        RECT 64.230 45.050 64.400 46.890 ;
        RECT 65.870 45.050 66.040 46.890 ;
        RECT 64.695 44.740 65.575 44.910 ;
        RECT 64.230 42.760 64.400 44.600 ;
        RECT 65.870 42.760 66.040 44.600 ;
        RECT 78.340 48.040 78.510 48.380 ;
        RECT 79.980 48.040 80.150 48.380 ;
        RECT 78.805 47.730 79.685 47.900 ;
        RECT 78.340 47.250 78.510 47.590 ;
        RECT 79.980 47.250 80.150 47.590 ;
        RECT 78.805 46.940 79.685 47.110 ;
        RECT 78.340 46.460 78.510 46.800 ;
        RECT 79.980 46.460 80.150 46.800 ;
        RECT 78.805 46.150 79.685 46.320 ;
        RECT 78.340 45.670 78.510 46.010 ;
        RECT 79.980 45.670 80.150 46.010 ;
        RECT 78.805 45.360 79.685 45.530 ;
        RECT 78.340 44.880 78.510 45.220 ;
        RECT 79.980 44.880 80.150 45.220 ;
        RECT 78.805 44.570 79.685 44.740 ;
        RECT 78.340 44.090 78.510 44.430 ;
        RECT 79.980 44.090 80.150 44.430 ;
        RECT 78.805 43.780 79.685 43.950 ;
        RECT 64.695 42.450 65.575 42.620 ;
        RECT 64.230 40.470 64.400 42.310 ;
        RECT 65.870 40.470 66.040 42.310 ;
        RECT 64.695 40.160 65.575 40.330 ;
        RECT 64.230 38.180 64.400 40.020 ;
        RECT 65.870 38.180 66.040 40.020 ;
        RECT 64.695 37.870 65.575 38.040 ;
        RECT 64.230 35.890 64.400 37.730 ;
        RECT 65.870 35.890 66.040 37.730 ;
        RECT 64.695 35.580 65.575 35.750 ;
        RECT 73.620 42.150 74.500 42.320 ;
        RECT 73.200 40.170 73.370 42.010 ;
        RECT 74.750 40.170 74.920 42.010 ;
        RECT 73.620 39.860 74.500 40.030 ;
        RECT 73.200 37.880 73.370 39.720 ;
        RECT 74.750 37.880 74.920 39.720 ;
        RECT 73.620 37.570 74.500 37.740 ;
        RECT 73.200 35.590 73.370 37.430 ;
        RECT 74.750 35.590 74.920 37.430 ;
        RECT 73.620 35.280 74.500 35.450 ;
        RECT 62.650 33.600 62.990 33.770 ;
        RECT 62.340 30.970 62.510 33.350 ;
        RECT 63.130 30.970 63.300 33.350 ;
        RECT 62.650 30.550 62.990 30.720 ;
        RECT 64.580 33.600 64.920 33.770 ;
        RECT 64.270 30.970 64.440 33.350 ;
        RECT 65.060 30.970 65.230 33.350 ;
        RECT 64.580 30.550 64.920 30.720 ;
        RECT 73.200 33.300 73.370 35.140 ;
        RECT 74.750 33.300 74.920 35.140 ;
        RECT 73.620 32.990 74.500 33.160 ;
        RECT 73.200 31.010 73.370 32.850 ;
        RECT 74.750 31.010 74.920 32.850 ;
        RECT 78.340 43.300 78.510 43.640 ;
        RECT 79.980 43.300 80.150 43.640 ;
        RECT 78.805 42.990 79.685 43.160 ;
        RECT 78.340 42.510 78.510 42.850 ;
        RECT 79.980 42.510 80.150 42.850 ;
        RECT 78.805 42.200 79.685 42.370 ;
        RECT 78.340 41.720 78.510 42.060 ;
        RECT 79.980 41.720 80.150 42.060 ;
        RECT 78.805 41.410 79.685 41.580 ;
        RECT 78.340 40.930 78.510 41.270 ;
        RECT 79.980 40.930 80.150 41.270 ;
        RECT 78.805 40.620 79.685 40.790 ;
        RECT 78.340 40.140 78.510 40.480 ;
        RECT 79.980 40.140 80.150 40.480 ;
        RECT 78.805 39.830 79.685 40.000 ;
        RECT 78.340 39.350 78.510 39.690 ;
        RECT 79.980 39.350 80.150 39.690 ;
        RECT 78.805 39.040 79.685 39.210 ;
        RECT 78.340 38.560 78.510 38.900 ;
        RECT 79.980 38.560 80.150 38.900 ;
        RECT 78.805 38.250 79.685 38.420 ;
        RECT 78.340 37.770 78.510 38.110 ;
        RECT 79.980 37.770 80.150 38.110 ;
        RECT 78.805 37.460 79.685 37.630 ;
        RECT 78.340 36.980 78.510 37.320 ;
        RECT 79.980 36.980 80.150 37.320 ;
        RECT 78.805 36.670 79.685 36.840 ;
        RECT 78.340 36.190 78.510 36.530 ;
        RECT 79.980 36.190 80.150 36.530 ;
        RECT 78.805 35.880 79.685 36.050 ;
        RECT 78.340 35.400 78.510 35.740 ;
        RECT 79.980 35.400 80.150 35.740 ;
        RECT 78.805 35.090 79.685 35.260 ;
        RECT 78.340 34.610 78.510 34.950 ;
        RECT 79.980 34.610 80.150 34.950 ;
        RECT 78.805 34.300 79.685 34.470 ;
        RECT 78.340 33.820 78.510 34.160 ;
        RECT 79.980 33.820 80.150 34.160 ;
        RECT 78.805 33.510 79.685 33.680 ;
        RECT 100.310 47.075 100.500 49.060 ;
        RECT 100.310 42.280 100.500 44.265 ;
        RECT 95.850 39.280 97.690 39.450 ;
        RECT 98.140 39.280 99.980 39.450 ;
        RECT 100.430 39.280 102.270 39.450 ;
        RECT 102.720 39.280 104.560 39.450 ;
        RECT 95.540 38.150 95.710 39.030 ;
        RECT 97.830 38.150 98.000 39.030 ;
        RECT 100.120 38.150 100.290 39.030 ;
        RECT 102.410 38.150 102.580 39.030 ;
        RECT 104.700 38.150 104.870 39.030 ;
        RECT 95.850 37.730 97.690 37.900 ;
        RECT 98.140 37.730 99.980 37.900 ;
        RECT 100.430 37.730 102.270 37.900 ;
        RECT 102.720 37.730 104.560 37.900 ;
        RECT 95.250 34.630 105.560 36.550 ;
        RECT 117.270 50.160 146.730 50.740 ;
        RECT 117.270 45.670 122.740 50.160 ;
        RECT 124.265 48.920 125.145 49.090 ;
        RECT 123.800 46.940 123.970 48.780 ;
        RECT 125.440 46.940 125.610 48.780 ;
        RECT 124.265 46.630 125.145 46.800 ;
        RECT 123.800 44.650 123.970 46.490 ;
        RECT 125.440 44.650 125.610 46.490 ;
        RECT 124.265 44.340 125.145 44.510 ;
        RECT 123.800 42.360 123.970 44.200 ;
        RECT 125.440 42.360 125.610 44.200 ;
        RECT 124.265 42.050 125.145 42.220 ;
        RECT 123.800 40.070 123.970 41.910 ;
        RECT 125.440 40.070 125.610 41.910 ;
        RECT 124.265 39.760 125.145 39.930 ;
        RECT 123.800 37.780 123.970 39.620 ;
        RECT 125.440 37.780 125.610 39.620 ;
        RECT 124.265 37.470 125.145 37.640 ;
        RECT 123.800 35.490 123.970 37.330 ;
        RECT 125.440 35.490 125.610 37.330 ;
        RECT 124.265 35.180 125.145 35.350 ;
        RECT 126.925 48.920 127.805 49.090 ;
        RECT 126.460 46.940 126.630 48.780 ;
        RECT 128.100 46.940 128.270 48.780 ;
        RECT 129.260 47.790 139.570 50.160 ;
        RECT 141.035 48.910 141.915 49.080 ;
        RECT 140.570 48.430 140.740 48.770 ;
        RECT 142.210 48.430 142.380 48.770 ;
        RECT 141.035 48.120 141.915 48.290 ;
        RECT 126.925 46.630 127.805 46.800 ;
        RECT 126.460 44.650 126.630 46.490 ;
        RECT 128.100 44.650 128.270 46.490 ;
        RECT 126.925 44.340 127.805 44.510 ;
        RECT 126.460 42.360 126.630 44.200 ;
        RECT 128.100 42.360 128.270 44.200 ;
        RECT 140.570 47.640 140.740 47.980 ;
        RECT 142.210 47.640 142.380 47.980 ;
        RECT 141.035 47.330 141.915 47.500 ;
        RECT 140.570 46.850 140.740 47.190 ;
        RECT 142.210 46.850 142.380 47.190 ;
        RECT 141.035 46.540 141.915 46.710 ;
        RECT 140.570 46.060 140.740 46.400 ;
        RECT 142.210 46.060 142.380 46.400 ;
        RECT 141.035 45.750 141.915 45.920 ;
        RECT 140.570 45.270 140.740 45.610 ;
        RECT 142.210 45.270 142.380 45.610 ;
        RECT 141.035 44.960 141.915 45.130 ;
        RECT 140.570 44.480 140.740 44.820 ;
        RECT 142.210 44.480 142.380 44.820 ;
        RECT 141.035 44.170 141.915 44.340 ;
        RECT 140.570 43.690 140.740 44.030 ;
        RECT 142.210 43.690 142.380 44.030 ;
        RECT 141.035 43.380 141.915 43.550 ;
        RECT 126.925 42.050 127.805 42.220 ;
        RECT 126.460 40.070 126.630 41.910 ;
        RECT 128.100 40.070 128.270 41.910 ;
        RECT 126.925 39.760 127.805 39.930 ;
        RECT 126.460 37.780 126.630 39.620 ;
        RECT 128.100 37.780 128.270 39.620 ;
        RECT 126.925 37.470 127.805 37.640 ;
        RECT 126.460 35.490 126.630 37.330 ;
        RECT 128.100 35.490 128.270 37.330 ;
        RECT 126.925 35.180 127.805 35.350 ;
        RECT 135.850 41.750 136.730 41.920 ;
        RECT 135.430 39.770 135.600 41.610 ;
        RECT 136.980 39.770 137.150 41.610 ;
        RECT 135.850 39.460 136.730 39.630 ;
        RECT 135.430 37.480 135.600 39.320 ;
        RECT 136.980 37.480 137.150 39.320 ;
        RECT 135.850 37.170 136.730 37.340 ;
        RECT 135.430 35.190 135.600 37.030 ;
        RECT 136.980 35.190 137.150 37.030 ;
        RECT 135.850 34.880 136.730 35.050 ;
        RECT 73.620 30.700 74.500 30.870 ;
        RECT 73.200 28.720 73.370 30.560 ;
        RECT 74.750 28.720 74.920 30.560 ;
        RECT 73.620 28.410 74.500 28.580 ;
        RECT 55.910 26.660 57.750 26.830 ;
        RECT 58.200 26.660 60.040 26.830 ;
        RECT 60.490 26.660 62.330 26.830 ;
        RECT 62.780 26.660 64.620 26.830 ;
        RECT 55.600 25.530 55.770 26.410 ;
        RECT 57.890 25.530 58.060 26.410 ;
        RECT 60.180 25.530 60.350 26.410 ;
        RECT 62.470 25.530 62.640 26.410 ;
        RECT 64.760 25.530 64.930 26.410 ;
        RECT 73.200 26.430 73.370 28.270 ;
        RECT 74.750 26.430 74.920 28.270 ;
        RECT 73.620 26.120 74.500 26.290 ;
        RECT 55.910 25.110 57.750 25.280 ;
        RECT 58.200 25.110 60.040 25.280 ;
        RECT 60.490 25.110 62.330 25.280 ;
        RECT 62.780 25.110 64.620 25.280 ;
        RECT 70.540 24.250 84.430 25.350 ;
        RECT 56.040 22.730 84.440 24.250 ;
        RECT 124.880 33.200 125.220 33.370 ;
        RECT 124.570 30.570 124.740 32.950 ;
        RECT 125.360 30.570 125.530 32.950 ;
        RECT 124.880 30.150 125.220 30.320 ;
        RECT 126.810 33.200 127.150 33.370 ;
        RECT 126.500 30.570 126.670 32.950 ;
        RECT 127.290 30.570 127.460 32.950 ;
        RECT 126.810 30.150 127.150 30.320 ;
        RECT 135.430 32.900 135.600 34.740 ;
        RECT 136.980 32.900 137.150 34.740 ;
        RECT 135.850 32.590 136.730 32.760 ;
        RECT 135.430 30.610 135.600 32.450 ;
        RECT 136.980 30.610 137.150 32.450 ;
        RECT 140.570 42.900 140.740 43.240 ;
        RECT 142.210 42.900 142.380 43.240 ;
        RECT 141.035 42.590 141.915 42.760 ;
        RECT 140.570 42.110 140.740 42.450 ;
        RECT 142.210 42.110 142.380 42.450 ;
        RECT 141.035 41.800 141.915 41.970 ;
        RECT 140.570 41.320 140.740 41.660 ;
        RECT 142.210 41.320 142.380 41.660 ;
        RECT 141.035 41.010 141.915 41.180 ;
        RECT 140.570 40.530 140.740 40.870 ;
        RECT 142.210 40.530 142.380 40.870 ;
        RECT 141.035 40.220 141.915 40.390 ;
        RECT 140.570 39.740 140.740 40.080 ;
        RECT 142.210 39.740 142.380 40.080 ;
        RECT 141.035 39.430 141.915 39.600 ;
        RECT 140.570 38.950 140.740 39.290 ;
        RECT 142.210 38.950 142.380 39.290 ;
        RECT 141.035 38.640 141.915 38.810 ;
        RECT 140.570 38.160 140.740 38.500 ;
        RECT 142.210 38.160 142.380 38.500 ;
        RECT 141.035 37.850 141.915 38.020 ;
        RECT 140.570 37.370 140.740 37.710 ;
        RECT 142.210 37.370 142.380 37.710 ;
        RECT 141.035 37.060 141.915 37.230 ;
        RECT 140.570 36.580 140.740 36.920 ;
        RECT 142.210 36.580 142.380 36.920 ;
        RECT 141.035 36.270 141.915 36.440 ;
        RECT 140.570 35.790 140.740 36.130 ;
        RECT 142.210 35.790 142.380 36.130 ;
        RECT 141.035 35.480 141.915 35.650 ;
        RECT 140.570 35.000 140.740 35.340 ;
        RECT 142.210 35.000 142.380 35.340 ;
        RECT 141.035 34.690 141.915 34.860 ;
        RECT 140.570 34.210 140.740 34.550 ;
        RECT 142.210 34.210 142.380 34.550 ;
        RECT 141.035 33.900 141.915 34.070 ;
        RECT 140.570 33.420 140.740 33.760 ;
        RECT 142.210 33.420 142.380 33.760 ;
        RECT 141.035 33.110 141.915 33.280 ;
        RECT 135.850 30.300 136.730 30.470 ;
        RECT 135.430 28.320 135.600 30.160 ;
        RECT 136.980 28.320 137.150 30.160 ;
        RECT 135.850 28.010 136.730 28.180 ;
        RECT 118.140 26.260 119.980 26.430 ;
        RECT 120.430 26.260 122.270 26.430 ;
        RECT 122.720 26.260 124.560 26.430 ;
        RECT 125.010 26.260 126.850 26.430 ;
        RECT 117.830 25.130 118.000 26.010 ;
        RECT 120.120 25.130 120.290 26.010 ;
        RECT 122.410 25.130 122.580 26.010 ;
        RECT 124.700 25.130 124.870 26.010 ;
        RECT 126.990 25.130 127.160 26.010 ;
        RECT 135.430 26.030 135.600 27.870 ;
        RECT 136.980 26.030 137.150 27.870 ;
        RECT 135.850 25.720 136.730 25.890 ;
        RECT 118.140 24.710 119.980 24.880 ;
        RECT 120.430 24.710 122.270 24.880 ;
        RECT 122.720 24.710 124.560 24.880 ;
        RECT 125.010 24.710 126.850 24.880 ;
        RECT 132.770 23.850 146.660 24.950 ;
        RECT 118.270 22.330 146.670 23.850 ;
      LAYER met1 ;
        RECT 11.120 213.390 150.500 213.870 ;
        RECT 65.025 213.190 65.315 213.235 ;
        RECT 65.470 213.190 65.790 213.250 ;
        RECT 65.025 213.050 65.790 213.190 ;
        RECT 65.025 213.005 65.315 213.050 ;
        RECT 65.470 212.990 65.790 213.050 ;
        RECT 105.950 212.990 106.270 213.250 ;
        RECT 106.040 212.510 106.180 212.990 ;
        RECT 106.040 212.370 110.780 212.510 ;
        RECT 64.090 211.970 64.410 212.230 ;
        RECT 86.630 211.970 86.950 212.230 ;
        RECT 95.830 212.170 96.150 212.230 ;
        RECT 96.305 212.170 96.595 212.215 ;
        RECT 95.830 212.030 96.595 212.170 ;
        RECT 95.830 211.970 96.150 212.030 ;
        RECT 96.305 211.985 96.595 212.030 ;
        RECT 104.570 211.970 104.890 212.230 ;
        RECT 110.640 212.215 110.780 212.370 ;
        RECT 109.185 212.170 109.475 212.215 ;
        RECT 109.185 212.030 109.860 212.170 ;
        RECT 109.185 211.985 109.475 212.030 ;
        RECT 87.565 211.490 87.855 211.535 ;
        RECT 89.390 211.490 89.710 211.550 ;
        RECT 87.565 211.350 89.710 211.490 ;
        RECT 87.565 211.305 87.855 211.350 ;
        RECT 89.390 211.290 89.710 211.350 ;
        RECT 97.225 211.490 97.515 211.535 ;
        RECT 99.050 211.490 99.370 211.550 ;
        RECT 97.225 211.350 99.370 211.490 ;
        RECT 97.225 211.305 97.515 211.350 ;
        RECT 99.050 211.290 99.370 211.350 ;
        RECT 107.790 211.290 108.110 211.550 ;
        RECT 108.710 211.290 109.030 211.550 ;
        RECT 109.720 211.535 109.860 212.030 ;
        RECT 110.565 211.985 110.855 212.215 ;
        RECT 116.070 212.170 116.390 212.230 ;
        RECT 117.465 212.170 117.755 212.215 ;
        RECT 116.070 212.030 117.755 212.170 ;
        RECT 116.070 211.970 116.390 212.030 ;
        RECT 117.465 211.985 117.755 212.030 ;
        RECT 126.190 212.170 126.510 212.230 ;
        RECT 128.505 212.170 128.795 212.215 ;
        RECT 126.190 212.030 128.795 212.170 ;
        RECT 126.190 211.970 126.510 212.030 ;
        RECT 128.505 211.985 128.795 212.030 ;
        RECT 136.310 212.170 136.630 212.230 ;
        RECT 137.245 212.170 137.535 212.215 ;
        RECT 136.310 212.030 137.535 212.170 ;
        RECT 136.310 211.970 136.630 212.030 ;
        RECT 137.245 211.985 137.535 212.030 ;
        RECT 109.645 211.305 109.935 211.535 ;
        RECT 116.530 211.290 116.850 211.550 ;
        RECT 127.570 211.290 127.890 211.550 ;
        RECT 137.690 211.290 138.010 211.550 ;
        RECT 11.120 210.670 151.295 211.150 ;
        RECT 42.025 210.285 42.315 210.515 ;
        RECT 81.125 210.470 81.415 210.515 ;
        RECT 84.345 210.470 84.635 210.515 ;
        RECT 86.630 210.470 86.950 210.530 ;
        RECT 81.125 210.330 84.100 210.470 ;
        RECT 81.125 210.285 81.415 210.330 ;
        RECT 14.870 210.130 15.190 210.190 ;
        RECT 15.345 210.130 15.635 210.175 ;
        RECT 14.870 209.990 15.635 210.130 ;
        RECT 14.870 209.930 15.190 209.990 ;
        RECT 15.345 209.945 15.635 209.990 ;
        RECT 24.990 210.130 25.310 210.190 ;
        RECT 27.305 210.130 27.595 210.175 ;
        RECT 24.990 209.990 27.595 210.130 ;
        RECT 24.990 209.930 25.310 209.990 ;
        RECT 27.305 209.945 27.595 209.990 ;
        RECT 31.445 210.130 31.735 210.175 ;
        RECT 34.205 210.130 34.495 210.175 ;
        RECT 35.110 210.130 35.430 210.190 ;
        RECT 31.445 209.990 33.040 210.130 ;
        RECT 31.445 209.945 31.735 209.990 ;
        RECT 32.900 209.850 33.040 209.990 ;
        RECT 34.205 209.990 35.430 210.130 ;
        RECT 42.100 210.130 42.240 210.285 ;
        RECT 42.100 209.990 49.600 210.130 ;
        RECT 34.205 209.945 34.495 209.990 ;
        RECT 35.110 209.930 35.430 209.990 ;
        RECT 17.185 209.790 17.475 209.835 ;
        RECT 19.470 209.790 19.790 209.850 ;
        RECT 21.310 209.835 21.630 209.850 ;
        RECT 17.185 209.650 19.790 209.790 ;
        RECT 17.185 209.605 17.475 209.650 ;
        RECT 19.470 209.590 19.790 209.650 ;
        RECT 21.280 209.605 21.630 209.835 ;
        RECT 29.145 209.605 29.435 209.835 ;
        RECT 32.365 209.605 32.655 209.835 ;
        RECT 21.310 209.590 21.630 209.605 ;
        RECT 19.930 209.250 20.250 209.510 ;
        RECT 20.825 209.450 21.115 209.495 ;
        RECT 22.015 209.450 22.305 209.495 ;
        RECT 24.535 209.450 24.825 209.495 ;
        RECT 20.825 209.310 24.825 209.450 ;
        RECT 20.825 209.265 21.115 209.310 ;
        RECT 22.015 209.265 22.305 209.310 ;
        RECT 24.535 209.265 24.825 209.310 ;
        RECT 20.430 209.110 20.720 209.155 ;
        RECT 22.530 209.110 22.820 209.155 ;
        RECT 24.100 209.110 24.390 209.155 ;
        RECT 20.430 208.970 24.390 209.110 ;
        RECT 29.220 209.110 29.360 209.605 ;
        RECT 30.050 209.450 30.370 209.510 ;
        RECT 32.440 209.450 32.580 209.605 ;
        RECT 32.810 209.590 33.130 209.850 ;
        RECT 33.745 209.605 34.035 209.835 ;
        RECT 33.820 209.450 33.960 209.605 ;
        RECT 36.030 209.590 36.350 209.850 ;
        RECT 37.870 209.790 38.190 209.850 ;
        RECT 38.345 209.790 38.635 209.835 ;
        RECT 37.870 209.650 38.635 209.790 ;
        RECT 37.870 209.590 38.190 209.650 ;
        RECT 38.345 209.605 38.635 209.650 ;
        RECT 40.185 209.790 40.475 209.835 ;
        RECT 43.390 209.790 43.710 209.850 ;
        RECT 40.185 209.650 43.710 209.790 ;
        RECT 40.185 209.605 40.475 209.650 ;
        RECT 43.390 209.590 43.710 209.650 ;
        RECT 44.325 209.790 44.615 209.835 ;
        RECT 46.165 209.790 46.455 209.835 ;
        RECT 47.990 209.790 48.310 209.850 ;
        RECT 49.460 209.835 49.600 209.990 ;
        RECT 55.900 209.990 64.320 210.130 ;
        RECT 55.900 209.850 56.040 209.990 ;
        RECT 44.325 209.650 45.920 209.790 ;
        RECT 44.325 209.605 44.615 209.650 ;
        RECT 30.050 209.310 33.960 209.450 ;
        RECT 38.790 209.450 39.110 209.510 ;
        RECT 39.725 209.450 40.015 209.495 ;
        RECT 38.790 209.310 40.015 209.450 ;
        RECT 30.050 209.250 30.370 209.310 ;
        RECT 38.790 209.250 39.110 209.310 ;
        RECT 39.725 209.265 40.015 209.310 ;
        RECT 42.930 209.110 43.250 209.170 ;
        RECT 29.220 208.970 43.250 209.110 ;
        RECT 20.430 208.925 20.720 208.970 ;
        RECT 22.530 208.925 22.820 208.970 ;
        RECT 24.100 208.925 24.390 208.970 ;
        RECT 42.930 208.910 43.250 208.970 ;
        RECT 43.405 209.110 43.695 209.155 ;
        RECT 44.770 209.110 45.090 209.170 ;
        RECT 43.405 208.970 45.090 209.110 ;
        RECT 43.405 208.925 43.695 208.970 ;
        RECT 44.770 208.910 45.090 208.970 ;
        RECT 45.780 208.830 45.920 209.650 ;
        RECT 46.165 209.650 48.310 209.790 ;
        RECT 46.165 209.605 46.455 209.650 ;
        RECT 47.990 209.590 48.310 209.650 ;
        RECT 49.385 209.605 49.675 209.835 ;
        RECT 53.050 209.590 53.370 209.850 ;
        RECT 55.365 209.790 55.655 209.835 ;
        RECT 55.810 209.790 56.130 209.850 ;
        RECT 55.365 209.650 56.130 209.790 ;
        RECT 55.365 209.605 55.655 209.650 ;
        RECT 55.810 209.590 56.130 209.650 ;
        RECT 56.700 209.790 56.990 209.835 ;
        RECT 58.110 209.790 58.430 209.850 ;
        RECT 64.180 209.835 64.320 209.990 ;
        RECT 74.300 209.990 83.180 210.130 ;
        RECT 56.700 209.650 58.430 209.790 ;
        RECT 56.700 209.605 56.990 209.650 ;
        RECT 58.110 209.590 58.430 209.650 ;
        RECT 64.105 209.605 64.395 209.835 ;
        RECT 64.550 209.790 64.870 209.850 ;
        RECT 74.300 209.835 74.440 209.990 ;
        RECT 65.385 209.790 65.675 209.835 ;
        RECT 71.925 209.790 72.215 209.835 ;
        RECT 64.550 209.650 65.675 209.790 ;
        RECT 64.550 209.590 64.870 209.650 ;
        RECT 65.385 209.605 65.675 209.650 ;
        RECT 71.080 209.650 72.215 209.790 ;
        RECT 46.625 209.450 46.915 209.495 ;
        RECT 47.530 209.450 47.850 209.510 ;
        RECT 46.625 209.310 47.850 209.450 ;
        RECT 46.625 209.265 46.915 209.310 ;
        RECT 47.530 209.250 47.850 209.310 ;
        RECT 48.925 209.265 49.215 209.495 ;
        RECT 51.225 209.450 51.515 209.495 ;
        RECT 52.605 209.450 52.895 209.495 ;
        RECT 51.225 209.310 52.895 209.450 ;
        RECT 51.225 209.265 51.515 209.310 ;
        RECT 52.605 209.265 52.895 209.310 ;
        RECT 56.245 209.450 56.535 209.495 ;
        RECT 57.435 209.450 57.725 209.495 ;
        RECT 59.955 209.450 60.245 209.495 ;
        RECT 56.245 209.310 60.245 209.450 ;
        RECT 56.245 209.265 56.535 209.310 ;
        RECT 57.435 209.265 57.725 209.310 ;
        RECT 59.955 209.265 60.245 209.310 ;
        RECT 64.985 209.450 65.275 209.495 ;
        RECT 66.175 209.450 66.465 209.495 ;
        RECT 68.695 209.450 68.985 209.495 ;
        RECT 64.985 209.310 68.985 209.450 ;
        RECT 64.985 209.265 65.275 209.310 ;
        RECT 66.175 209.265 66.465 209.310 ;
        RECT 68.695 209.265 68.985 209.310 ;
        RECT 48.005 209.110 48.295 209.155 ;
        RECT 49.000 209.110 49.140 209.265 ;
        RECT 48.005 208.970 49.140 209.110 ;
        RECT 55.850 209.110 56.140 209.155 ;
        RECT 57.950 209.110 58.240 209.155 ;
        RECT 59.520 209.110 59.810 209.155 ;
        RECT 55.850 208.970 59.810 209.110 ;
        RECT 48.005 208.925 48.295 208.970 ;
        RECT 55.850 208.925 56.140 208.970 ;
        RECT 57.950 208.925 58.240 208.970 ;
        RECT 59.520 208.925 59.810 208.970 ;
        RECT 64.090 208.910 64.410 209.170 ;
        RECT 71.080 209.155 71.220 209.650 ;
        RECT 71.925 209.605 72.215 209.650 ;
        RECT 74.225 209.605 74.515 209.835 ;
        RECT 74.670 209.790 74.990 209.850 ;
        RECT 75.505 209.790 75.795 209.835 ;
        RECT 74.670 209.650 75.795 209.790 ;
        RECT 83.040 209.790 83.180 209.990 ;
        RECT 83.410 209.930 83.730 210.190 ;
        RECT 83.960 210.130 84.100 210.330 ;
        RECT 84.345 210.330 86.950 210.470 ;
        RECT 84.345 210.285 84.635 210.330 ;
        RECT 86.630 210.270 86.950 210.330 ;
        RECT 103.665 210.470 103.955 210.515 ;
        RECT 104.570 210.470 104.890 210.530 ;
        RECT 103.665 210.330 104.890 210.470 ;
        RECT 103.665 210.285 103.955 210.330 ;
        RECT 104.570 210.270 104.890 210.330 ;
        RECT 116.530 210.270 116.850 210.530 ;
        RECT 85.265 210.130 85.555 210.175 ;
        RECT 83.960 209.990 85.555 210.130 ;
        RECT 85.265 209.945 85.555 209.990 ;
        RECT 85.710 210.130 86.030 210.190 ;
        RECT 87.105 210.130 87.395 210.175 ;
        RECT 105.460 210.130 105.750 210.175 ;
        RECT 107.790 210.130 108.110 210.190 ;
        RECT 85.710 209.990 87.395 210.130 ;
        RECT 85.710 209.930 86.030 209.990 ;
        RECT 87.105 209.945 87.395 209.990 ;
        RECT 89.020 209.990 96.980 210.130 ;
        RECT 84.330 209.790 84.650 209.850 ;
        RECT 83.040 209.650 84.650 209.790 ;
        RECT 74.670 209.590 74.990 209.650 ;
        RECT 75.505 209.605 75.795 209.650 ;
        RECT 84.330 209.590 84.650 209.650 ;
        RECT 75.105 209.450 75.395 209.495 ;
        RECT 76.295 209.450 76.585 209.495 ;
        RECT 78.815 209.450 79.105 209.495 ;
        RECT 75.105 209.310 79.105 209.450 ;
        RECT 84.420 209.450 84.560 209.590 ;
        RECT 89.020 209.510 89.160 209.990 ;
        RECT 89.390 209.790 89.710 209.850 ;
        RECT 96.840 209.835 96.980 209.990 ;
        RECT 105.460 209.990 108.110 210.130 ;
        RECT 105.460 209.945 105.750 209.990 ;
        RECT 107.790 209.930 108.110 209.990 ;
        RECT 90.225 209.790 90.515 209.835 ;
        RECT 89.390 209.650 90.515 209.790 ;
        RECT 89.390 209.590 89.710 209.650 ;
        RECT 90.225 209.605 90.515 209.650 ;
        RECT 96.765 209.605 97.055 209.835 ;
        RECT 98.100 209.790 98.390 209.835 ;
        RECT 99.970 209.790 100.290 209.850 ;
        RECT 111.485 209.790 111.775 209.835 ;
        RECT 98.100 209.650 100.290 209.790 ;
        RECT 98.100 209.605 98.390 209.650 ;
        RECT 99.970 209.590 100.290 209.650 ;
        RECT 111.100 209.650 111.775 209.790 ;
        RECT 88.930 209.450 89.250 209.510 ;
        RECT 84.420 209.310 89.250 209.450 ;
        RECT 75.105 209.265 75.395 209.310 ;
        RECT 76.295 209.265 76.585 209.310 ;
        RECT 78.815 209.265 79.105 209.310 ;
        RECT 88.930 209.250 89.250 209.310 ;
        RECT 89.825 209.450 90.115 209.495 ;
        RECT 91.015 209.450 91.305 209.495 ;
        RECT 93.535 209.450 93.825 209.495 ;
        RECT 89.825 209.310 93.825 209.450 ;
        RECT 89.825 209.265 90.115 209.310 ;
        RECT 91.015 209.265 91.305 209.310 ;
        RECT 93.535 209.265 93.825 209.310 ;
        RECT 97.645 209.450 97.935 209.495 ;
        RECT 98.835 209.450 99.125 209.495 ;
        RECT 101.355 209.450 101.645 209.495 ;
        RECT 97.645 209.310 101.645 209.450 ;
        RECT 97.645 209.265 97.935 209.310 ;
        RECT 98.835 209.265 99.125 209.310 ;
        RECT 101.355 209.265 101.645 209.310 ;
        RECT 104.125 209.265 104.415 209.495 ;
        RECT 105.005 209.450 105.295 209.495 ;
        RECT 106.195 209.450 106.485 209.495 ;
        RECT 108.715 209.450 109.005 209.495 ;
        RECT 105.005 209.310 109.005 209.450 ;
        RECT 105.005 209.265 105.295 209.310 ;
        RECT 106.195 209.265 106.485 209.310 ;
        RECT 108.715 209.265 109.005 209.310 ;
        RECT 64.590 209.110 64.880 209.155 ;
        RECT 66.690 209.110 66.980 209.155 ;
        RECT 68.260 209.110 68.550 209.155 ;
        RECT 64.590 208.970 68.550 209.110 ;
        RECT 64.590 208.925 64.880 208.970 ;
        RECT 66.690 208.925 66.980 208.970 ;
        RECT 68.260 208.925 68.550 208.970 ;
        RECT 71.005 208.925 71.295 209.155 ;
        RECT 74.710 209.110 75.000 209.155 ;
        RECT 76.810 209.110 77.100 209.155 ;
        RECT 78.380 209.110 78.670 209.155 ;
        RECT 74.710 208.970 78.670 209.110 ;
        RECT 74.710 208.925 75.000 208.970 ;
        RECT 76.810 208.925 77.100 208.970 ;
        RECT 78.380 208.925 78.670 208.970 ;
        RECT 79.270 209.110 79.590 209.170 ;
        RECT 81.585 209.110 81.875 209.155 ;
        RECT 79.270 208.970 81.875 209.110 ;
        RECT 79.270 208.910 79.590 208.970 ;
        RECT 81.585 208.925 81.875 208.970 ;
        RECT 89.430 209.110 89.720 209.155 ;
        RECT 91.530 209.110 91.820 209.155 ;
        RECT 93.100 209.110 93.390 209.155 ;
        RECT 89.430 208.970 93.390 209.110 ;
        RECT 89.430 208.925 89.720 208.970 ;
        RECT 91.530 208.925 91.820 208.970 ;
        RECT 93.100 208.925 93.390 208.970 ;
        RECT 97.250 209.110 97.540 209.155 ;
        RECT 99.350 209.110 99.640 209.155 ;
        RECT 100.920 209.110 101.210 209.155 ;
        RECT 97.250 208.970 101.210 209.110 ;
        RECT 97.250 208.925 97.540 208.970 ;
        RECT 99.350 208.925 99.640 208.970 ;
        RECT 100.920 208.925 101.210 208.970 ;
        RECT 26.830 208.570 27.150 208.830 ;
        RECT 30.510 208.570 30.830 208.830 ;
        RECT 33.270 208.570 33.590 208.830 ;
        RECT 37.425 208.770 37.715 208.815 ;
        RECT 38.330 208.770 38.650 208.830 ;
        RECT 37.425 208.630 38.650 208.770 ;
        RECT 37.425 208.585 37.715 208.630 ;
        RECT 38.330 208.570 38.650 208.630 ;
        RECT 45.690 208.570 46.010 208.830 ;
        RECT 54.445 208.770 54.735 208.815 ;
        RECT 61.790 208.770 62.110 208.830 ;
        RECT 54.445 208.630 62.110 208.770 ;
        RECT 54.445 208.585 54.735 208.630 ;
        RECT 61.790 208.570 62.110 208.630 ;
        RECT 62.265 208.770 62.555 208.815 ;
        RECT 64.180 208.770 64.320 208.910 ;
        RECT 62.265 208.630 64.320 208.770 ;
        RECT 73.305 208.770 73.595 208.815 ;
        RECT 75.590 208.770 75.910 208.830 ;
        RECT 73.305 208.630 75.910 208.770 ;
        RECT 62.265 208.585 62.555 208.630 ;
        RECT 73.305 208.585 73.595 208.630 ;
        RECT 75.590 208.570 75.910 208.630 ;
        RECT 82.490 208.770 82.810 208.830 ;
        RECT 83.425 208.770 83.715 208.815 ;
        RECT 82.490 208.630 83.715 208.770 ;
        RECT 82.490 208.570 82.810 208.630 ;
        RECT 83.425 208.585 83.715 208.630 ;
        RECT 83.870 208.770 84.190 208.830 ;
        RECT 95.845 208.770 96.135 208.815 ;
        RECT 83.870 208.630 96.135 208.770 ;
        RECT 104.200 208.770 104.340 209.265 ;
        RECT 111.100 209.155 111.240 209.650 ;
        RECT 111.485 209.605 111.775 209.650 ;
        RECT 113.785 209.790 114.075 209.835 ;
        RECT 116.620 209.790 116.760 210.270 ;
        RECT 113.785 209.650 116.760 209.790 ;
        RECT 121.705 209.790 121.995 209.835 ;
        RECT 122.510 209.790 122.830 209.850 ;
        RECT 124.810 209.835 125.130 209.850 ;
        RECT 121.705 209.650 122.830 209.790 ;
        RECT 113.785 209.605 114.075 209.650 ;
        RECT 121.705 209.605 121.995 209.650 ;
        RECT 122.510 209.590 122.830 209.650 ;
        RECT 124.780 209.605 125.130 209.835 ;
        RECT 124.810 209.590 125.130 209.605 ;
        RECT 118.395 209.450 118.685 209.495 ;
        RECT 120.915 209.450 121.205 209.495 ;
        RECT 122.105 209.450 122.395 209.495 ;
        RECT 118.395 209.310 122.395 209.450 ;
        RECT 118.395 209.265 118.685 209.310 ;
        RECT 120.915 209.265 121.205 209.310 ;
        RECT 122.105 209.265 122.395 209.310 ;
        RECT 122.985 209.450 123.275 209.495 ;
        RECT 123.445 209.450 123.735 209.495 ;
        RECT 122.985 209.310 123.735 209.450 ;
        RECT 122.985 209.265 123.275 209.310 ;
        RECT 123.445 209.265 123.735 209.310 ;
        RECT 124.325 209.450 124.615 209.495 ;
        RECT 125.515 209.450 125.805 209.495 ;
        RECT 128.035 209.450 128.325 209.495 ;
        RECT 124.325 209.310 128.325 209.450 ;
        RECT 124.325 209.265 124.615 209.310 ;
        RECT 125.515 209.265 125.805 209.310 ;
        RECT 128.035 209.265 128.325 209.310 ;
        RECT 104.610 209.110 104.900 209.155 ;
        RECT 106.710 209.110 107.000 209.155 ;
        RECT 108.280 209.110 108.570 209.155 ;
        RECT 104.610 208.970 108.570 209.110 ;
        RECT 104.610 208.925 104.900 208.970 ;
        RECT 106.710 208.925 107.000 208.970 ;
        RECT 108.280 208.925 108.570 208.970 ;
        RECT 111.025 208.925 111.315 209.155 ;
        RECT 111.470 209.110 111.790 209.170 ;
        RECT 116.085 209.110 116.375 209.155 ;
        RECT 111.470 208.970 116.375 209.110 ;
        RECT 111.470 208.910 111.790 208.970 ;
        RECT 116.085 208.925 116.375 208.970 ;
        RECT 118.830 209.110 119.120 209.155 ;
        RECT 120.400 209.110 120.690 209.155 ;
        RECT 122.500 209.110 122.790 209.155 ;
        RECT 118.830 208.970 122.790 209.110 ;
        RECT 118.830 208.925 119.120 208.970 ;
        RECT 120.400 208.925 120.690 208.970 ;
        RECT 122.500 208.925 122.790 208.970 ;
        RECT 123.060 208.830 123.200 209.265 ;
        RECT 123.930 209.110 124.220 209.155 ;
        RECT 126.030 209.110 126.320 209.155 ;
        RECT 127.600 209.110 127.890 209.155 ;
        RECT 123.930 208.970 127.890 209.110 ;
        RECT 123.930 208.925 124.220 208.970 ;
        RECT 126.030 208.925 126.320 208.970 ;
        RECT 127.600 208.925 127.890 208.970 ;
        RECT 105.490 208.770 105.810 208.830 ;
        RECT 104.200 208.630 105.810 208.770 ;
        RECT 83.870 208.570 84.190 208.630 ;
        RECT 95.845 208.585 96.135 208.630 ;
        RECT 105.490 208.570 105.810 208.630 ;
        RECT 111.930 208.570 112.250 208.830 ;
        RECT 112.850 208.770 113.170 208.830 ;
        RECT 113.325 208.770 113.615 208.815 ;
        RECT 112.850 208.630 113.615 208.770 ;
        RECT 112.850 208.570 113.170 208.630 ;
        RECT 113.325 208.585 113.615 208.630 ;
        RECT 122.970 208.570 123.290 208.830 ;
        RECT 130.330 208.570 130.650 208.830 ;
        RECT 11.120 207.950 150.500 208.430 ;
        RECT 21.310 207.750 21.630 207.810 ;
        RECT 22.245 207.750 22.535 207.795 ;
        RECT 21.310 207.610 22.535 207.750 ;
        RECT 21.310 207.550 21.630 207.610 ;
        RECT 22.245 207.565 22.535 207.610 ;
        RECT 25.465 207.750 25.755 207.795 ;
        RECT 30.970 207.750 31.290 207.810 ;
        RECT 25.465 207.610 31.290 207.750 ;
        RECT 25.465 207.565 25.755 207.610 ;
        RECT 30.970 207.550 31.290 207.610 ;
        RECT 47.530 207.550 47.850 207.810 ;
        RECT 53.065 207.750 53.355 207.795 ;
        RECT 55.350 207.750 55.670 207.810 ;
        RECT 53.065 207.610 55.670 207.750 ;
        RECT 53.065 207.565 53.355 207.610 ;
        RECT 55.350 207.550 55.670 207.610 ;
        RECT 61.790 207.550 62.110 207.810 ;
        RECT 65.025 207.750 65.315 207.795 ;
        RECT 64.180 207.610 65.315 207.750 ;
        RECT 24.545 207.225 24.835 207.455 ;
        RECT 23.165 206.730 23.455 206.775 ;
        RECT 24.620 206.730 24.760 207.225 ;
        RECT 26.830 207.210 27.150 207.470 ;
        RECT 32.810 207.410 33.130 207.470 ;
        RECT 29.680 207.270 33.130 207.410 ;
        RECT 26.920 207.070 27.060 207.210 ;
        RECT 26.920 206.930 28.900 207.070 ;
        RECT 23.165 206.590 24.760 206.730 ;
        RECT 26.830 206.730 27.150 206.790 ;
        RECT 28.760 206.775 28.900 206.930 ;
        RECT 27.305 206.730 27.595 206.775 ;
        RECT 26.830 206.590 27.595 206.730 ;
        RECT 23.165 206.545 23.455 206.590 ;
        RECT 26.830 206.530 27.150 206.590 ;
        RECT 27.305 206.545 27.595 206.590 ;
        RECT 28.685 206.545 28.975 206.775 ;
        RECT 29.680 206.110 29.820 207.270 ;
        RECT 32.810 207.210 33.130 207.270 ;
        RECT 35.570 207.410 35.860 207.455 ;
        RECT 37.140 207.410 37.430 207.455 ;
        RECT 39.240 207.410 39.530 207.455 ;
        RECT 35.570 207.270 39.530 207.410 ;
        RECT 35.570 207.225 35.860 207.270 ;
        RECT 37.140 207.225 37.430 207.270 ;
        RECT 39.240 207.225 39.530 207.270 ;
        RECT 47.070 207.210 47.390 207.470 ;
        RECT 35.135 207.070 35.425 207.115 ;
        RECT 37.655 207.070 37.945 207.115 ;
        RECT 38.845 207.070 39.135 207.115 ;
        RECT 35.135 206.930 39.135 207.070 ;
        RECT 35.135 206.885 35.425 206.930 ;
        RECT 37.655 206.885 37.945 206.930 ;
        RECT 38.845 206.885 39.135 206.930 ;
        RECT 38.330 206.775 38.650 206.790 ;
        RECT 30.065 206.545 30.355 206.775 ;
        RECT 38.330 206.730 38.680 206.775 ;
        RECT 38.330 206.590 38.845 206.730 ;
        RECT 38.330 206.545 38.680 206.590 ;
        RECT 30.140 206.110 30.280 206.545 ;
        RECT 38.330 206.530 38.650 206.545 ;
        RECT 39.710 206.530 40.030 206.790 ;
        RECT 52.130 206.530 52.450 206.790 ;
        RECT 61.880 206.730 62.020 207.550 ;
        RECT 64.180 207.410 64.320 207.610 ;
        RECT 65.025 207.565 65.315 207.610 ;
        RECT 73.765 207.750 74.055 207.795 ;
        RECT 74.670 207.750 74.990 207.810 ;
        RECT 73.765 207.610 74.990 207.750 ;
        RECT 73.765 207.565 74.055 207.610 ;
        RECT 74.670 207.550 74.990 207.610 ;
        RECT 83.410 207.550 83.730 207.810 ;
        RECT 99.970 207.550 100.290 207.810 ;
        RECT 122.510 207.750 122.830 207.810 ;
        RECT 123.445 207.750 123.735 207.795 ;
        RECT 103.740 207.610 116.760 207.750 ;
        RECT 67.325 207.410 67.615 207.455 ;
        RECT 64.180 207.270 67.615 207.410 ;
        RECT 64.180 207.130 64.320 207.270 ;
        RECT 67.325 207.225 67.615 207.270 ;
        RECT 85.750 207.410 86.040 207.455 ;
        RECT 87.850 207.410 88.140 207.455 ;
        RECT 89.420 207.410 89.710 207.455 ;
        RECT 85.750 207.270 89.710 207.410 ;
        RECT 85.750 207.225 86.040 207.270 ;
        RECT 87.850 207.225 88.140 207.270 ;
        RECT 89.420 207.225 89.710 207.270 ;
        RECT 92.150 207.410 92.470 207.470 ;
        RECT 103.740 207.410 103.880 207.610 ;
        RECT 92.150 207.270 96.060 207.410 ;
        RECT 92.150 207.210 92.470 207.270 ;
        RECT 64.090 206.870 64.410 207.130 ;
        RECT 66.865 206.885 67.155 207.115 ;
        RECT 70.085 207.070 70.375 207.115 ;
        RECT 84.330 207.070 84.650 207.130 ;
        RECT 95.920 207.115 96.060 207.270 ;
        RECT 97.760 207.270 103.880 207.410 ;
        RECT 104.150 207.410 104.440 207.455 ;
        RECT 106.250 207.410 106.540 207.455 ;
        RECT 107.820 207.410 108.110 207.455 ;
        RECT 104.150 207.270 108.110 207.410 ;
        RECT 85.265 207.070 85.555 207.115 ;
        RECT 70.085 206.930 72.140 207.070 ;
        RECT 70.085 206.885 70.375 206.930 ;
        RECT 64.565 206.730 64.855 206.775 ;
        RECT 66.940 206.730 67.080 206.885 ;
        RECT 61.880 206.590 66.160 206.730 ;
        RECT 66.940 206.590 70.300 206.730 ;
        RECT 64.565 206.545 64.855 206.590 ;
        RECT 44.770 206.390 45.090 206.450 ;
        RECT 45.245 206.390 45.535 206.435 ;
        RECT 44.770 206.250 45.535 206.390 ;
        RECT 66.020 206.390 66.160 206.590 ;
        RECT 69.165 206.390 69.455 206.435 ;
        RECT 66.020 206.250 69.455 206.390 ;
        RECT 70.160 206.390 70.300 206.590 ;
        RECT 70.530 206.530 70.850 206.790 ;
        RECT 72.000 206.775 72.140 206.930 ;
        RECT 84.330 206.930 85.555 207.070 ;
        RECT 84.330 206.870 84.650 206.930 ;
        RECT 85.265 206.885 85.555 206.930 ;
        RECT 86.145 207.070 86.435 207.115 ;
        RECT 87.335 207.070 87.625 207.115 ;
        RECT 89.855 207.070 90.145 207.115 ;
        RECT 86.145 206.930 90.145 207.070 ;
        RECT 86.145 206.885 86.435 206.930 ;
        RECT 87.335 206.885 87.625 206.930 ;
        RECT 89.855 206.885 90.145 206.930 ;
        RECT 95.845 206.885 96.135 207.115 ;
        RECT 71.465 206.545 71.755 206.775 ;
        RECT 71.925 206.545 72.215 206.775 ;
        RECT 71.540 206.390 71.680 206.545 ;
        RECT 72.370 206.530 72.690 206.790 ;
        RECT 81.585 206.730 81.875 206.775 ;
        RECT 82.030 206.730 82.350 206.790 ;
        RECT 83.885 206.730 84.175 206.775 ;
        RECT 81.585 206.590 84.175 206.730 ;
        RECT 81.585 206.545 81.875 206.590 ;
        RECT 82.030 206.530 82.350 206.590 ;
        RECT 83.885 206.545 84.175 206.590 ;
        RECT 84.790 206.530 85.110 206.790 ;
        RECT 91.690 206.730 92.010 206.790 ;
        RECT 97.760 206.775 97.900 207.270 ;
        RECT 104.150 207.225 104.440 207.270 ;
        RECT 106.250 207.225 106.540 207.270 ;
        RECT 107.820 207.225 108.110 207.270 ;
        RECT 111.970 207.410 112.260 207.455 ;
        RECT 114.070 207.410 114.360 207.455 ;
        RECT 115.640 207.410 115.930 207.455 ;
        RECT 111.970 207.270 115.930 207.410 ;
        RECT 111.970 207.225 112.260 207.270 ;
        RECT 114.070 207.225 114.360 207.270 ;
        RECT 115.640 207.225 115.930 207.270 ;
        RECT 104.545 207.070 104.835 207.115 ;
        RECT 105.735 207.070 106.025 207.115 ;
        RECT 108.255 207.070 108.545 207.115 ;
        RECT 104.545 206.930 108.545 207.070 ;
        RECT 104.545 206.885 104.835 206.930 ;
        RECT 105.735 206.885 106.025 206.930 ;
        RECT 108.255 206.885 108.545 206.930 ;
        RECT 112.365 207.070 112.655 207.115 ;
        RECT 113.555 207.070 113.845 207.115 ;
        RECT 116.075 207.070 116.365 207.115 ;
        RECT 112.365 206.930 116.365 207.070 ;
        RECT 112.365 206.885 112.655 206.930 ;
        RECT 113.555 206.885 113.845 206.930 ;
        RECT 116.075 206.885 116.365 206.930 ;
        RECT 97.685 206.730 97.975 206.775 ;
        RECT 91.690 206.590 97.975 206.730 ;
        RECT 91.690 206.530 92.010 206.590 ;
        RECT 97.685 206.545 97.975 206.590 ;
        RECT 99.050 206.730 99.370 206.790 ;
        RECT 99.525 206.730 99.815 206.775 ;
        RECT 99.050 206.590 99.815 206.730 ;
        RECT 99.050 206.530 99.370 206.590 ;
        RECT 99.525 206.545 99.815 206.590 ;
        RECT 103.665 206.730 103.955 206.775 ;
        RECT 110.550 206.730 110.870 206.790 ;
        RECT 112.850 206.775 113.170 206.790 ;
        RECT 111.485 206.730 111.775 206.775 ;
        RECT 112.820 206.730 113.170 206.775 ;
        RECT 103.665 206.590 111.775 206.730 ;
        RECT 112.655 206.590 113.170 206.730 ;
        RECT 103.665 206.545 103.955 206.590 ;
        RECT 105.580 206.450 105.720 206.590 ;
        RECT 110.550 206.530 110.870 206.590 ;
        RECT 111.485 206.545 111.775 206.590 ;
        RECT 112.820 206.545 113.170 206.590 ;
        RECT 112.850 206.530 113.170 206.545 ;
        RECT 70.160 206.250 71.680 206.390 ;
        RECT 44.770 206.190 45.090 206.250 ;
        RECT 45.245 206.205 45.535 206.250 ;
        RECT 69.165 206.205 69.455 206.250 ;
        RECT 82.505 206.205 82.795 206.435 ;
        RECT 84.345 206.390 84.635 206.435 ;
        RECT 86.490 206.390 86.780 206.435 ;
        RECT 84.345 206.250 86.780 206.390 ;
        RECT 84.345 206.205 84.635 206.250 ;
        RECT 86.490 206.205 86.780 206.250 ;
        RECT 105.000 206.205 105.290 206.435 ;
        RECT 25.465 206.050 25.755 206.095 ;
        RECT 27.765 206.050 28.055 206.095 ;
        RECT 25.465 205.910 28.055 206.050 ;
        RECT 25.465 205.865 25.755 205.910 ;
        RECT 27.765 205.865 28.055 205.910 ;
        RECT 29.590 205.850 29.910 206.110 ;
        RECT 30.050 205.850 30.370 206.110 ;
        RECT 45.690 206.050 46.010 206.110 ;
        RECT 65.470 206.050 65.790 206.110 ;
        RECT 45.690 205.910 65.790 206.050 ;
        RECT 45.690 205.850 46.010 205.910 ;
        RECT 65.470 205.850 65.790 205.910 ;
        RECT 68.230 205.850 68.550 206.110 ;
        RECT 68.705 206.050 68.995 206.095 ;
        RECT 71.450 206.050 71.770 206.110 ;
        RECT 68.705 205.910 71.770 206.050 ;
        RECT 68.705 205.865 68.995 205.910 ;
        RECT 71.450 205.850 71.770 205.910 ;
        RECT 77.890 206.050 78.210 206.110 ;
        RECT 82.580 206.050 82.720 206.205 ;
        RECT 83.870 206.050 84.190 206.110 ;
        RECT 77.890 205.910 84.190 206.050 ;
        RECT 77.890 205.850 78.210 205.910 ;
        RECT 83.870 205.850 84.190 205.910 ;
        RECT 93.070 205.850 93.390 206.110 ;
        RECT 98.605 206.050 98.895 206.095 ;
        RECT 99.050 206.050 99.370 206.110 ;
        RECT 98.605 205.910 99.370 206.050 ;
        RECT 105.120 206.050 105.260 206.205 ;
        RECT 105.490 206.190 105.810 206.450 ;
        RECT 108.710 206.190 109.030 206.450 ;
        RECT 116.620 206.390 116.760 207.610 ;
        RECT 122.510 207.610 123.735 207.750 ;
        RECT 122.510 207.550 122.830 207.610 ;
        RECT 123.445 207.565 123.735 207.610 ;
        RECT 124.365 207.750 124.655 207.795 ;
        RECT 124.810 207.750 125.130 207.810 ;
        RECT 124.365 207.610 125.130 207.750 ;
        RECT 124.365 207.565 124.655 207.610 ;
        RECT 124.810 207.550 125.130 207.610 ;
        RECT 130.330 207.550 130.650 207.810 ;
        RECT 118.385 207.410 118.675 207.455 ;
        RECT 118.385 207.270 120.440 207.410 ;
        RECT 118.385 207.225 118.675 207.270 ;
        RECT 120.300 207.115 120.440 207.270 ;
        RECT 120.225 206.885 120.515 207.115 ;
        RECT 130.420 207.070 130.560 207.550 ;
        RECT 132.645 207.070 132.935 207.115 ;
        RECT 130.420 206.930 132.935 207.070 ;
        RECT 132.645 206.885 132.935 206.930 ;
        RECT 124.825 206.730 125.115 206.775 ;
        RECT 127.570 206.730 127.890 206.790 ;
        RECT 124.825 206.590 127.890 206.730 ;
        RECT 124.825 206.545 125.115 206.590 ;
        RECT 127.570 206.530 127.890 206.590 ;
        RECT 127.110 206.390 127.430 206.450 ;
        RECT 137.690 206.390 138.010 206.450 ;
        RECT 116.620 206.250 138.010 206.390 ;
        RECT 127.110 206.190 127.430 206.250 ;
        RECT 137.690 206.190 138.010 206.250 ;
        RECT 108.800 206.050 108.940 206.190 ;
        RECT 105.120 205.910 108.940 206.050 ;
        RECT 110.090 206.050 110.410 206.110 ;
        RECT 110.565 206.050 110.855 206.095 ;
        RECT 110.090 205.910 110.855 206.050 ;
        RECT 98.605 205.865 98.895 205.910 ;
        RECT 99.050 205.850 99.370 205.910 ;
        RECT 110.090 205.850 110.410 205.910 ;
        RECT 110.565 205.865 110.855 205.910 ;
        RECT 129.410 206.050 129.730 206.110 ;
        RECT 129.885 206.050 130.175 206.095 ;
        RECT 129.410 205.910 130.175 206.050 ;
        RECT 129.410 205.850 129.730 205.910 ;
        RECT 129.885 205.865 130.175 205.910 ;
        RECT 11.120 205.230 151.295 205.710 ;
        RECT 31.115 205.030 31.405 205.075 ;
        RECT 33.270 205.030 33.590 205.090 ;
        RECT 31.115 204.890 33.590 205.030 ;
        RECT 31.115 204.845 31.405 204.890 ;
        RECT 33.270 204.830 33.590 204.890 ;
        RECT 38.790 204.830 39.110 205.090 ;
        RECT 44.770 205.030 45.090 205.090 ;
        RECT 45.245 205.030 45.535 205.075 ;
        RECT 46.150 205.030 46.470 205.090 ;
        RECT 44.770 204.890 46.470 205.030 ;
        RECT 44.770 204.830 45.090 204.890 ;
        RECT 45.245 204.845 45.535 204.890 ;
        RECT 46.150 204.830 46.470 204.890 ;
        RECT 47.070 205.030 47.390 205.090 ;
        RECT 48.465 205.030 48.755 205.075 ;
        RECT 60.425 205.030 60.715 205.075 ;
        RECT 64.090 205.030 64.410 205.090 ;
        RECT 47.070 204.890 48.755 205.030 ;
        RECT 47.070 204.830 47.390 204.890 ;
        RECT 48.465 204.845 48.755 204.890 ;
        RECT 56.590 204.890 59.260 205.030 ;
        RECT 30.065 204.690 30.355 204.735 ;
        RECT 56.590 204.690 56.730 204.890 ;
        RECT 30.065 204.550 31.200 204.690 ;
        RECT 30.065 204.505 30.355 204.550 ;
        RECT 31.060 204.070 31.200 204.550 ;
        RECT 44.860 204.550 48.680 204.690 ;
        RECT 42.470 204.350 42.790 204.410 ;
        RECT 44.860 204.395 45.000 204.550 ;
        RECT 45.320 204.395 45.920 204.400 ;
        RECT 44.785 204.350 45.075 204.395 ;
        RECT 42.470 204.210 45.075 204.350 ;
        RECT 42.470 204.150 42.790 204.210 ;
        RECT 44.785 204.165 45.075 204.210 ;
        RECT 45.320 204.260 45.995 204.395 ;
        RECT 30.970 203.810 31.290 204.070 ;
        RECT 37.870 203.810 38.190 204.070 ;
        RECT 41.090 203.810 41.410 204.070 ;
        RECT 45.320 204.010 45.460 204.260 ;
        RECT 45.705 204.165 45.995 204.260 ;
        RECT 46.150 204.150 46.470 204.410 ;
        RECT 47.530 204.150 47.850 204.410 ;
        RECT 48.005 204.350 48.295 204.395 ;
        RECT 48.540 204.350 48.680 204.550 ;
        RECT 49.000 204.550 56.730 204.690 ;
        RECT 49.000 204.395 49.140 204.550 ;
        RECT 48.005 204.210 48.680 204.350 ;
        RECT 48.005 204.165 48.295 204.210 ;
        RECT 48.925 204.165 49.215 204.395 ;
        RECT 54.905 204.165 55.195 204.395 ;
        RECT 49.000 204.010 49.140 204.165 ;
        RECT 45.320 203.870 49.140 204.010 ;
        RECT 54.445 203.825 54.735 204.055 ;
        RECT 54.980 204.010 55.120 204.165 ;
        RECT 58.570 204.150 58.890 204.410 ;
        RECT 54.980 203.870 56.500 204.010 ;
        RECT 31.905 203.670 32.195 203.715 ;
        RECT 37.960 203.670 38.100 203.810 ;
        RECT 31.905 203.530 38.100 203.670 ;
        RECT 39.725 203.670 40.015 203.715 ;
        RECT 40.170 203.670 40.490 203.730 ;
        RECT 39.725 203.530 40.490 203.670 ;
        RECT 31.905 203.485 32.195 203.530 ;
        RECT 39.725 203.485 40.015 203.530 ;
        RECT 40.170 203.470 40.490 203.530 ;
        RECT 46.165 203.485 46.455 203.715 ;
        RECT 30.510 203.330 30.830 203.390 ;
        RECT 30.985 203.330 31.275 203.375 ;
        RECT 30.510 203.190 31.275 203.330 ;
        RECT 46.240 203.330 46.380 203.485 ;
        RECT 54.520 203.330 54.660 203.825 ;
        RECT 46.240 203.190 54.660 203.330 ;
        RECT 56.360 203.330 56.500 203.870 ;
        RECT 58.125 203.825 58.415 204.055 ;
        RECT 59.120 204.010 59.260 204.890 ;
        RECT 60.425 204.890 64.410 205.030 ;
        RECT 60.425 204.845 60.715 204.890 ;
        RECT 64.090 204.830 64.410 204.890 ;
        RECT 68.230 205.030 68.550 205.090 ;
        RECT 68.230 204.890 71.220 205.030 ;
        RECT 68.230 204.830 68.550 204.890 ;
        RECT 64.180 204.350 64.320 204.830 ;
        RECT 71.080 204.410 71.220 204.890 ;
        RECT 72.370 204.830 72.690 205.090 ;
        RECT 79.270 204.830 79.590 205.090 ;
        RECT 82.030 204.830 82.350 205.090 ;
        RECT 82.505 205.030 82.795 205.075 ;
        RECT 84.790 205.030 85.110 205.090 ;
        RECT 82.505 204.890 85.110 205.030 ;
        RECT 82.505 204.845 82.795 204.890 ;
        RECT 84.790 204.830 85.110 204.890 ;
        RECT 93.070 204.830 93.390 205.090 ;
        RECT 69.165 204.350 69.455 204.395 ;
        RECT 64.180 204.210 69.455 204.350 ;
        RECT 69.165 204.165 69.455 204.210 ;
        RECT 69.610 204.150 69.930 204.410 ;
        RECT 70.070 204.350 70.390 204.410 ;
        RECT 70.545 204.350 70.835 204.395 ;
        RECT 70.070 204.210 70.835 204.350 ;
        RECT 70.070 204.150 70.390 204.210 ;
        RECT 70.545 204.165 70.835 204.210 ;
        RECT 70.990 204.150 71.310 204.410 ;
        RECT 71.450 204.150 71.770 204.410 ;
        RECT 59.120 203.870 67.540 204.010 ;
        RECT 56.745 203.670 57.035 203.715 ;
        RECT 58.200 203.670 58.340 203.825 ;
        RECT 67.400 203.730 67.540 203.870 ;
        RECT 66.390 203.670 66.710 203.730 ;
        RECT 56.745 203.530 58.340 203.670 ;
        RECT 58.660 203.530 66.710 203.670 ;
        RECT 56.745 203.485 57.035 203.530 ;
        RECT 58.660 203.330 58.800 203.530 ;
        RECT 66.390 203.470 66.710 203.530 ;
        RECT 67.310 203.470 67.630 203.730 ;
        RECT 71.540 203.670 71.680 204.150 ;
        RECT 71.925 204.010 72.215 204.055 ;
        RECT 72.460 204.010 72.600 204.830 ;
        RECT 77.445 204.690 77.735 204.735 ;
        RECT 77.890 204.690 78.210 204.750 ;
        RECT 93.160 204.690 93.300 204.830 ;
        RECT 77.445 204.550 78.210 204.690 ;
        RECT 77.445 204.505 77.735 204.550 ;
        RECT 77.890 204.490 78.210 204.550 ;
        RECT 78.595 204.350 78.885 204.565 ;
        RECT 83.960 204.550 93.300 204.690 ;
        RECT 83.960 204.395 84.100 204.550 ;
        RECT 81.125 204.350 81.415 204.395 ;
        RECT 78.595 204.335 83.640 204.350 ;
        RECT 78.600 204.210 83.640 204.335 ;
        RECT 81.125 204.165 81.415 204.210 ;
        RECT 71.925 203.870 72.600 204.010 ;
        RECT 71.925 203.825 72.215 203.870 ;
        RECT 80.205 203.825 80.495 204.055 ;
        RECT 82.030 204.010 82.350 204.070 ;
        RECT 83.500 204.055 83.640 204.210 ;
        RECT 83.885 204.165 84.175 204.395 ;
        RECT 88.930 204.350 89.250 204.410 ;
        RECT 90.785 204.350 91.075 204.395 ;
        RECT 88.930 204.210 91.075 204.350 ;
        RECT 88.930 204.150 89.250 204.210 ;
        RECT 90.785 204.165 91.075 204.210 ;
        RECT 91.230 204.350 91.550 204.410 ;
        RECT 112.390 204.395 112.710 204.410 ;
        RECT 92.065 204.350 92.355 204.395 ;
        RECT 91.230 204.210 92.355 204.350 ;
        RECT 91.230 204.150 91.550 204.210 ;
        RECT 92.065 204.165 92.355 204.210 ;
        RECT 112.390 204.165 112.740 204.395 ;
        RECT 112.390 204.150 112.710 204.165 ;
        RECT 82.505 204.010 82.795 204.055 ;
        RECT 82.030 203.870 82.795 204.010 ;
        RECT 73.750 203.670 74.070 203.730 ;
        RECT 71.540 203.530 74.070 203.670 ;
        RECT 73.750 203.470 74.070 203.530 ;
        RECT 56.360 203.190 58.800 203.330 ;
        RECT 78.350 203.330 78.670 203.390 ;
        RECT 80.280 203.330 80.420 203.825 ;
        RECT 82.030 203.810 82.350 203.870 ;
        RECT 82.505 203.825 82.795 203.870 ;
        RECT 83.425 204.010 83.715 204.055 ;
        RECT 84.330 204.010 84.650 204.070 ;
        RECT 83.425 203.870 84.650 204.010 ;
        RECT 83.425 203.825 83.715 203.870 ;
        RECT 84.330 203.810 84.650 203.870 ;
        RECT 91.665 204.010 91.955 204.055 ;
        RECT 92.855 204.010 93.145 204.055 ;
        RECT 95.375 204.010 95.665 204.055 ;
        RECT 91.665 203.870 95.665 204.010 ;
        RECT 91.665 203.825 91.955 203.870 ;
        RECT 92.855 203.825 93.145 203.870 ;
        RECT 95.375 203.825 95.665 203.870 ;
        RECT 109.195 204.010 109.485 204.055 ;
        RECT 111.715 204.010 112.005 204.055 ;
        RECT 112.905 204.010 113.195 204.055 ;
        RECT 109.195 203.870 113.195 204.010 ;
        RECT 109.195 203.825 109.485 203.870 ;
        RECT 111.715 203.825 112.005 203.870 ;
        RECT 112.905 203.825 113.195 203.870 ;
        RECT 113.785 203.825 114.075 204.055 ;
        RECT 91.270 203.670 91.560 203.715 ;
        RECT 93.370 203.670 93.660 203.715 ;
        RECT 94.940 203.670 95.230 203.715 ;
        RECT 91.270 203.530 95.230 203.670 ;
        RECT 91.270 203.485 91.560 203.530 ;
        RECT 93.370 203.485 93.660 203.530 ;
        RECT 94.940 203.485 95.230 203.530 ;
        RECT 97.685 203.485 97.975 203.715 ;
        RECT 92.150 203.330 92.470 203.390 ;
        RECT 78.350 203.190 92.470 203.330 ;
        RECT 30.510 203.130 30.830 203.190 ;
        RECT 30.985 203.145 31.275 203.190 ;
        RECT 78.350 203.130 78.670 203.190 ;
        RECT 92.150 203.130 92.470 203.190 ;
        RECT 92.610 203.330 92.930 203.390 ;
        RECT 97.760 203.330 97.900 203.485 ;
        RECT 106.870 203.470 107.190 203.730 ;
        RECT 109.630 203.670 109.920 203.715 ;
        RECT 111.200 203.670 111.490 203.715 ;
        RECT 113.300 203.670 113.590 203.715 ;
        RECT 109.630 203.530 113.590 203.670 ;
        RECT 109.630 203.485 109.920 203.530 ;
        RECT 111.200 203.485 111.490 203.530 ;
        RECT 113.300 203.485 113.590 203.530 ;
        RECT 99.510 203.330 99.830 203.390 ;
        RECT 92.610 203.190 99.830 203.330 ;
        RECT 92.610 203.130 92.930 203.190 ;
        RECT 99.510 203.130 99.830 203.190 ;
        RECT 110.550 203.330 110.870 203.390 ;
        RECT 113.860 203.330 114.000 203.825 ;
        RECT 110.550 203.190 114.000 203.330 ;
        RECT 110.550 203.130 110.870 203.190 ;
        RECT 11.120 202.510 150.500 202.990 ;
        RECT 27.380 202.170 37.180 202.310 ;
        RECT 17.210 201.970 17.500 202.015 ;
        RECT 19.310 201.970 19.600 202.015 ;
        RECT 20.880 201.970 21.170 202.015 ;
        RECT 17.210 201.830 21.170 201.970 ;
        RECT 17.210 201.785 17.500 201.830 ;
        RECT 19.310 201.785 19.600 201.830 ;
        RECT 20.880 201.785 21.170 201.830 ;
        RECT 23.625 201.970 23.915 202.015 ;
        RECT 27.380 201.970 27.520 202.170 ;
        RECT 23.625 201.830 27.520 201.970 ;
        RECT 23.625 201.785 23.915 201.830 ;
        RECT 27.380 201.675 27.520 201.830 ;
        RECT 29.630 201.970 29.920 202.015 ;
        RECT 31.730 201.970 32.020 202.015 ;
        RECT 33.300 201.970 33.590 202.015 ;
        RECT 29.630 201.830 33.590 201.970 ;
        RECT 29.630 201.785 29.920 201.830 ;
        RECT 31.730 201.785 32.020 201.830 ;
        RECT 33.300 201.785 33.590 201.830 ;
        RECT 17.605 201.630 17.895 201.675 ;
        RECT 18.795 201.630 19.085 201.675 ;
        RECT 21.315 201.630 21.605 201.675 ;
        RECT 17.605 201.490 21.605 201.630 ;
        RECT 17.605 201.445 17.895 201.490 ;
        RECT 18.795 201.445 19.085 201.490 ;
        RECT 21.315 201.445 21.605 201.490 ;
        RECT 22.090 201.490 24.300 201.630 ;
        RECT 15.330 201.290 15.650 201.350 ;
        RECT 16.725 201.290 17.015 201.335 ;
        RECT 19.930 201.290 20.250 201.350 ;
        RECT 22.090 201.290 22.230 201.490 ;
        RECT 15.330 201.150 22.230 201.290 ;
        RECT 15.330 201.090 15.650 201.150 ;
        RECT 16.725 201.105 17.015 201.150 ;
        RECT 19.930 201.090 20.250 201.150 ;
        RECT 18.060 200.950 18.350 200.995 ;
        RECT 20.390 200.950 20.710 201.010 ;
        RECT 18.060 200.810 20.710 200.950 ;
        RECT 24.160 200.950 24.300 201.490 ;
        RECT 27.305 201.445 27.595 201.675 ;
        RECT 30.025 201.630 30.315 201.675 ;
        RECT 31.215 201.630 31.505 201.675 ;
        RECT 33.735 201.630 34.025 201.675 ;
        RECT 30.025 201.490 34.025 201.630 ;
        RECT 30.025 201.445 30.315 201.490 ;
        RECT 31.215 201.445 31.505 201.490 ;
        RECT 33.735 201.445 34.025 201.490 ;
        RECT 37.040 201.630 37.180 202.170 ;
        RECT 38.330 202.110 38.650 202.370 ;
        RECT 40.185 202.310 40.475 202.355 ;
        RECT 41.090 202.310 41.410 202.370 ;
        RECT 40.185 202.170 41.410 202.310 ;
        RECT 40.185 202.125 40.475 202.170 ;
        RECT 41.090 202.110 41.410 202.170 ;
        RECT 47.990 202.310 48.310 202.370 ;
        RECT 50.305 202.310 50.595 202.355 ;
        RECT 47.990 202.170 50.595 202.310 ;
        RECT 47.990 202.110 48.310 202.170 ;
        RECT 50.305 202.125 50.595 202.170 ;
        RECT 67.785 202.125 68.075 202.355 ;
        RECT 38.420 201.970 38.560 202.110 ;
        RECT 40.645 201.970 40.935 202.015 ;
        RECT 38.420 201.830 40.935 201.970 ;
        RECT 40.645 201.785 40.935 201.830 ;
        RECT 37.040 201.490 40.400 201.630 ;
        RECT 29.145 201.290 29.435 201.335 ;
        RECT 37.040 201.290 37.180 201.490 ;
        RECT 37.425 201.290 37.715 201.335 ;
        RECT 29.145 201.150 33.040 201.290 ;
        RECT 37.040 201.150 37.715 201.290 ;
        RECT 29.145 201.105 29.435 201.150 ;
        RECT 29.220 200.950 29.360 201.105 ;
        RECT 24.160 200.810 29.360 200.950 ;
        RECT 30.480 200.950 30.770 200.995 ;
        RECT 31.890 200.950 32.210 201.010 ;
        RECT 30.480 200.810 32.210 200.950 ;
        RECT 32.900 200.950 33.040 201.150 ;
        RECT 37.425 201.105 37.715 201.150 ;
        RECT 39.710 201.090 40.030 201.350 ;
        RECT 39.800 200.950 39.940 201.090 ;
        RECT 32.900 200.810 39.940 200.950 ;
        RECT 40.260 200.950 40.400 201.490 ;
        RECT 41.180 201.290 41.320 202.110 ;
        RECT 42.010 201.970 42.330 202.030 ;
        RECT 42.945 201.970 43.235 202.015 ;
        RECT 42.010 201.830 43.235 201.970 ;
        RECT 42.010 201.770 42.330 201.830 ;
        RECT 42.945 201.785 43.235 201.830 ;
        RECT 43.390 201.770 43.710 202.030 ;
        RECT 63.185 201.970 63.475 202.015 ;
        RECT 65.010 201.970 65.330 202.030 ;
        RECT 67.860 201.970 68.000 202.125 ;
        RECT 70.990 202.110 71.310 202.370 ;
        RECT 73.750 202.110 74.070 202.370 ;
        RECT 84.805 202.310 85.095 202.355 ;
        RECT 89.865 202.310 90.155 202.355 ;
        RECT 91.230 202.310 91.550 202.370 ;
        RECT 84.805 202.170 89.620 202.310 ;
        RECT 84.805 202.125 85.095 202.170 ;
        RECT 77.890 201.970 78.210 202.030 ;
        RECT 63.185 201.830 78.210 201.970 ;
        RECT 63.185 201.785 63.475 201.830 ;
        RECT 65.010 201.770 65.330 201.830 ;
        RECT 77.890 201.770 78.210 201.830 ;
        RECT 42.945 201.290 43.235 201.335 ;
        RECT 41.180 201.150 43.235 201.290 ;
        RECT 43.480 201.290 43.620 201.770 ;
        RECT 63.645 201.445 63.935 201.675 ;
        RECT 82.490 201.630 82.810 201.690 ;
        RECT 84.880 201.630 85.020 202.125 ;
        RECT 85.725 201.785 86.015 202.015 ;
        RECT 89.480 201.970 89.620 202.170 ;
        RECT 89.865 202.170 91.550 202.310 ;
        RECT 89.865 202.125 90.155 202.170 ;
        RECT 91.230 202.110 91.550 202.170 ;
        RECT 112.390 202.310 112.710 202.370 ;
        RECT 112.865 202.310 113.155 202.355 ;
        RECT 112.390 202.170 113.155 202.310 ;
        RECT 112.390 202.110 112.710 202.170 ;
        RECT 112.865 202.125 113.155 202.170 ;
        RECT 99.050 201.970 99.370 202.030 ;
        RECT 89.480 201.830 99.370 201.970 ;
        RECT 65.560 201.490 69.380 201.630 ;
        RECT 44.325 201.290 44.615 201.335 ;
        RECT 43.480 201.150 44.615 201.290 ;
        RECT 42.945 201.105 43.235 201.150 ;
        RECT 44.325 201.105 44.615 201.150 ;
        RECT 47.990 201.290 48.310 201.350 ;
        RECT 51.225 201.290 51.515 201.335 ;
        RECT 47.990 201.150 51.515 201.290 ;
        RECT 47.990 201.090 48.310 201.150 ;
        RECT 51.225 201.105 51.515 201.150 ;
        RECT 51.670 201.290 51.990 201.350 ;
        RECT 52.605 201.290 52.895 201.335 ;
        RECT 51.670 201.150 52.895 201.290 ;
        RECT 63.720 201.290 63.860 201.445 ;
        RECT 65.025 201.290 65.315 201.335 ;
        RECT 63.720 201.150 65.315 201.290 ;
        RECT 51.670 201.090 51.990 201.150 ;
        RECT 52.605 201.105 52.895 201.150 ;
        RECT 65.025 201.105 65.315 201.150 ;
        RECT 42.470 200.950 42.790 201.010 ;
        RECT 40.260 200.810 42.790 200.950 ;
        RECT 18.060 200.765 18.350 200.810 ;
        RECT 20.390 200.750 20.710 200.810 ;
        RECT 30.480 200.765 30.770 200.810 ;
        RECT 31.890 200.750 32.210 200.810 ;
        RECT 42.470 200.750 42.790 200.810 ;
        RECT 47.070 200.950 47.390 201.010 ;
        RECT 61.345 200.950 61.635 200.995 ;
        RECT 65.560 200.950 65.700 201.490 ;
        RECT 69.240 201.335 69.380 201.490 ;
        RECT 70.390 201.490 85.020 201.630 ;
        RECT 66.405 201.105 66.695 201.335 ;
        RECT 69.165 201.105 69.455 201.335 ;
        RECT 47.070 200.810 65.700 200.950 ;
        RECT 66.480 200.950 66.620 201.105 ;
        RECT 69.610 201.090 69.930 201.350 ;
        RECT 69.700 200.950 69.840 201.090 ;
        RECT 66.480 200.810 69.840 200.950 ;
        RECT 47.070 200.750 47.390 200.810 ;
        RECT 61.345 200.765 61.635 200.810 ;
        RECT 24.070 200.610 24.390 200.670 ;
        RECT 24.545 200.610 24.835 200.655 ;
        RECT 24.070 200.470 24.835 200.610 ;
        RECT 24.070 200.410 24.390 200.470 ;
        RECT 24.545 200.425 24.835 200.470 ;
        RECT 36.045 200.610 36.335 200.655 ;
        RECT 38.330 200.610 38.650 200.670 ;
        RECT 36.045 200.470 38.650 200.610 ;
        RECT 36.045 200.425 36.335 200.470 ;
        RECT 38.330 200.410 38.650 200.470 ;
        RECT 39.725 200.610 40.015 200.655 ;
        RECT 40.170 200.610 40.490 200.670 ;
        RECT 43.865 200.610 44.155 200.655 ;
        RECT 39.725 200.470 44.155 200.610 ;
        RECT 39.725 200.425 40.015 200.470 ;
        RECT 40.170 200.410 40.490 200.470 ;
        RECT 43.865 200.425 44.155 200.470 ;
        RECT 52.130 200.610 52.450 200.670 ;
        RECT 64.105 200.610 64.395 200.655 ;
        RECT 52.130 200.470 64.395 200.610 ;
        RECT 52.130 200.410 52.450 200.470 ;
        RECT 64.105 200.425 64.395 200.470 ;
        RECT 65.945 200.610 66.235 200.655 ;
        RECT 66.865 200.610 67.155 200.655 ;
        RECT 65.945 200.470 67.155 200.610 ;
        RECT 65.945 200.425 66.235 200.470 ;
        RECT 66.865 200.425 67.155 200.470 ;
        RECT 67.770 200.610 68.090 200.670 ;
        RECT 70.390 200.610 70.530 201.490 ;
        RECT 82.490 201.430 82.810 201.490 ;
        RECT 72.845 201.290 73.135 201.335 ;
        RECT 73.305 201.290 73.595 201.335 ;
        RECT 71.540 201.150 73.595 201.290 ;
        RECT 71.540 201.010 71.680 201.150 ;
        RECT 72.845 201.105 73.135 201.150 ;
        RECT 73.305 201.105 73.595 201.150 ;
        RECT 74.225 201.290 74.515 201.335 ;
        RECT 78.350 201.290 78.670 201.350 ;
        RECT 74.225 201.150 78.670 201.290 ;
        RECT 74.225 201.105 74.515 201.150 ;
        RECT 71.450 200.750 71.770 201.010 ;
        RECT 71.910 200.950 72.230 201.010 ;
        RECT 74.300 200.950 74.440 201.105 ;
        RECT 78.350 201.090 78.670 201.150 ;
        RECT 82.950 201.090 83.270 201.350 ;
        RECT 85.800 201.290 85.940 201.785 ;
        RECT 99.050 201.770 99.370 201.830 ;
        RECT 104.570 201.970 104.860 202.015 ;
        RECT 106.140 201.970 106.430 202.015 ;
        RECT 108.240 201.970 108.530 202.015 ;
        RECT 104.570 201.830 108.530 201.970 ;
        RECT 104.570 201.785 104.860 201.830 ;
        RECT 106.140 201.785 106.430 201.830 ;
        RECT 108.240 201.785 108.530 201.830 ;
        RECT 115.190 201.970 115.480 202.015 ;
        RECT 117.290 201.970 117.580 202.015 ;
        RECT 118.860 201.970 119.150 202.015 ;
        RECT 115.190 201.830 119.150 201.970 ;
        RECT 115.190 201.785 115.480 201.830 ;
        RECT 117.290 201.785 117.580 201.830 ;
        RECT 118.860 201.785 119.150 201.830 ;
        RECT 104.135 201.630 104.425 201.675 ;
        RECT 106.655 201.630 106.945 201.675 ;
        RECT 107.845 201.630 108.135 201.675 ;
        RECT 110.550 201.630 110.870 201.690 ;
        RECT 114.705 201.630 114.995 201.675 ;
        RECT 104.135 201.490 108.135 201.630 ;
        RECT 104.135 201.445 104.425 201.490 ;
        RECT 106.655 201.445 106.945 201.490 ;
        RECT 107.845 201.445 108.135 201.490 ;
        RECT 108.800 201.490 114.995 201.630 ;
        RECT 88.945 201.290 89.235 201.335 ;
        RECT 85.800 201.150 89.235 201.290 ;
        RECT 88.945 201.105 89.235 201.150 ;
        RECT 99.985 201.290 100.275 201.335 ;
        RECT 100.430 201.290 100.750 201.350 ;
        RECT 99.985 201.150 100.750 201.290 ;
        RECT 99.985 201.105 100.275 201.150 ;
        RECT 100.430 201.090 100.750 201.150 ;
        RECT 108.250 201.290 108.570 201.350 ;
        RECT 108.800 201.335 108.940 201.490 ;
        RECT 110.550 201.430 110.870 201.490 ;
        RECT 114.705 201.445 114.995 201.490 ;
        RECT 115.585 201.630 115.875 201.675 ;
        RECT 116.775 201.630 117.065 201.675 ;
        RECT 119.295 201.630 119.585 201.675 ;
        RECT 115.585 201.490 119.585 201.630 ;
        RECT 115.585 201.445 115.875 201.490 ;
        RECT 116.775 201.445 117.065 201.490 ;
        RECT 119.295 201.445 119.585 201.490 ;
        RECT 108.725 201.290 109.015 201.335 ;
        RECT 108.250 201.150 109.015 201.290 ;
        RECT 108.250 201.090 108.570 201.150 ;
        RECT 108.725 201.105 109.015 201.150 ;
        RECT 110.090 201.090 110.410 201.350 ;
        RECT 114.780 201.290 114.920 201.445 ;
        RECT 122.970 201.290 123.290 201.350 ;
        RECT 127.570 201.290 127.890 201.350 ;
        RECT 114.780 201.150 127.890 201.290 ;
        RECT 122.970 201.090 123.290 201.150 ;
        RECT 127.570 201.090 127.890 201.150 ;
        RECT 107.390 200.950 107.680 200.995 ;
        RECT 71.910 200.810 74.440 200.950 ;
        RECT 100.980 200.810 107.680 200.950 ;
        RECT 71.910 200.750 72.230 200.810 ;
        RECT 67.770 200.470 70.530 200.610 ;
        RECT 67.770 200.410 68.090 200.470 ;
        RECT 84.790 200.410 85.110 200.670 ;
        RECT 100.980 200.655 101.120 200.810 ;
        RECT 107.390 200.765 107.680 200.810 ;
        RECT 116.040 200.950 116.330 200.995 ;
        RECT 116.990 200.950 117.310 201.010 ;
        RECT 116.040 200.810 117.310 200.950 ;
        RECT 116.040 200.765 116.330 200.810 ;
        RECT 116.990 200.750 117.310 200.810 ;
        RECT 100.905 200.425 101.195 200.655 ;
        RECT 101.810 200.410 102.130 200.670 ;
        RECT 121.590 200.410 121.910 200.670 ;
        RECT 11.120 199.790 151.295 200.270 ;
        RECT 20.390 199.590 20.710 199.650 ;
        RECT 20.390 199.450 22.230 199.590 ;
        RECT 20.390 199.390 20.710 199.450 ;
        RECT 22.090 198.230 22.230 199.450 ;
        RECT 24.070 199.390 24.390 199.650 ;
        RECT 26.830 199.590 27.150 199.650 ;
        RECT 25.080 199.450 27.150 199.590 ;
        RECT 25.080 199.250 25.220 199.450 ;
        RECT 26.830 199.390 27.150 199.450 ;
        RECT 27.685 199.590 27.975 199.635 ;
        RECT 30.050 199.590 30.370 199.650 ;
        RECT 27.685 199.450 31.660 199.590 ;
        RECT 27.685 199.405 27.975 199.450 ;
        RECT 30.050 199.390 30.370 199.450 ;
        RECT 24.620 199.110 25.220 199.250 ;
        RECT 24.620 198.955 24.760 199.110 ;
        RECT 23.165 198.725 23.455 198.955 ;
        RECT 24.545 198.725 24.835 198.955 ;
        RECT 23.240 198.570 23.380 198.725 ;
        RECT 24.990 198.710 25.310 198.970 ;
        RECT 25.465 198.910 25.755 198.955 ;
        RECT 26.920 198.910 27.060 199.390 ;
        RECT 28.685 199.065 28.975 199.295 ;
        RECT 31.520 199.250 31.660 199.450 ;
        RECT 31.890 199.390 32.210 199.650 ;
        RECT 47.990 199.390 48.310 199.650 ;
        RECT 49.845 199.590 50.135 199.635 ;
        RECT 51.670 199.590 51.990 199.650 ;
        RECT 49.845 199.450 51.990 199.590 ;
        RECT 49.845 199.405 50.135 199.450 ;
        RECT 51.670 199.390 51.990 199.450 ;
        RECT 52.130 199.390 52.450 199.650 ;
        RECT 53.050 199.590 53.370 199.650 ;
        RECT 53.985 199.590 54.275 199.635 ;
        RECT 53.050 199.450 54.275 199.590 ;
        RECT 53.050 199.390 53.370 199.450 ;
        RECT 53.985 199.405 54.275 199.450 ;
        RECT 69.610 199.390 69.930 199.650 ;
        RECT 80.190 199.635 80.510 199.650 ;
        RECT 76.600 199.450 79.960 199.590 ;
        RECT 31.520 199.110 35.800 199.250 ;
        RECT 28.760 198.910 28.900 199.065 ;
        RECT 35.660 198.970 35.800 199.110 ;
        RECT 48.540 199.110 50.060 199.250 ;
        RECT 25.465 198.770 27.060 198.910 ;
        RECT 27.380 198.770 28.900 198.910 ;
        RECT 25.465 198.725 25.755 198.770 ;
        RECT 27.380 198.630 27.520 198.770 ;
        RECT 32.810 198.710 33.130 198.970 ;
        RECT 35.570 198.710 35.890 198.970 ;
        RECT 48.540 198.955 48.680 199.110 ;
        RECT 49.920 198.970 50.060 199.110 ;
        RECT 47.545 198.725 47.835 198.955 ;
        RECT 48.465 198.725 48.755 198.955 ;
        RECT 48.925 198.725 49.215 198.955 ;
        RECT 23.240 198.430 26.140 198.570 ;
        RECT 26.000 198.275 26.140 198.430 ;
        RECT 26.385 198.385 26.675 198.615 ;
        RECT 23.165 198.230 23.455 198.275 ;
        RECT 22.090 198.090 23.455 198.230 ;
        RECT 23.165 198.045 23.455 198.090 ;
        RECT 25.925 198.045 26.215 198.275 ;
        RECT 26.460 198.230 26.600 198.385 ;
        RECT 27.290 198.370 27.610 198.630 ;
        RECT 41.550 198.570 41.870 198.630 ;
        RECT 47.620 198.570 47.760 198.725 ;
        RECT 49.000 198.570 49.140 198.725 ;
        RECT 49.830 198.710 50.150 198.970 ;
        RECT 52.220 198.955 52.360 199.390 ;
        RECT 66.390 199.250 66.710 199.310 ;
        RECT 76.600 199.295 76.740 199.450 ;
        RECT 76.525 199.250 76.815 199.295 ;
        RECT 66.390 199.110 76.815 199.250 ;
        RECT 66.390 199.050 66.710 199.110 ;
        RECT 76.525 199.065 76.815 199.110 ;
        RECT 77.605 199.250 77.895 199.295 ;
        RECT 78.350 199.250 78.670 199.310 ;
        RECT 77.605 199.110 78.670 199.250 ;
        RECT 77.605 199.065 77.895 199.110 ;
        RECT 78.350 199.050 78.670 199.110 ;
        RECT 79.285 199.065 79.575 199.295 ;
        RECT 79.820 199.250 79.960 199.450 ;
        RECT 80.190 199.405 80.575 199.635 ;
        RECT 81.125 199.590 81.415 199.635 ;
        RECT 82.490 199.590 82.810 199.650 ;
        RECT 81.125 199.450 83.180 199.590 ;
        RECT 81.125 199.405 81.415 199.450 ;
        RECT 80.190 199.390 80.510 199.405 ;
        RECT 82.490 199.390 82.810 199.450 ;
        RECT 83.040 199.295 83.180 199.450 ;
        RECT 84.790 199.390 85.110 199.650 ;
        RECT 100.430 199.390 100.750 199.650 ;
        RECT 116.990 199.390 117.310 199.650 ;
        RECT 79.820 199.110 82.720 199.250 ;
        RECT 52.145 198.725 52.435 198.955 ;
        RECT 71.925 198.910 72.215 198.955 ;
        RECT 71.080 198.770 72.215 198.910 ;
        RECT 71.080 198.630 71.220 198.770 ;
        RECT 71.925 198.725 72.215 198.770 ;
        RECT 76.970 198.710 77.290 198.970 ;
        RECT 41.550 198.430 49.140 198.570 ;
        RECT 41.550 198.370 41.870 198.430 ;
        RECT 51.670 198.370 51.990 198.630 ;
        RECT 70.990 198.370 71.310 198.630 ;
        RECT 77.060 198.230 77.200 198.710 ;
        RECT 79.360 198.570 79.500 199.065 ;
        RECT 82.580 198.910 82.720 199.110 ;
        RECT 82.965 199.065 83.255 199.295 ;
        RECT 83.885 199.250 84.175 199.295 ;
        RECT 92.610 199.250 92.930 199.310 ;
        RECT 99.970 199.295 100.290 199.310 ;
        RECT 83.885 199.110 92.930 199.250 ;
        RECT 83.885 199.065 84.175 199.110 ;
        RECT 83.960 198.910 84.100 199.065 ;
        RECT 92.610 199.050 92.930 199.110 ;
        RECT 98.605 199.065 98.895 199.295 ;
        RECT 99.685 199.065 100.290 199.295 ;
        RECT 82.580 198.770 84.100 198.910 ;
        RECT 92.150 198.710 92.470 198.970 ;
        RECT 98.680 198.910 98.820 199.065 ;
        RECT 99.970 199.050 100.290 199.065 ;
        RECT 101.350 199.250 101.670 199.310 ;
        RECT 127.570 199.250 127.890 199.310 ;
        RECT 101.350 199.110 114.920 199.250 ;
        RECT 101.350 199.050 101.670 199.110 ;
        RECT 106.410 198.955 106.730 198.970 ;
        RECT 114.780 198.955 114.920 199.110 ;
        RECT 127.570 199.110 130.100 199.250 ;
        RECT 127.570 199.050 127.890 199.110 ;
        RECT 100.905 198.910 101.195 198.955 ;
        RECT 98.680 198.770 101.195 198.910 ;
        RECT 100.905 198.725 101.195 198.770 ;
        RECT 106.380 198.725 106.730 198.955 ;
        RECT 114.705 198.725 114.995 198.955 ;
        RECT 106.410 198.710 106.730 198.725 ;
        RECT 81.110 198.570 81.430 198.630 ;
        RECT 26.460 198.090 77.200 198.230 ;
        RECT 77.980 198.430 81.430 198.570 ;
        RECT 27.765 197.890 28.055 197.935 ;
        RECT 30.050 197.890 30.370 197.950 ;
        RECT 35.110 197.890 35.430 197.950 ;
        RECT 27.765 197.750 35.430 197.890 ;
        RECT 27.765 197.705 28.055 197.750 ;
        RECT 30.050 197.690 30.370 197.750 ;
        RECT 35.110 197.690 35.430 197.750 ;
        RECT 35.570 197.890 35.890 197.950 ;
        RECT 56.270 197.890 56.590 197.950 ;
        RECT 35.570 197.750 56.590 197.890 ;
        RECT 35.570 197.690 35.890 197.750 ;
        RECT 56.270 197.690 56.590 197.750 ;
        RECT 71.465 197.890 71.755 197.935 ;
        RECT 71.910 197.890 72.230 197.950 ;
        RECT 71.465 197.750 72.230 197.890 ;
        RECT 71.465 197.705 71.755 197.750 ;
        RECT 71.910 197.690 72.230 197.750 ;
        RECT 73.750 197.890 74.070 197.950 ;
        RECT 77.445 197.890 77.735 197.935 ;
        RECT 77.980 197.890 78.120 198.430 ;
        RECT 81.110 198.370 81.430 198.430 ;
        RECT 82.950 198.370 83.270 198.630 ;
        RECT 92.625 198.570 92.915 198.615 ;
        RECT 101.810 198.570 102.130 198.630 ;
        RECT 103.665 198.570 103.955 198.615 ;
        RECT 92.625 198.430 103.955 198.570 ;
        RECT 92.625 198.385 92.915 198.430 ;
        RECT 101.810 198.370 102.130 198.430 ;
        RECT 103.665 198.385 103.955 198.430 ;
        RECT 105.045 198.385 105.335 198.615 ;
        RECT 105.925 198.570 106.215 198.615 ;
        RECT 107.115 198.570 107.405 198.615 ;
        RECT 109.635 198.570 109.925 198.615 ;
        RECT 105.925 198.430 109.925 198.570 ;
        RECT 114.780 198.570 114.920 198.725 ;
        RECT 115.610 198.710 115.930 198.970 ;
        RECT 116.545 198.910 116.835 198.955 ;
        RECT 117.925 198.910 118.215 198.955 ;
        RECT 116.545 198.770 118.215 198.910 ;
        RECT 116.545 198.725 116.835 198.770 ;
        RECT 117.925 198.725 118.215 198.770 ;
        RECT 128.605 198.910 128.895 198.955 ;
        RECT 129.410 198.910 129.730 198.970 ;
        RECT 129.960 198.955 130.100 199.110 ;
        RECT 128.605 198.770 129.730 198.910 ;
        RECT 128.605 198.725 128.895 198.770 ;
        RECT 129.410 198.710 129.730 198.770 ;
        RECT 129.885 198.725 130.175 198.955 ;
        RECT 124.350 198.570 124.670 198.630 ;
        RECT 114.780 198.430 124.670 198.570 ;
        RECT 105.925 198.385 106.215 198.430 ;
        RECT 107.115 198.385 107.405 198.430 ;
        RECT 109.635 198.385 109.925 198.430 ;
        RECT 78.365 198.230 78.655 198.275 ;
        RECT 83.040 198.230 83.180 198.370 ;
        RECT 78.365 198.090 83.180 198.230 ;
        RECT 78.365 198.045 78.655 198.090 ;
        RECT 73.750 197.750 78.120 197.890 ;
        RECT 78.810 197.890 79.130 197.950 ;
        RECT 80.205 197.890 80.495 197.935 ;
        RECT 78.810 197.750 80.495 197.890 ;
        RECT 73.750 197.690 74.070 197.750 ;
        RECT 77.445 197.705 77.735 197.750 ;
        RECT 78.810 197.690 79.130 197.750 ;
        RECT 80.205 197.705 80.495 197.750 ;
        RECT 93.990 197.690 94.310 197.950 ;
        RECT 99.050 197.890 99.370 197.950 ;
        RECT 99.525 197.890 99.815 197.935 ;
        RECT 99.050 197.750 99.815 197.890 ;
        RECT 105.120 197.890 105.260 198.385 ;
        RECT 124.350 198.370 124.670 198.430 ;
        RECT 125.295 198.570 125.585 198.615 ;
        RECT 127.815 198.570 128.105 198.615 ;
        RECT 129.005 198.570 129.295 198.615 ;
        RECT 125.295 198.430 129.295 198.570 ;
        RECT 125.295 198.385 125.585 198.430 ;
        RECT 127.815 198.385 128.105 198.430 ;
        RECT 129.005 198.385 129.295 198.430 ;
        RECT 105.530 198.230 105.820 198.275 ;
        RECT 107.630 198.230 107.920 198.275 ;
        RECT 109.200 198.230 109.490 198.275 ;
        RECT 105.530 198.090 109.490 198.230 ;
        RECT 105.530 198.045 105.820 198.090 ;
        RECT 107.630 198.045 107.920 198.090 ;
        RECT 109.200 198.045 109.490 198.090 ;
        RECT 125.730 198.230 126.020 198.275 ;
        RECT 127.300 198.230 127.590 198.275 ;
        RECT 129.400 198.230 129.690 198.275 ;
        RECT 125.730 198.090 129.690 198.230 ;
        RECT 125.730 198.045 126.020 198.090 ;
        RECT 127.300 198.045 127.590 198.090 ;
        RECT 129.400 198.045 129.690 198.090 ;
        RECT 108.250 197.890 108.570 197.950 ;
        RECT 105.120 197.750 108.570 197.890 ;
        RECT 99.050 197.690 99.370 197.750 ;
        RECT 99.525 197.705 99.815 197.750 ;
        RECT 108.250 197.690 108.570 197.750 ;
        RECT 111.945 197.890 112.235 197.935 ;
        RECT 113.310 197.890 113.630 197.950 ;
        RECT 111.945 197.750 113.630 197.890 ;
        RECT 111.945 197.705 112.235 197.750 ;
        RECT 113.310 197.690 113.630 197.750 ;
        RECT 122.970 197.690 123.290 197.950 ;
        RECT 11.120 197.070 150.500 197.550 ;
        RECT 41.550 196.870 41.870 196.930 ;
        RECT 39.800 196.730 41.870 196.870 ;
        RECT 27.290 196.530 27.610 196.590 ;
        RECT 39.800 196.575 39.940 196.730 ;
        RECT 41.550 196.670 41.870 196.730 ;
        RECT 43.390 196.870 43.710 196.930 ;
        RECT 44.325 196.870 44.615 196.915 ;
        RECT 43.390 196.730 44.615 196.870 ;
        RECT 43.390 196.670 43.710 196.730 ;
        RECT 44.325 196.685 44.615 196.730 ;
        RECT 57.650 196.870 57.970 196.930 ;
        RECT 59.505 196.870 59.795 196.915 ;
        RECT 67.770 196.870 68.090 196.930 ;
        RECT 57.650 196.730 68.090 196.870 ;
        RECT 57.650 196.670 57.970 196.730 ;
        RECT 59.505 196.685 59.795 196.730 ;
        RECT 67.770 196.670 68.090 196.730 ;
        RECT 70.990 196.670 71.310 196.930 ;
        RECT 79.270 196.670 79.590 196.930 ;
        RECT 82.030 196.870 82.350 196.930 ;
        RECT 84.345 196.870 84.635 196.915 ;
        RECT 82.030 196.730 84.635 196.870 ;
        RECT 82.030 196.670 82.350 196.730 ;
        RECT 84.345 196.685 84.635 196.730 ;
        RECT 99.970 196.870 100.290 196.930 ;
        RECT 102.745 196.870 103.035 196.915 ;
        RECT 104.570 196.870 104.890 196.930 ;
        RECT 99.970 196.730 104.890 196.870 ;
        RECT 99.970 196.670 100.290 196.730 ;
        RECT 102.745 196.685 103.035 196.730 ;
        RECT 104.570 196.670 104.890 196.730 ;
        RECT 106.410 196.670 106.730 196.930 ;
        RECT 115.610 196.870 115.930 196.930 ;
        RECT 116.085 196.870 116.375 196.915 ;
        RECT 115.610 196.730 116.375 196.870 ;
        RECT 115.610 196.670 115.930 196.730 ;
        RECT 116.085 196.685 116.375 196.730 ;
        RECT 120.685 196.870 120.975 196.915 ;
        RECT 121.590 196.870 121.910 196.930 ;
        RECT 120.685 196.730 121.910 196.870 ;
        RECT 120.685 196.685 120.975 196.730 ;
        RECT 121.590 196.670 121.910 196.730 ;
        RECT 39.725 196.530 40.015 196.575 ;
        RECT 27.290 196.390 40.015 196.530 ;
        RECT 27.290 196.330 27.610 196.390 ;
        RECT 39.725 196.345 40.015 196.390 ;
        RECT 61.370 196.530 61.660 196.575 ;
        RECT 63.470 196.530 63.760 196.575 ;
        RECT 65.040 196.530 65.330 196.575 ;
        RECT 61.370 196.390 65.330 196.530 ;
        RECT 61.370 196.345 61.660 196.390 ;
        RECT 63.470 196.345 63.760 196.390 ;
        RECT 65.040 196.345 65.330 196.390 ;
        RECT 66.850 196.530 67.170 196.590 ;
        RECT 71.080 196.530 71.220 196.670 ;
        RECT 66.850 196.390 71.220 196.530 ;
        RECT 66.850 196.330 67.170 196.390 ;
        RECT 40.645 196.190 40.935 196.235 ;
        RECT 43.405 196.190 43.695 196.235 ;
        RECT 43.865 196.190 44.155 196.235 ;
        RECT 60.885 196.190 61.175 196.235 ;
        RECT 40.645 196.050 42.700 196.190 ;
        RECT 40.645 196.005 40.935 196.050 ;
        RECT 41.105 195.665 41.395 195.895 ;
        RECT 42.560 195.850 42.700 196.050 ;
        RECT 43.405 196.050 44.155 196.190 ;
        RECT 43.405 196.005 43.695 196.050 ;
        RECT 43.865 196.005 44.155 196.050 ;
        RECT 55.900 196.050 61.175 196.190 ;
        RECT 55.900 195.910 56.040 196.050 ;
        RECT 60.885 196.005 61.175 196.050 ;
        RECT 61.765 196.190 62.055 196.235 ;
        RECT 62.955 196.190 63.245 196.235 ;
        RECT 65.475 196.190 65.765 196.235 ;
        RECT 61.765 196.050 65.765 196.190 ;
        RECT 61.765 196.005 62.055 196.050 ;
        RECT 62.955 196.005 63.245 196.050 ;
        RECT 65.475 196.005 65.765 196.050 ;
        RECT 70.070 195.990 70.390 196.250 ;
        RECT 79.360 196.190 79.500 196.670 ;
        RECT 82.490 196.330 82.810 196.590 ;
        RECT 89.890 196.530 90.180 196.575 ;
        RECT 91.990 196.530 92.280 196.575 ;
        RECT 93.560 196.530 93.850 196.575 ;
        RECT 89.890 196.390 93.850 196.530 ;
        RECT 89.890 196.345 90.180 196.390 ;
        RECT 91.990 196.345 92.280 196.390 ;
        RECT 93.560 196.345 93.850 196.390 ;
        RECT 88.930 196.190 89.250 196.250 ;
        RECT 89.405 196.190 89.695 196.235 ;
        RECT 77.980 196.050 79.500 196.190 ;
        RECT 84.880 196.050 88.700 196.190 ;
        RECT 77.980 195.910 78.120 196.050 ;
        RECT 44.785 195.850 45.075 195.895 ;
        RECT 42.560 195.710 45.075 195.850 ;
        RECT 44.785 195.665 45.075 195.710 ;
        RECT 45.245 195.665 45.535 195.895 ;
        RECT 37.870 195.510 38.190 195.570 ;
        RECT 38.345 195.510 38.635 195.555 ;
        RECT 41.180 195.510 41.320 195.665 ;
        RECT 37.870 195.370 41.320 195.510 ;
        RECT 37.870 195.310 38.190 195.370 ;
        RECT 38.345 195.325 38.635 195.370 ;
        RECT 44.770 195.170 45.090 195.230 ;
        RECT 45.320 195.170 45.460 195.665 ;
        RECT 55.810 195.650 56.130 195.910 ;
        RECT 56.270 195.850 56.590 195.910 ;
        RECT 57.665 195.850 57.955 195.895 ;
        RECT 56.270 195.710 57.955 195.850 ;
        RECT 56.270 195.650 56.590 195.710 ;
        RECT 57.665 195.665 57.955 195.710 ;
        RECT 63.630 195.850 63.950 195.910 ;
        RECT 71.450 195.850 71.770 195.910 ;
        RECT 63.630 195.710 71.770 195.850 ;
        RECT 63.630 195.650 63.950 195.710 ;
        RECT 71.450 195.650 71.770 195.710 ;
        RECT 71.910 195.850 72.230 195.910 ;
        RECT 72.385 195.850 72.675 195.895 ;
        RECT 71.910 195.710 72.675 195.850 ;
        RECT 71.910 195.650 72.230 195.710 ;
        RECT 72.385 195.665 72.675 195.710 ;
        RECT 77.890 195.650 78.210 195.910 ;
        RECT 78.350 195.850 78.670 195.910 ;
        RECT 80.205 195.850 80.495 195.895 ;
        RECT 78.350 195.710 80.495 195.850 ;
        RECT 78.350 195.650 78.670 195.710 ;
        RECT 80.205 195.665 80.495 195.710 ;
        RECT 59.505 195.510 59.795 195.555 ;
        RECT 61.330 195.510 61.650 195.570 ;
        RECT 62.250 195.555 62.570 195.570 ;
        RECT 59.505 195.370 61.650 195.510 ;
        RECT 59.505 195.325 59.795 195.370 ;
        RECT 61.330 195.310 61.650 195.370 ;
        RECT 62.220 195.325 62.570 195.555 ;
        RECT 62.250 195.310 62.570 195.325 ;
        RECT 78.810 195.310 79.130 195.570 ;
        RECT 81.110 195.510 81.430 195.570 ;
        RECT 84.880 195.510 85.020 196.050 ;
        RECT 88.025 195.850 88.315 195.895 ;
        RECT 81.110 195.370 85.020 195.510 ;
        RECT 85.340 195.710 88.315 195.850 ;
        RECT 88.560 195.850 88.700 196.050 ;
        RECT 88.930 196.050 89.695 196.190 ;
        RECT 88.930 195.990 89.250 196.050 ;
        RECT 89.405 196.005 89.695 196.050 ;
        RECT 90.285 196.190 90.575 196.235 ;
        RECT 91.475 196.190 91.765 196.235 ;
        RECT 93.995 196.190 94.285 196.235 ;
        RECT 90.285 196.050 94.285 196.190 ;
        RECT 90.285 196.005 90.575 196.050 ;
        RECT 91.475 196.005 91.765 196.050 ;
        RECT 93.995 196.005 94.285 196.050 ;
        RECT 112.390 196.190 112.710 196.250 ;
        RECT 112.865 196.190 113.155 196.235 ;
        RECT 112.390 196.050 113.155 196.190 ;
        RECT 112.390 195.990 112.710 196.050 ;
        RECT 112.865 196.005 113.155 196.050 ;
        RECT 118.370 196.190 118.690 196.250 ;
        RECT 121.605 196.190 121.895 196.235 ;
        RECT 118.370 196.050 121.895 196.190 ;
        RECT 118.370 195.990 118.690 196.050 ;
        RECT 121.605 196.005 121.895 196.050 ;
        RECT 107.345 195.850 107.635 195.895 ;
        RECT 88.560 195.710 96.520 195.850 ;
        RECT 81.110 195.310 81.430 195.370 ;
        RECT 44.770 195.030 45.460 195.170 ;
        RECT 44.770 194.970 45.090 195.030 ;
        RECT 60.410 194.970 60.730 195.230 ;
        RECT 63.170 195.170 63.490 195.230 ;
        RECT 66.850 195.170 67.170 195.230 ;
        RECT 67.785 195.170 68.075 195.215 ;
        RECT 63.170 195.030 68.075 195.170 ;
        RECT 63.170 194.970 63.490 195.030 ;
        RECT 66.850 194.970 67.170 195.030 ;
        RECT 67.785 194.985 68.075 195.030 ;
        RECT 79.270 195.170 79.590 195.230 ;
        RECT 85.340 195.215 85.480 195.710 ;
        RECT 88.025 195.665 88.315 195.710 ;
        RECT 90.630 195.510 90.920 195.555 ;
        RECT 89.020 195.370 90.920 195.510 ;
        RECT 89.020 195.215 89.160 195.370 ;
        RECT 90.630 195.325 90.920 195.370 ;
        RECT 96.380 195.215 96.520 195.710 ;
        RECT 103.740 195.710 107.635 195.850 ;
        RECT 99.050 195.510 99.370 195.570 ;
        RECT 101.825 195.510 102.115 195.555 ;
        RECT 99.050 195.370 102.115 195.510 ;
        RECT 99.050 195.310 99.370 195.370 ;
        RECT 101.825 195.325 102.115 195.370 ;
        RECT 79.745 195.170 80.035 195.215 ;
        RECT 79.270 195.030 80.035 195.170 ;
        RECT 79.270 194.970 79.590 195.030 ;
        RECT 79.745 194.985 80.035 195.030 ;
        RECT 82.045 195.170 82.335 195.215 ;
        RECT 84.345 195.170 84.635 195.215 ;
        RECT 82.045 195.030 84.635 195.170 ;
        RECT 82.045 194.985 82.335 195.030 ;
        RECT 84.345 194.985 84.635 195.030 ;
        RECT 85.265 194.985 85.555 195.215 ;
        RECT 88.945 194.985 89.235 195.215 ;
        RECT 96.305 195.170 96.595 195.215 ;
        RECT 100.890 195.170 101.210 195.230 ;
        RECT 96.305 195.030 101.210 195.170 ;
        RECT 96.305 194.985 96.595 195.030 ;
        RECT 100.890 194.970 101.210 195.030 ;
        RECT 102.270 195.170 102.590 195.230 ;
        RECT 103.740 195.215 103.880 195.710 ;
        RECT 107.345 195.665 107.635 195.710 ;
        RECT 117.450 195.850 117.770 195.910 ;
        RECT 120.225 195.850 120.515 195.895 ;
        RECT 117.450 195.710 120.515 195.850 ;
        RECT 117.450 195.650 117.770 195.710 ;
        RECT 120.225 195.665 120.515 195.710 ;
        RECT 105.045 195.325 105.335 195.555 ;
        RECT 105.965 195.510 106.255 195.555 ;
        RECT 106.410 195.510 106.730 195.570 ;
        RECT 114.245 195.510 114.535 195.555 ;
        RECT 105.965 195.370 114.535 195.510 ;
        RECT 105.965 195.325 106.255 195.370 ;
        RECT 102.825 195.170 103.115 195.215 ;
        RECT 102.270 195.030 103.115 195.170 ;
        RECT 102.270 194.970 102.590 195.030 ;
        RECT 102.825 194.985 103.115 195.030 ;
        RECT 103.665 194.985 103.955 195.215 ;
        RECT 104.125 195.170 104.415 195.215 ;
        RECT 104.570 195.170 104.890 195.230 ;
        RECT 104.125 195.030 104.890 195.170 ;
        RECT 105.120 195.170 105.260 195.325 ;
        RECT 106.410 195.310 106.730 195.370 ;
        RECT 114.245 195.325 114.535 195.370 ;
        RECT 105.490 195.170 105.810 195.230 ;
        RECT 111.470 195.170 111.790 195.230 ;
        RECT 105.120 195.030 111.790 195.170 ;
        RECT 104.125 194.985 104.415 195.030 ;
        RECT 104.570 194.970 104.890 195.030 ;
        RECT 105.490 194.970 105.810 195.030 ;
        RECT 111.470 194.970 111.790 195.030 ;
        RECT 113.770 194.970 114.090 195.230 ;
        RECT 121.590 194.970 121.910 195.230 ;
        RECT 11.120 194.350 151.295 194.830 ;
        RECT 30.065 194.150 30.355 194.195 ;
        RECT 32.365 194.150 32.655 194.195 ;
        RECT 30.065 194.010 32.655 194.150 ;
        RECT 30.065 193.965 30.355 194.010 ;
        RECT 32.365 193.965 32.655 194.010 ;
        RECT 35.110 194.150 35.430 194.210 ;
        RECT 47.070 194.150 47.390 194.210 ;
        RECT 35.110 194.010 47.390 194.150 ;
        RECT 15.880 193.670 22.230 193.810 ;
        RECT 14.870 193.270 15.190 193.530 ;
        RECT 15.330 193.130 15.650 193.190 ;
        RECT 15.880 193.175 16.020 193.670 ;
        RECT 17.140 193.470 17.430 193.515 ;
        RECT 19.010 193.470 19.330 193.530 ;
        RECT 17.140 193.330 19.330 193.470 ;
        RECT 22.090 193.470 22.230 193.670 ;
        RECT 23.165 193.470 23.455 193.515 ;
        RECT 22.090 193.330 23.455 193.470 ;
        RECT 17.140 193.285 17.430 193.330 ;
        RECT 19.010 193.270 19.330 193.330 ;
        RECT 23.165 193.285 23.455 193.330 ;
        RECT 24.500 193.470 24.790 193.515 ;
        RECT 25.910 193.470 26.230 193.530 ;
        RECT 24.500 193.330 26.230 193.470 ;
        RECT 24.500 193.285 24.790 193.330 ;
        RECT 25.910 193.270 26.230 193.330 ;
        RECT 26.830 193.470 27.150 193.530 ;
        RECT 31.445 193.470 31.735 193.515 ;
        RECT 26.830 193.330 31.735 193.470 ;
        RECT 26.830 193.270 27.150 193.330 ;
        RECT 31.445 193.285 31.735 193.330 ;
        RECT 31.905 193.285 32.195 193.515 ;
        RECT 32.440 193.470 32.580 193.965 ;
        RECT 35.110 193.950 35.430 194.010 ;
        RECT 43.020 193.855 43.160 194.010 ;
        RECT 47.070 193.950 47.390 194.010 ;
        RECT 49.845 194.150 50.135 194.195 ;
        RECT 51.670 194.150 51.990 194.210 ;
        RECT 49.845 194.010 51.990 194.150 ;
        RECT 49.845 193.965 50.135 194.010 ;
        RECT 51.670 193.950 51.990 194.010 ;
        RECT 54.430 194.150 54.750 194.210 ;
        RECT 57.075 194.150 57.365 194.195 ;
        RECT 54.430 194.010 57.365 194.150 ;
        RECT 54.430 193.950 54.750 194.010 ;
        RECT 57.075 193.965 57.365 194.010 ;
        RECT 60.410 193.950 60.730 194.210 ;
        RECT 61.330 193.950 61.650 194.210 ;
        RECT 61.805 194.150 62.095 194.195 ;
        RECT 62.250 194.150 62.570 194.210 ;
        RECT 61.805 194.010 62.570 194.150 ;
        RECT 61.805 193.965 62.095 194.010 ;
        RECT 62.250 193.950 62.570 194.010 ;
        RECT 63.185 193.965 63.475 194.195 ;
        RECT 64.090 194.150 64.410 194.210 ;
        RECT 73.290 194.150 73.610 194.210 ;
        RECT 64.090 194.010 73.610 194.150 ;
        RECT 38.420 193.670 42.240 193.810 ;
        RECT 34.205 193.470 34.495 193.515 ;
        RECT 32.440 193.330 34.495 193.470 ;
        RECT 34.205 193.285 34.495 193.330 ;
        RECT 15.805 193.130 16.095 193.175 ;
        RECT 15.330 192.990 16.095 193.130 ;
        RECT 15.330 192.930 15.650 192.990 ;
        RECT 15.805 192.945 16.095 192.990 ;
        RECT 16.685 193.130 16.975 193.175 ;
        RECT 17.875 193.130 18.165 193.175 ;
        RECT 20.395 193.130 20.685 193.175 ;
        RECT 16.685 192.990 20.685 193.130 ;
        RECT 16.685 192.945 16.975 192.990 ;
        RECT 17.875 192.945 18.165 192.990 ;
        RECT 20.395 192.945 20.685 192.990 ;
        RECT 24.045 193.130 24.335 193.175 ;
        RECT 25.235 193.130 25.525 193.175 ;
        RECT 27.755 193.130 28.045 193.175 ;
        RECT 24.045 192.990 28.045 193.130 ;
        RECT 24.045 192.945 24.335 192.990 ;
        RECT 25.235 192.945 25.525 192.990 ;
        RECT 27.755 192.945 28.045 192.990 ;
        RECT 16.290 192.790 16.580 192.835 ;
        RECT 18.390 192.790 18.680 192.835 ;
        RECT 19.960 192.790 20.250 192.835 ;
        RECT 16.290 192.650 20.250 192.790 ;
        RECT 16.290 192.605 16.580 192.650 ;
        RECT 18.390 192.605 18.680 192.650 ;
        RECT 19.960 192.605 20.250 192.650 ;
        RECT 23.650 192.790 23.940 192.835 ;
        RECT 25.750 192.790 26.040 192.835 ;
        RECT 27.320 192.790 27.610 192.835 ;
        RECT 23.650 192.650 27.610 192.790 ;
        RECT 23.650 192.605 23.940 192.650 ;
        RECT 25.750 192.605 26.040 192.650 ;
        RECT 27.320 192.605 27.610 192.650 ;
        RECT 30.525 192.605 30.815 192.835 ;
        RECT 31.980 192.790 32.120 193.285 ;
        RECT 35.110 193.130 35.430 193.190 ;
        RECT 37.870 193.130 38.190 193.190 ;
        RECT 38.420 193.175 38.560 193.670 ;
        RECT 39.265 193.470 39.555 193.515 ;
        RECT 40.170 193.470 40.490 193.530 ;
        RECT 39.265 193.330 41.780 193.470 ;
        RECT 39.265 193.285 39.555 193.330 ;
        RECT 40.170 193.270 40.490 193.330 ;
        RECT 38.345 193.130 38.635 193.175 ;
        RECT 35.110 192.990 38.635 193.130 ;
        RECT 35.110 192.930 35.430 192.990 ;
        RECT 37.870 192.930 38.190 192.990 ;
        RECT 38.345 192.945 38.635 192.990 ;
        RECT 38.805 192.945 39.095 193.175 ;
        RECT 39.725 193.130 40.015 193.175 ;
        RECT 39.340 192.990 40.015 193.130 ;
        RECT 31.980 192.650 38.560 192.790 ;
        RECT 13.950 192.250 14.270 192.510 ;
        RECT 22.705 192.450 22.995 192.495 ;
        RECT 29.590 192.450 29.910 192.510 ;
        RECT 30.600 192.450 30.740 192.605 ;
        RECT 38.420 192.510 38.560 192.650 ;
        RECT 38.880 192.510 39.020 192.945 ;
        RECT 39.340 192.850 39.480 192.990 ;
        RECT 39.725 192.945 40.015 192.990 ;
        RECT 39.250 192.590 39.570 192.850 ;
        RECT 41.640 192.835 41.780 193.330 ;
        RECT 42.100 193.130 42.240 193.670 ;
        RECT 42.945 193.625 43.235 193.855 ;
        RECT 58.125 193.625 58.415 193.855 ;
        RECT 44.785 193.470 45.075 193.515 ;
        RECT 47.070 193.470 47.390 193.530 ;
        RECT 44.785 193.330 47.390 193.470 ;
        RECT 44.785 193.285 45.075 193.330 ;
        RECT 47.070 193.270 47.390 193.330 ;
        RECT 48.005 193.285 48.295 193.515 ;
        RECT 55.825 193.470 56.115 193.515 ;
        RECT 58.200 193.470 58.340 193.625 ;
        RECT 55.825 193.330 58.340 193.470 ;
        RECT 60.500 193.470 60.640 193.950 ;
        RECT 61.420 193.810 61.560 193.950 ;
        RECT 63.260 193.810 63.400 193.965 ;
        RECT 64.090 193.950 64.410 194.010 ;
        RECT 73.290 193.950 73.610 194.010 ;
        RECT 77.890 193.950 78.210 194.210 ;
        RECT 78.350 194.150 78.670 194.210 ;
        RECT 78.825 194.150 79.115 194.195 ;
        RECT 78.350 194.010 79.115 194.150 ;
        RECT 78.350 193.950 78.670 194.010 ;
        RECT 78.825 193.965 79.115 194.010 ;
        RECT 79.270 194.150 79.590 194.210 ;
        RECT 81.585 194.150 81.875 194.195 ;
        RECT 79.270 194.010 81.875 194.150 ;
        RECT 61.420 193.670 63.400 193.810 ;
        RECT 66.020 193.670 67.080 193.810 ;
        RECT 60.885 193.470 61.175 193.515 ;
        RECT 60.500 193.330 61.175 193.470 ;
        RECT 55.825 193.285 56.115 193.330 ;
        RECT 44.325 193.130 44.615 193.175 ;
        RECT 42.100 192.990 44.615 193.130 ;
        RECT 44.325 192.945 44.615 192.990 ;
        RECT 46.625 193.130 46.915 193.175 ;
        RECT 47.545 193.130 47.835 193.175 ;
        RECT 46.625 192.990 47.835 193.130 ;
        RECT 46.625 192.945 46.915 192.990 ;
        RECT 47.545 192.945 47.835 192.990 ;
        RECT 39.800 192.650 41.320 192.790 ;
        RECT 22.705 192.310 30.740 192.450 ;
        RECT 33.285 192.450 33.575 192.495 ;
        RECT 34.650 192.450 34.970 192.510 ;
        RECT 33.285 192.310 34.970 192.450 ;
        RECT 22.705 192.265 22.995 192.310 ;
        RECT 29.590 192.250 29.910 192.310 ;
        RECT 33.285 192.265 33.575 192.310 ;
        RECT 34.650 192.250 34.970 192.310 ;
        RECT 35.110 192.250 35.430 192.510 ;
        RECT 37.410 192.250 37.730 192.510 ;
        RECT 38.330 192.250 38.650 192.510 ;
        RECT 38.790 192.450 39.110 192.510 ;
        RECT 39.800 192.450 39.940 192.650 ;
        RECT 38.790 192.310 39.940 192.450 ;
        RECT 38.790 192.250 39.110 192.310 ;
        RECT 40.630 192.250 40.950 192.510 ;
        RECT 41.180 192.450 41.320 192.650 ;
        RECT 41.565 192.605 41.855 192.835 ;
        RECT 44.770 192.790 45.090 192.850 ;
        RECT 48.080 192.790 48.220 193.285 ;
        RECT 58.200 193.130 58.340 193.330 ;
        RECT 60.885 193.285 61.175 193.330 ;
        RECT 64.570 193.500 64.860 193.515 ;
        RECT 66.020 193.500 66.160 193.670 ;
        RECT 64.570 193.360 66.160 193.500 ;
        RECT 64.570 193.285 64.860 193.360 ;
        RECT 66.390 193.270 66.710 193.530 ;
        RECT 63.170 193.130 63.490 193.190 ;
        RECT 58.200 192.990 63.490 193.130 ;
        RECT 63.170 192.930 63.490 192.990 ;
        RECT 63.630 192.930 63.950 193.190 ;
        RECT 64.090 192.930 64.410 193.190 ;
        RECT 65.025 192.945 65.315 193.175 ;
        RECT 65.485 192.945 65.775 193.175 ;
        RECT 66.940 193.130 67.080 193.670 ;
        RECT 67.310 193.470 67.630 193.530 ;
        RECT 70.545 193.470 70.835 193.515 ;
        RECT 67.310 193.330 70.835 193.470 ;
        RECT 67.310 193.270 67.630 193.330 ;
        RECT 70.545 193.285 70.835 193.330 ;
        RECT 71.005 193.470 71.295 193.515 ;
        RECT 73.750 193.470 74.070 193.530 ;
        RECT 77.980 193.515 78.120 193.950 ;
        RECT 71.005 193.330 74.070 193.470 ;
        RECT 71.005 193.285 71.295 193.330 ;
        RECT 73.750 193.270 74.070 193.330 ;
        RECT 77.905 193.285 78.195 193.515 ;
        RECT 78.900 193.470 79.040 193.965 ;
        RECT 79.270 193.950 79.590 194.010 ;
        RECT 81.585 193.965 81.875 194.010 ;
        RECT 85.265 193.965 85.555 194.195 ;
        RECT 86.170 194.150 86.490 194.210 ;
        RECT 86.170 194.010 102.040 194.150 ;
        RECT 85.340 193.810 85.480 193.965 ;
        RECT 86.170 193.950 86.490 194.010 ;
        RECT 90.170 193.810 90.460 193.855 ;
        RECT 85.340 193.670 90.460 193.810 ;
        RECT 90.170 193.625 90.460 193.670 ;
        RECT 99.600 193.670 101.580 193.810 ;
        RECT 79.745 193.470 80.035 193.515 ;
        RECT 84.345 193.470 84.635 193.515 ;
        RECT 78.900 193.330 80.035 193.470 ;
        RECT 79.745 193.285 80.035 193.330 ;
        RECT 82.580 193.330 84.635 193.470 ;
        RECT 68.690 193.130 69.010 193.190 ;
        RECT 66.940 192.990 69.010 193.130 ;
        RECT 44.770 192.650 48.220 192.790 ;
        RECT 48.540 192.650 55.580 192.790 ;
        RECT 44.770 192.590 45.090 192.650 ;
        RECT 47.070 192.450 47.390 192.510 ;
        RECT 48.540 192.450 48.680 192.650 ;
        RECT 41.180 192.310 48.680 192.450 ;
        RECT 47.070 192.250 47.390 192.310 ;
        RECT 53.510 192.250 53.830 192.510 ;
        RECT 55.440 192.495 55.580 192.650 ;
        RECT 56.270 192.590 56.590 192.850 ;
        RECT 63.720 192.790 63.860 192.930 ;
        RECT 56.820 192.650 63.860 192.790 ;
        RECT 55.365 192.450 55.655 192.495 ;
        RECT 56.820 192.450 56.960 192.650 ;
        RECT 55.365 192.310 56.960 192.450 ;
        RECT 57.190 192.450 57.510 192.510 ;
        RECT 61.790 192.450 62.110 192.510 ;
        RECT 65.100 192.450 65.240 192.945 ;
        RECT 65.560 192.790 65.700 192.945 ;
        RECT 68.690 192.930 69.010 192.990 ;
        RECT 72.370 193.130 72.690 193.190 ;
        RECT 76.985 193.130 77.275 193.175 ;
        RECT 78.810 193.130 79.130 193.190 ;
        RECT 72.370 192.990 82.260 193.130 ;
        RECT 72.370 192.930 72.690 192.990 ;
        RECT 76.985 192.945 77.275 192.990 ;
        RECT 78.810 192.930 79.130 192.990 ;
        RECT 66.850 192.790 67.170 192.850 ;
        RECT 65.560 192.650 67.170 192.790 ;
        RECT 66.850 192.590 67.170 192.650 ;
        RECT 57.190 192.310 65.240 192.450 ;
        RECT 55.365 192.265 55.655 192.310 ;
        RECT 57.190 192.250 57.510 192.310 ;
        RECT 61.790 192.250 62.110 192.310 ;
        RECT 67.310 192.250 67.630 192.510 ;
        RECT 77.890 192.450 78.210 192.510 ;
        RECT 81.570 192.450 81.890 192.510 ;
        RECT 77.890 192.310 81.890 192.450 ;
        RECT 82.120 192.450 82.260 192.990 ;
        RECT 82.580 192.835 82.720 193.330 ;
        RECT 84.345 193.285 84.635 193.330 ;
        RECT 88.930 193.270 89.250 193.530 ;
        RECT 98.145 193.470 98.435 193.515 ;
        RECT 98.590 193.470 98.910 193.530 ;
        RECT 99.600 193.515 99.740 193.670 ;
        RECT 101.440 193.530 101.580 193.670 ;
        RECT 98.145 193.330 98.910 193.470 ;
        RECT 98.145 193.285 98.435 193.330 ;
        RECT 98.590 193.270 98.910 193.330 ;
        RECT 99.065 193.285 99.355 193.515 ;
        RECT 99.525 193.285 99.815 193.515 ;
        RECT 89.825 193.130 90.115 193.175 ;
        RECT 91.015 193.130 91.305 193.175 ;
        RECT 93.535 193.130 93.825 193.175 ;
        RECT 89.825 192.990 93.825 193.130 ;
        RECT 99.140 193.130 99.280 193.285 ;
        RECT 100.890 193.270 101.210 193.530 ;
        RECT 101.350 193.270 101.670 193.530 ;
        RECT 101.900 193.470 102.040 194.010 ;
        RECT 102.270 193.950 102.590 194.210 ;
        RECT 103.205 194.150 103.495 194.195 ;
        RECT 108.265 194.150 108.555 194.195 ;
        RECT 103.205 194.010 108.555 194.150 ;
        RECT 103.205 193.965 103.495 194.010 ;
        RECT 108.265 193.965 108.555 194.010 ;
        RECT 110.565 194.150 110.855 194.195 ;
        RECT 120.670 194.150 120.990 194.210 ;
        RECT 110.565 194.010 120.990 194.150 ;
        RECT 110.565 193.965 110.855 194.010 ;
        RECT 120.670 193.950 120.990 194.010 ;
        RECT 121.590 193.950 121.910 194.210 ;
        RECT 118.460 193.670 121.360 193.810 ;
        RECT 102.910 193.470 103.200 193.515 ;
        RECT 101.900 193.330 103.200 193.470 ;
        RECT 102.910 193.285 103.200 193.330 ;
        RECT 110.090 193.270 110.410 193.530 ;
        RECT 116.530 193.470 116.850 193.530 ;
        RECT 118.460 193.515 118.600 193.670 ;
        RECT 121.220 193.530 121.360 193.670 ;
        RECT 118.385 193.470 118.675 193.515 ;
        RECT 116.530 193.330 118.675 193.470 ;
        RECT 116.530 193.270 116.850 193.330 ;
        RECT 118.385 193.285 118.675 193.330 ;
        RECT 118.845 193.285 119.135 193.515 ;
        RECT 119.765 193.470 120.055 193.515 ;
        RECT 119.380 193.330 120.055 193.470 ;
        RECT 102.270 193.130 102.590 193.190 ;
        RECT 99.140 192.990 102.590 193.130 ;
        RECT 89.825 192.945 90.115 192.990 ;
        RECT 91.015 192.945 91.305 192.990 ;
        RECT 93.535 192.945 93.825 192.990 ;
        RECT 102.270 192.930 102.590 192.990 ;
        RECT 105.505 193.130 105.795 193.175 ;
        RECT 106.410 193.130 106.730 193.190 ;
        RECT 105.505 192.990 106.730 193.130 ;
        RECT 105.505 192.945 105.795 192.990 ;
        RECT 106.410 192.930 106.730 192.990 ;
        RECT 111.010 192.930 111.330 193.190 ;
        RECT 82.505 192.605 82.795 192.835 ;
        RECT 89.430 192.790 89.720 192.835 ;
        RECT 91.530 192.790 91.820 192.835 ;
        RECT 93.100 192.790 93.390 192.835 ;
        RECT 105.045 192.790 105.335 192.835 ;
        RECT 113.310 192.790 113.630 192.850 ;
        RECT 117.450 192.790 117.770 192.850 ;
        RECT 118.920 192.790 119.060 193.285 ;
        RECT 119.380 193.190 119.520 193.330 ;
        RECT 119.765 193.285 120.055 193.330 ;
        RECT 121.130 193.270 121.450 193.530 ;
        RECT 121.680 193.470 121.820 193.950 ;
        RECT 124.440 193.670 125.500 193.810 ;
        RECT 124.440 193.530 124.580 193.670 ;
        RECT 123.905 193.470 124.195 193.515 ;
        RECT 121.680 193.330 124.195 193.470 ;
        RECT 123.905 193.285 124.195 193.330 ;
        RECT 124.350 193.270 124.670 193.530 ;
        RECT 125.360 193.515 125.500 193.670 ;
        RECT 124.825 193.285 125.115 193.515 ;
        RECT 125.285 193.285 125.575 193.515 ;
        RECT 119.290 193.130 119.610 193.190 ;
        RECT 121.605 193.130 121.895 193.175 ;
        RECT 119.290 192.990 121.895 193.130 ;
        RECT 119.290 192.930 119.610 192.990 ;
        RECT 121.605 192.945 121.895 192.990 ;
        RECT 122.985 192.790 123.275 192.835 ;
        RECT 123.890 192.790 124.210 192.850 ;
        RECT 124.900 192.790 125.040 193.285 ;
        RECT 126.190 193.270 126.510 193.530 ;
        RECT 128.920 193.470 129.210 193.515 ;
        RECT 130.790 193.470 131.110 193.530 ;
        RECT 128.920 193.330 131.110 193.470 ;
        RECT 128.920 193.285 129.210 193.330 ;
        RECT 130.790 193.270 131.110 193.330 ;
        RECT 127.570 192.930 127.890 193.190 ;
        RECT 128.465 193.130 128.755 193.175 ;
        RECT 129.655 193.130 129.945 193.175 ;
        RECT 132.175 193.130 132.465 193.175 ;
        RECT 128.465 192.990 132.465 193.130 ;
        RECT 128.465 192.945 128.755 192.990 ;
        RECT 129.655 192.945 129.945 192.990 ;
        RECT 132.175 192.945 132.465 192.990 ;
        RECT 89.430 192.650 93.390 192.790 ;
        RECT 89.430 192.605 89.720 192.650 ;
        RECT 91.530 192.605 91.820 192.650 ;
        RECT 93.100 192.605 93.390 192.650 ;
        RECT 96.840 192.650 121.360 192.790 ;
        RECT 96.840 192.510 96.980 192.650 ;
        RECT 105.045 192.605 105.335 192.650 ;
        RECT 113.310 192.590 113.630 192.650 ;
        RECT 117.450 192.590 117.770 192.650 ;
        RECT 93.530 192.450 93.850 192.510 ;
        RECT 95.845 192.450 96.135 192.495 ;
        RECT 82.120 192.310 96.135 192.450 ;
        RECT 77.890 192.250 78.210 192.310 ;
        RECT 81.570 192.250 81.890 192.310 ;
        RECT 93.530 192.250 93.850 192.310 ;
        RECT 95.845 192.265 96.135 192.310 ;
        RECT 96.750 192.250 97.070 192.510 ;
        RECT 99.970 192.250 100.290 192.510 ;
        RECT 100.430 192.250 100.750 192.510 ;
        RECT 120.670 192.250 120.990 192.510 ;
        RECT 121.220 192.495 121.360 192.650 ;
        RECT 122.985 192.650 125.040 192.790 ;
        RECT 128.070 192.790 128.360 192.835 ;
        RECT 130.170 192.790 130.460 192.835 ;
        RECT 131.740 192.790 132.030 192.835 ;
        RECT 128.070 192.650 132.030 192.790 ;
        RECT 122.985 192.605 123.275 192.650 ;
        RECT 123.890 192.590 124.210 192.650 ;
        RECT 128.070 192.605 128.360 192.650 ;
        RECT 130.170 192.605 130.460 192.650 ;
        RECT 131.740 192.605 132.030 192.650 ;
        RECT 121.145 192.265 121.435 192.495 ;
        RECT 124.350 192.250 124.670 192.510 ;
        RECT 127.125 192.450 127.415 192.495 ;
        RECT 129.410 192.450 129.730 192.510 ;
        RECT 127.125 192.310 129.730 192.450 ;
        RECT 127.125 192.265 127.415 192.310 ;
        RECT 129.410 192.250 129.730 192.310 ;
        RECT 131.250 192.450 131.570 192.510 ;
        RECT 134.485 192.450 134.775 192.495 ;
        RECT 131.250 192.310 134.775 192.450 ;
        RECT 131.250 192.250 131.570 192.310 ;
        RECT 134.485 192.265 134.775 192.310 ;
        RECT 11.120 191.630 150.500 192.110 ;
        RECT 19.010 191.430 19.330 191.490 ;
        RECT 21.785 191.430 22.075 191.475 ;
        RECT 19.010 191.290 22.075 191.430 ;
        RECT 19.010 191.230 19.330 191.290 ;
        RECT 21.785 191.245 22.075 191.290 ;
        RECT 26.830 191.230 27.150 191.490 ;
        RECT 29.590 191.230 29.910 191.490 ;
        RECT 32.365 191.430 32.655 191.475 ;
        RECT 32.810 191.430 33.130 191.490 ;
        RECT 32.365 191.290 33.130 191.430 ;
        RECT 32.365 191.245 32.655 191.290 ;
        RECT 32.810 191.230 33.130 191.290 ;
        RECT 33.285 191.430 33.575 191.475 ;
        RECT 37.410 191.430 37.730 191.490 ;
        RECT 33.285 191.290 37.730 191.430 ;
        RECT 33.285 191.245 33.575 191.290 ;
        RECT 37.410 191.230 37.730 191.290 ;
        RECT 38.790 191.230 39.110 191.490 ;
        RECT 40.645 191.430 40.935 191.475 ;
        RECT 44.770 191.430 45.090 191.490 ;
        RECT 40.645 191.290 45.090 191.430 ;
        RECT 40.645 191.245 40.935 191.290 ;
        RECT 44.770 191.230 45.090 191.290 ;
        RECT 53.510 191.230 53.830 191.490 ;
        RECT 53.970 191.430 54.290 191.490 ;
        RECT 65.930 191.430 66.250 191.490 ;
        RECT 53.970 191.290 66.250 191.430 ;
        RECT 53.970 191.230 54.290 191.290 ;
        RECT 65.930 191.230 66.250 191.290 ;
        RECT 71.910 191.430 72.230 191.490 ;
        RECT 78.810 191.430 79.130 191.490 ;
        RECT 71.910 191.290 79.130 191.430 ;
        RECT 71.910 191.230 72.230 191.290 ;
        RECT 78.810 191.230 79.130 191.290 ;
        RECT 86.630 191.430 86.950 191.490 ;
        RECT 88.930 191.430 89.250 191.490 ;
        RECT 86.630 191.290 89.250 191.430 ;
        RECT 86.630 191.230 86.950 191.290 ;
        RECT 88.930 191.230 89.250 191.290 ;
        RECT 108.250 191.230 108.570 191.490 ;
        RECT 111.010 191.230 111.330 191.490 ;
        RECT 126.190 191.430 126.510 191.490 ;
        RECT 127.585 191.430 127.875 191.475 ;
        RECT 126.190 191.290 127.875 191.430 ;
        RECT 126.190 191.230 126.510 191.290 ;
        RECT 127.585 191.245 127.875 191.290 ;
        RECT 129.410 191.230 129.730 191.490 ;
        RECT 130.790 191.230 131.110 191.490 ;
        RECT 13.070 191.090 13.360 191.135 ;
        RECT 15.170 191.090 15.460 191.135 ;
        RECT 16.740 191.090 17.030 191.135 ;
        RECT 13.070 190.950 17.030 191.090 ;
        RECT 13.070 190.905 13.360 190.950 ;
        RECT 15.170 190.905 15.460 190.950 ;
        RECT 16.740 190.905 17.030 190.950 ;
        RECT 19.485 190.905 19.775 191.135 ;
        RECT 13.465 190.750 13.755 190.795 ;
        RECT 14.655 190.750 14.945 190.795 ;
        RECT 17.175 190.750 17.465 190.795 ;
        RECT 13.465 190.610 17.465 190.750 ;
        RECT 19.560 190.750 19.700 190.905 ;
        RECT 26.920 190.750 27.060 191.230 ;
        RECT 29.680 190.750 29.820 191.230 ;
        RECT 38.880 190.750 39.020 191.230 ;
        RECT 53.600 190.750 53.740 191.230 ;
        RECT 54.430 191.090 54.750 191.150 ;
        RECT 86.170 191.090 86.490 191.150 ;
        RECT 54.430 190.950 86.490 191.090 ;
        RECT 54.430 190.890 54.750 190.950 ;
        RECT 86.170 190.890 86.490 190.950 ;
        RECT 92.150 191.090 92.470 191.150 ;
        RECT 96.750 191.090 97.070 191.150 ;
        RECT 92.150 190.950 97.440 191.090 ;
        RECT 92.150 190.890 92.470 190.950 ;
        RECT 96.750 190.890 97.070 190.950 ;
        RECT 57.190 190.750 57.510 190.810 ;
        RECT 19.560 190.610 27.060 190.750 ;
        RECT 28.760 190.610 29.820 190.750 ;
        RECT 30.140 190.610 39.020 190.750 ;
        RECT 39.340 190.610 53.740 190.750 ;
        RECT 54.060 190.610 57.510 190.750 ;
        RECT 13.465 190.565 13.755 190.610 ;
        RECT 14.655 190.565 14.945 190.610 ;
        RECT 17.175 190.565 17.465 190.610 ;
        RECT 12.585 190.410 12.875 190.455 ;
        RECT 15.330 190.410 15.650 190.470 ;
        RECT 21.400 190.455 21.540 190.610 ;
        RECT 12.585 190.270 15.650 190.410 ;
        RECT 12.585 190.225 12.875 190.270 ;
        RECT 13.950 190.115 14.270 190.130 ;
        RECT 13.920 190.070 14.270 190.115 ;
        RECT 13.755 189.930 14.270 190.070 ;
        RECT 13.920 189.885 14.270 189.930 ;
        RECT 13.950 189.870 14.270 189.885 ;
        RECT 14.500 189.790 14.640 190.270 ;
        RECT 15.330 190.210 15.650 190.270 ;
        RECT 21.325 190.410 21.615 190.455 ;
        RECT 21.325 190.270 21.725 190.410 ;
        RECT 21.325 190.225 21.615 190.270 ;
        RECT 22.690 190.210 23.010 190.470 ;
        RECT 28.760 190.455 28.900 190.610 ;
        RECT 28.685 190.225 28.975 190.455 ;
        RECT 29.145 190.410 29.435 190.455 ;
        RECT 29.590 190.410 29.910 190.470 ;
        RECT 29.145 190.270 29.910 190.410 ;
        RECT 29.145 190.225 29.435 190.270 ;
        RECT 29.590 190.210 29.910 190.270 ;
        RECT 26.830 190.070 27.150 190.130 ;
        RECT 30.140 190.070 30.280 190.610 ;
        RECT 34.650 190.410 34.970 190.470 ;
        RECT 39.340 190.455 39.480 190.610 ;
        RECT 35.125 190.410 35.415 190.455 ;
        RECT 34.650 190.270 35.415 190.410 ;
        RECT 34.650 190.210 34.970 190.270 ;
        RECT 35.125 190.225 35.415 190.270 ;
        RECT 39.265 190.225 39.555 190.455 ;
        RECT 40.630 190.210 40.950 190.470 ;
        RECT 53.510 190.410 53.830 190.470 ;
        RECT 54.060 190.455 54.200 190.610 ;
        RECT 57.190 190.550 57.510 190.610 ;
        RECT 73.290 190.750 73.610 190.810 ;
        RECT 77.430 190.750 77.750 190.810 ;
        RECT 73.290 190.610 78.580 190.750 ;
        RECT 73.290 190.550 73.610 190.610 ;
        RECT 77.430 190.550 77.750 190.610 ;
        RECT 53.985 190.410 54.275 190.455 ;
        RECT 53.510 190.270 54.275 190.410 ;
        RECT 53.510 190.210 53.830 190.270 ;
        RECT 53.985 190.225 54.275 190.270 ;
        RECT 54.430 190.410 54.750 190.470 ;
        RECT 54.905 190.410 55.195 190.455 ;
        RECT 54.430 190.270 55.195 190.410 ;
        RECT 54.430 190.210 54.750 190.270 ;
        RECT 54.905 190.225 55.195 190.270 ;
        RECT 55.350 190.210 55.670 190.470 ;
        RECT 70.085 190.410 70.375 190.455 ;
        RECT 71.045 190.410 71.335 190.465 ;
        RECT 73.750 190.410 74.070 190.470 ;
        RECT 78.440 190.455 78.580 190.610 ;
        RECT 93.160 190.610 96.525 190.750 ;
        RECT 70.085 190.270 70.485 190.410 ;
        RECT 71.045 190.270 74.070 190.410 ;
        RECT 70.085 190.225 70.375 190.270 ;
        RECT 71.045 190.235 71.335 190.270 ;
        RECT 39.725 190.070 40.015 190.115 ;
        RECT 26.830 189.930 30.280 190.070 ;
        RECT 31.520 189.930 40.015 190.070 ;
        RECT 26.830 189.870 27.150 189.930 ;
        RECT 14.410 189.530 14.730 189.790 ;
        RECT 20.390 189.530 20.710 189.790 ;
        RECT 26.370 189.730 26.690 189.790 ;
        RECT 31.520 189.775 31.660 189.930 ;
        RECT 39.725 189.885 40.015 189.930 ;
        RECT 47.530 190.070 47.850 190.130 ;
        RECT 70.160 190.070 70.300 190.225 ;
        RECT 73.750 190.210 74.070 190.270 ;
        RECT 78.365 190.225 78.655 190.455 ;
        RECT 72.370 190.070 72.690 190.130 ;
        RECT 47.530 189.930 72.690 190.070 ;
        RECT 47.530 189.870 47.850 189.930 ;
        RECT 72.370 189.870 72.690 189.930 ;
        RECT 73.290 190.070 73.610 190.130 ;
        RECT 92.610 190.070 92.930 190.130 ;
        RECT 93.160 190.070 93.300 190.610 ;
        RECT 93.990 190.410 94.310 190.470 ;
        RECT 96.385 190.455 96.525 190.610 ;
        RECT 97.300 190.455 97.440 190.950 ;
        RECT 120.300 190.950 129.180 191.090 ;
        RECT 102.270 190.750 102.590 190.810 ;
        RECT 112.390 190.750 112.710 190.810 ;
        RECT 116.530 190.750 116.850 190.810 ;
        RECT 120.300 190.750 120.440 190.950 ;
        RECT 102.270 190.610 116.850 190.750 ;
        RECT 102.270 190.550 102.590 190.610 ;
        RECT 112.390 190.550 112.710 190.610 ;
        RECT 116.530 190.550 116.850 190.610 ;
        RECT 119.380 190.610 120.440 190.750 ;
        RECT 120.670 190.750 120.990 190.810 ;
        RECT 120.670 190.610 121.360 190.750 ;
        RECT 95.845 190.410 96.135 190.455 ;
        RECT 93.990 190.270 96.135 190.410 ;
        RECT 93.990 190.210 94.310 190.270 ;
        RECT 95.845 190.225 96.135 190.270 ;
        RECT 96.310 190.225 96.600 190.455 ;
        RECT 97.225 190.225 97.515 190.455 ;
        RECT 98.375 190.410 98.665 190.455 ;
        RECT 103.190 190.410 103.510 190.470 ;
        RECT 98.375 190.270 103.510 190.410 ;
        RECT 98.375 190.225 98.665 190.270 ;
        RECT 103.190 190.210 103.510 190.270 ;
        RECT 112.865 190.410 113.155 190.455 ;
        RECT 113.310 190.410 113.630 190.470 ;
        RECT 117.465 190.410 117.755 190.455 ;
        RECT 112.865 190.270 117.755 190.410 ;
        RECT 112.865 190.225 113.155 190.270 ;
        RECT 113.310 190.210 113.630 190.270 ;
        RECT 117.465 190.225 117.755 190.270 ;
        RECT 117.910 190.410 118.230 190.470 ;
        RECT 119.380 190.455 119.520 190.610 ;
        RECT 120.670 190.550 120.990 190.610 ;
        RECT 117.910 190.270 118.830 190.410 ;
        RECT 117.910 190.210 118.230 190.270 ;
        RECT 73.290 189.930 93.300 190.070 ;
        RECT 73.290 189.870 73.610 189.930 ;
        RECT 92.610 189.870 92.930 189.930 ;
        RECT 95.370 189.870 95.690 190.130 ;
        RECT 97.670 189.870 97.990 190.130 ;
        RECT 101.825 190.070 102.115 190.115 ;
        RECT 98.220 189.930 102.115 190.070 ;
        RECT 118.690 190.070 118.830 190.270 ;
        RECT 119.305 190.225 119.595 190.455 ;
        RECT 119.380 190.070 119.520 190.225 ;
        RECT 120.210 190.210 120.530 190.470 ;
        RECT 121.220 190.455 121.360 190.610 ;
        RECT 121.145 190.225 121.435 190.455 ;
        RECT 122.985 190.410 123.275 190.455 ;
        RECT 124.350 190.410 124.670 190.470 ;
        RECT 122.985 190.270 124.670 190.410 ;
        RECT 122.985 190.225 123.275 190.270 ;
        RECT 124.350 190.210 124.670 190.270 ;
        RECT 125.270 190.410 125.590 190.470 ;
        RECT 129.040 190.455 129.180 190.950 ;
        RECT 129.500 190.750 129.640 191.230 ;
        RECT 129.500 190.610 131.940 190.750 ;
        RECT 128.505 190.410 128.795 190.455 ;
        RECT 125.270 190.270 128.795 190.410 ;
        RECT 125.270 190.210 125.590 190.270 ;
        RECT 128.505 190.225 128.795 190.270 ;
        RECT 128.965 190.410 129.255 190.455 ;
        RECT 128.965 190.270 130.100 190.410 ;
        RECT 128.965 190.225 129.255 190.270 ;
        RECT 122.065 190.070 122.355 190.115 ;
        RECT 118.690 189.930 119.520 190.070 ;
        RECT 121.220 189.930 122.355 190.070 ;
        RECT 27.765 189.730 28.055 189.775 ;
        RECT 26.370 189.590 28.055 189.730 ;
        RECT 26.370 189.530 26.690 189.590 ;
        RECT 27.765 189.545 28.055 189.590 ;
        RECT 31.445 189.545 31.735 189.775 ;
        RECT 33.285 189.730 33.575 189.775 ;
        RECT 52.590 189.730 52.910 189.790 ;
        RECT 33.285 189.590 52.910 189.730 ;
        RECT 33.285 189.545 33.575 189.590 ;
        RECT 52.590 189.530 52.910 189.590 ;
        RECT 53.050 189.530 53.370 189.790 ;
        RECT 56.285 189.730 56.575 189.775 ;
        RECT 56.730 189.730 57.050 189.790 ;
        RECT 56.285 189.590 57.050 189.730 ;
        RECT 56.285 189.545 56.575 189.590 ;
        RECT 56.730 189.530 57.050 189.590 ;
        RECT 66.390 189.730 66.710 189.790 ;
        RECT 69.610 189.730 69.930 189.790 ;
        RECT 66.390 189.590 69.930 189.730 ;
        RECT 66.390 189.530 66.710 189.590 ;
        RECT 69.610 189.530 69.930 189.590 ;
        RECT 70.990 189.730 71.310 189.790 ;
        RECT 76.510 189.730 76.830 189.790 ;
        RECT 70.990 189.590 76.830 189.730 ;
        RECT 70.990 189.530 71.310 189.590 ;
        RECT 76.510 189.530 76.830 189.590 ;
        RECT 79.270 189.530 79.590 189.790 ;
        RECT 95.460 189.730 95.600 189.870 ;
        RECT 98.220 189.730 98.360 189.930 ;
        RECT 101.825 189.885 102.115 189.930 ;
        RECT 121.220 189.790 121.360 189.930 ;
        RECT 122.065 189.885 122.355 189.930 ;
        RECT 122.525 189.885 122.815 190.115 ;
        RECT 123.980 189.930 128.720 190.070 ;
        RECT 95.460 189.590 98.360 189.730 ;
        RECT 99.050 189.530 99.370 189.790 ;
        RECT 120.685 189.730 120.975 189.775 ;
        RECT 121.130 189.730 121.450 189.790 ;
        RECT 120.685 189.590 121.450 189.730 ;
        RECT 120.685 189.545 120.975 189.590 ;
        RECT 121.130 189.530 121.450 189.590 ;
        RECT 121.590 189.730 121.910 189.790 ;
        RECT 122.600 189.730 122.740 189.885 ;
        RECT 123.980 189.775 124.120 189.930 ;
        RECT 121.590 189.590 122.740 189.730 ;
        RECT 121.590 189.530 121.910 189.590 ;
        RECT 123.905 189.545 124.195 189.775 ;
        RECT 128.580 189.730 128.720 189.930 ;
        RECT 129.425 189.885 129.715 190.115 ;
        RECT 129.960 190.070 130.100 190.270 ;
        RECT 130.330 190.210 130.650 190.470 ;
        RECT 131.250 190.210 131.570 190.470 ;
        RECT 131.800 190.455 131.940 190.610 ;
        RECT 131.725 190.225 132.015 190.455 ;
        RECT 131.340 190.070 131.480 190.210 ;
        RECT 129.960 189.930 131.480 190.070 ;
        RECT 129.500 189.730 129.640 189.885 ;
        RECT 128.580 189.590 129.640 189.730 ;
        RECT 11.120 188.910 151.295 189.390 ;
        RECT 13.965 188.710 14.255 188.755 ;
        RECT 14.870 188.710 15.190 188.770 ;
        RECT 13.965 188.570 15.190 188.710 ;
        RECT 13.965 188.525 14.255 188.570 ;
        RECT 14.870 188.510 15.190 188.570 ;
        RECT 25.465 188.525 25.755 188.755 ;
        RECT 17.170 188.170 17.490 188.430 ;
        RECT 18.265 188.370 18.555 188.415 ;
        RECT 19.010 188.370 19.330 188.430 ;
        RECT 24.530 188.415 24.850 188.430 ;
        RECT 18.265 188.230 19.330 188.370 ;
        RECT 18.265 188.185 18.555 188.230 ;
        RECT 19.010 188.170 19.330 188.230 ;
        RECT 23.625 188.185 23.915 188.415 ;
        RECT 24.530 188.185 24.915 188.415 ;
        RECT 16.265 187.690 16.555 187.735 ;
        RECT 20.390 187.690 20.710 187.750 ;
        RECT 16.265 187.550 20.710 187.690 ;
        RECT 23.700 187.690 23.840 188.185 ;
        RECT 24.530 188.170 24.850 188.185 ;
        RECT 25.540 188.030 25.680 188.525 ;
        RECT 25.910 188.510 26.230 188.770 ;
        RECT 52.605 188.710 52.895 188.755 ;
        RECT 54.065 188.710 54.355 188.755 ;
        RECT 52.605 188.570 54.355 188.710 ;
        RECT 52.605 188.525 52.895 188.570 ;
        RECT 54.065 188.525 54.355 188.570 ;
        RECT 54.905 188.710 55.195 188.755 ;
        RECT 55.350 188.710 55.670 188.770 ;
        RECT 61.790 188.710 62.110 188.770 ;
        RECT 62.265 188.710 62.555 188.755 ;
        RECT 54.905 188.570 55.670 188.710 ;
        RECT 54.905 188.525 55.195 188.570 ;
        RECT 55.350 188.510 55.670 188.570 ;
        RECT 55.900 188.570 61.560 188.710 ;
        RECT 30.970 188.370 31.290 188.430 ;
        RECT 52.130 188.370 52.450 188.430 ;
        RECT 53.065 188.370 53.355 188.415 ;
        RECT 29.220 188.230 53.355 188.370 ;
        RECT 26.845 188.030 27.135 188.075 ;
        RECT 25.540 187.890 27.135 188.030 ;
        RECT 26.845 187.845 27.135 187.890 ;
        RECT 29.220 187.690 29.360 188.230 ;
        RECT 30.970 188.170 31.290 188.230 ;
        RECT 52.130 188.170 52.450 188.230 ;
        RECT 53.065 188.185 53.355 188.230 ;
        RECT 53.510 188.170 53.830 188.430 ;
        RECT 55.900 188.370 56.040 188.570 ;
        RECT 56.730 188.415 57.050 188.430 ;
        RECT 56.700 188.370 57.050 188.415 ;
        RECT 54.060 188.230 56.040 188.370 ;
        RECT 56.535 188.230 57.050 188.370 ;
        RECT 30.510 187.830 30.830 188.090 ;
        RECT 31.430 188.030 31.750 188.090 ;
        RECT 35.110 188.030 35.430 188.090 ;
        RECT 31.430 187.890 35.430 188.030 ;
        RECT 31.430 187.830 31.750 187.890 ;
        RECT 35.110 187.830 35.430 187.890 ;
        RECT 41.550 187.830 41.870 188.090 ;
        RECT 47.530 188.030 47.850 188.090 ;
        RECT 50.305 188.030 50.595 188.075 ;
        RECT 47.530 187.890 50.595 188.030 ;
        RECT 47.530 187.830 47.850 187.890 ;
        RECT 50.305 187.845 50.595 187.890 ;
        RECT 51.670 187.830 51.990 188.090 ;
        RECT 52.605 188.030 52.895 188.075 ;
        RECT 53.600 188.030 53.740 188.170 ;
        RECT 52.605 187.890 53.740 188.030 ;
        RECT 52.605 187.845 52.895 187.890 ;
        RECT 23.700 187.550 29.360 187.690 ;
        RECT 16.265 187.505 16.555 187.550 ;
        RECT 20.390 187.490 20.710 187.550 ;
        RECT 42.010 187.490 42.330 187.750 ;
        RECT 49.830 187.690 50.150 187.750 ;
        RECT 54.060 187.690 54.200 188.230 ;
        RECT 56.700 188.185 57.050 188.230 ;
        RECT 56.730 188.170 57.050 188.185 ;
        RECT 55.365 188.030 55.655 188.075 ;
        RECT 55.810 188.030 56.130 188.090 ;
        RECT 55.365 187.890 56.130 188.030 ;
        RECT 61.420 188.030 61.560 188.570 ;
        RECT 61.790 188.570 62.555 188.710 ;
        RECT 61.790 188.510 62.110 188.570 ;
        RECT 62.265 188.525 62.555 188.570 ;
        RECT 65.010 188.710 65.330 188.770 ;
        RECT 67.770 188.710 68.090 188.770 ;
        RECT 73.290 188.710 73.610 188.770 ;
        RECT 65.010 188.570 68.090 188.710 ;
        RECT 65.010 188.510 65.330 188.570 ;
        RECT 67.770 188.510 68.090 188.570 ;
        RECT 68.320 188.570 73.610 188.710 ;
        RECT 63.980 188.370 64.270 188.415 ;
        RECT 65.100 188.370 65.240 188.510 ;
        RECT 68.320 188.370 68.460 188.570 ;
        RECT 73.290 188.510 73.610 188.570 ;
        RECT 73.765 188.525 74.055 188.755 ;
        RECT 73.840 188.370 73.980 188.525 ;
        RECT 77.430 188.510 77.750 188.770 ;
        RECT 78.350 188.710 78.670 188.770 ;
        RECT 77.980 188.570 78.670 188.710 ;
        RECT 77.980 188.415 78.120 188.570 ;
        RECT 78.350 188.510 78.670 188.570 ;
        RECT 78.810 188.710 79.130 188.770 ;
        RECT 94.925 188.710 95.215 188.755 ;
        RECT 97.670 188.710 97.990 188.770 ;
        RECT 78.810 188.570 81.340 188.710 ;
        RECT 78.810 188.510 79.130 188.570 ;
        RECT 63.980 188.230 65.240 188.370 ;
        RECT 66.940 188.230 68.460 188.370 ;
        RECT 68.600 188.230 71.220 188.370 ;
        RECT 73.840 188.230 74.440 188.370 ;
        RECT 63.980 188.185 64.270 188.230 ;
        RECT 64.565 188.030 64.855 188.075 ;
        RECT 66.940 188.030 67.080 188.230 ;
        RECT 61.420 187.890 67.080 188.030 ;
        RECT 67.310 188.030 67.630 188.090 ;
        RECT 68.600 188.075 68.740 188.230 ;
        RECT 71.080 188.090 71.220 188.230 ;
        RECT 67.785 188.030 68.075 188.075 ;
        RECT 67.310 187.890 68.075 188.030 ;
        RECT 55.365 187.845 55.655 187.890 ;
        RECT 55.810 187.830 56.130 187.890 ;
        RECT 64.565 187.845 64.855 187.890 ;
        RECT 67.310 187.830 67.630 187.890 ;
        RECT 67.785 187.845 68.075 187.890 ;
        RECT 68.525 187.845 68.815 188.075 ;
        RECT 69.150 187.830 69.470 188.090 ;
        RECT 69.610 187.830 69.930 188.090 ;
        RECT 70.070 188.075 70.390 188.090 ;
        RECT 70.070 187.845 70.595 188.075 ;
        RECT 70.070 187.830 70.390 187.845 ;
        RECT 70.990 187.830 71.310 188.090 ;
        RECT 72.830 188.075 73.150 188.090 ;
        RECT 71.465 187.845 71.755 188.075 ;
        RECT 72.810 188.030 73.150 188.075 ;
        RECT 72.810 187.890 73.310 188.030 ;
        RECT 72.810 187.845 73.150 187.890 ;
        RECT 49.830 187.550 54.200 187.690 ;
        RECT 56.245 187.690 56.535 187.735 ;
        RECT 57.435 187.690 57.725 187.735 ;
        RECT 59.955 187.690 60.245 187.735 ;
        RECT 56.245 187.550 60.245 187.690 ;
        RECT 49.830 187.490 50.150 187.550 ;
        RECT 56.245 187.505 56.535 187.550 ;
        RECT 57.435 187.505 57.725 187.550 ;
        RECT 59.955 187.505 60.245 187.550 ;
        RECT 65.010 187.490 65.330 187.750 ;
        RECT 66.405 187.690 66.695 187.735 ;
        RECT 66.850 187.690 67.170 187.750 ;
        RECT 66.405 187.550 67.170 187.690 ;
        RECT 66.405 187.505 66.695 187.550 ;
        RECT 66.850 187.490 67.170 187.550 ;
        RECT 71.485 187.410 71.625 187.845 ;
        RECT 72.830 187.830 73.150 187.845 ;
        RECT 73.750 187.830 74.070 188.090 ;
        RECT 74.300 188.075 74.440 188.230 ;
        RECT 77.905 188.185 78.195 188.415 ;
        RECT 74.255 187.845 74.545 188.075 ;
        RECT 75.130 188.030 75.450 188.090 ;
        RECT 81.200 188.075 81.340 188.570 ;
        RECT 94.925 188.570 97.990 188.710 ;
        RECT 94.925 188.525 95.215 188.570 ;
        RECT 82.965 188.370 83.255 188.415 ;
        RECT 83.410 188.370 83.730 188.430 ;
        RECT 82.965 188.230 83.730 188.370 ;
        RECT 82.965 188.185 83.255 188.230 ;
        RECT 83.410 188.170 83.730 188.230 ;
        RECT 83.885 188.370 84.175 188.415 ;
        RECT 84.790 188.370 85.110 188.430 ;
        RECT 83.885 188.230 85.110 188.370 ;
        RECT 83.885 188.185 84.175 188.230 ;
        RECT 84.790 188.170 85.110 188.230 ;
        RECT 86.170 188.170 86.490 188.430 ;
        RECT 95.000 188.370 95.140 188.525 ;
        RECT 97.670 188.510 97.990 188.570 ;
        RECT 100.445 188.525 100.735 188.755 ;
        RECT 113.310 188.710 113.630 188.770 ;
        RECT 116.085 188.710 116.375 188.755 ;
        RECT 113.310 188.570 116.375 188.710 ;
        RECT 94.080 188.230 95.140 188.370 ;
        RECT 98.605 188.370 98.895 188.415 ;
        RECT 100.520 188.370 100.660 188.525 ;
        RECT 113.310 188.510 113.630 188.570 ;
        RECT 116.085 188.525 116.375 188.570 ;
        RECT 116.530 188.510 116.850 188.770 ;
        RECT 105.965 188.370 106.255 188.415 ;
        RECT 117.910 188.370 118.230 188.430 ;
        RECT 98.605 188.230 100.660 188.370 ;
        RECT 101.210 188.230 106.255 188.370 ;
        RECT 76.065 188.030 76.355 188.075 ;
        RECT 75.130 187.890 76.355 188.030 ;
        RECT 75.130 187.830 75.450 187.890 ;
        RECT 76.065 187.845 76.355 187.890 ;
        RECT 76.600 187.890 77.820 188.030 ;
        RECT 72.385 187.690 72.675 187.735 ;
        RECT 73.840 187.690 73.980 187.830 ;
        RECT 76.600 187.690 76.740 187.890 ;
        RECT 72.385 187.550 73.980 187.690 ;
        RECT 76.140 187.550 76.740 187.690 ;
        RECT 77.680 187.690 77.820 187.890 ;
        RECT 80.205 187.845 80.495 188.075 ;
        RECT 81.125 187.845 81.415 188.075 ;
        RECT 80.280 187.690 80.420 187.845 ;
        RECT 82.490 187.830 82.810 188.090 ;
        RECT 85.265 188.030 85.555 188.075 ;
        RECT 86.260 188.030 86.400 188.170 ;
        RECT 85.265 187.890 86.400 188.030 ;
        RECT 85.265 187.845 85.555 187.890 ;
        RECT 88.025 187.845 88.315 188.075 ;
        RECT 82.030 187.690 82.350 187.750 ;
        RECT 77.680 187.550 82.350 187.690 ;
        RECT 72.385 187.505 72.675 187.550 ;
        RECT 14.885 187.350 15.175 187.395 ;
        RECT 19.025 187.350 19.315 187.395 ;
        RECT 22.690 187.350 23.010 187.410 ;
        RECT 14.885 187.210 16.940 187.350 ;
        RECT 14.885 187.165 15.175 187.210 ;
        RECT 16.800 187.070 16.940 187.210 ;
        RECT 19.025 187.210 23.010 187.350 ;
        RECT 19.025 187.165 19.315 187.210 ;
        RECT 22.690 187.150 23.010 187.210 ;
        RECT 43.405 187.350 43.695 187.395 ;
        RECT 55.850 187.350 56.140 187.395 ;
        RECT 57.950 187.350 58.240 187.395 ;
        RECT 59.520 187.350 59.810 187.395 ;
        RECT 43.405 187.210 54.660 187.350 ;
        RECT 43.405 187.165 43.695 187.210 ;
        RECT 16.710 187.010 17.030 187.070 ;
        RECT 18.105 187.010 18.395 187.055 ;
        RECT 16.710 186.870 18.395 187.010 ;
        RECT 16.710 186.810 17.030 186.870 ;
        RECT 18.105 186.825 18.395 186.870 ;
        RECT 24.545 187.010 24.835 187.055 ;
        RECT 27.290 187.010 27.610 187.070 ;
        RECT 24.545 186.870 27.610 187.010 ;
        RECT 24.545 186.825 24.835 186.870 ;
        RECT 27.290 186.810 27.610 186.870 ;
        RECT 30.970 186.810 31.290 187.070 ;
        RECT 53.050 187.010 53.370 187.070 ;
        RECT 53.985 187.010 54.275 187.055 ;
        RECT 53.050 186.870 54.275 187.010 ;
        RECT 54.520 187.010 54.660 187.210 ;
        RECT 55.850 187.210 59.810 187.350 ;
        RECT 55.850 187.165 56.140 187.210 ;
        RECT 57.950 187.165 58.240 187.210 ;
        RECT 59.520 187.165 59.810 187.210 ;
        RECT 71.005 187.165 71.295 187.395 ;
        RECT 58.570 187.010 58.890 187.070 ;
        RECT 54.520 186.870 58.890 187.010 ;
        RECT 53.050 186.810 53.370 186.870 ;
        RECT 53.985 186.825 54.275 186.870 ;
        RECT 58.570 186.810 58.890 186.870 ;
        RECT 61.790 187.010 62.110 187.070 ;
        RECT 63.185 187.010 63.475 187.055 ;
        RECT 61.790 186.870 63.475 187.010 ;
        RECT 61.790 186.810 62.110 186.870 ;
        RECT 63.185 186.825 63.475 186.870 ;
        RECT 66.390 187.010 66.710 187.070 ;
        RECT 71.080 187.010 71.220 187.165 ;
        RECT 71.450 187.150 71.770 187.410 ;
        RECT 74.210 187.150 74.530 187.410 ;
        RECT 66.390 186.870 71.220 187.010 ;
        RECT 72.845 187.010 73.135 187.055 ;
        RECT 76.140 187.010 76.280 187.550 ;
        RECT 82.030 187.490 82.350 187.550 ;
        RECT 78.350 187.350 78.670 187.410 ;
        RECT 79.285 187.350 79.575 187.395 ;
        RECT 88.100 187.350 88.240 187.845 ;
        RECT 92.150 187.830 92.470 188.090 ;
        RECT 92.610 188.030 92.930 188.090 ;
        RECT 94.080 188.075 94.220 188.230 ;
        RECT 98.605 188.185 98.895 188.230 ;
        RECT 92.610 187.890 93.125 188.030 ;
        RECT 92.610 187.830 92.930 187.890 ;
        RECT 94.005 187.845 94.295 188.075 ;
        RECT 94.450 187.830 94.770 188.090 ;
        RECT 94.910 188.030 95.230 188.090 ;
        RECT 97.225 188.030 97.515 188.075 ;
        RECT 94.910 187.890 97.515 188.030 ;
        RECT 94.910 187.830 95.230 187.890 ;
        RECT 97.225 187.845 97.515 187.890 ;
        RECT 97.685 188.030 97.975 188.075 ;
        RECT 99.970 188.030 100.290 188.090 ;
        RECT 97.685 187.890 100.290 188.030 ;
        RECT 97.685 187.845 97.975 187.890 ;
        RECT 99.970 187.830 100.290 187.890 ;
        RECT 100.430 188.030 100.750 188.090 ;
        RECT 101.210 188.075 101.350 188.230 ;
        RECT 105.965 188.185 106.255 188.230 ;
        RECT 115.700 188.230 118.230 188.370 ;
        RECT 101.135 188.030 101.425 188.075 ;
        RECT 100.430 187.890 101.425 188.030 ;
        RECT 100.430 187.830 100.750 187.890 ;
        RECT 101.135 187.845 101.425 187.890 ;
        RECT 101.810 187.830 102.130 188.090 ;
        RECT 102.270 187.830 102.590 188.090 ;
        RECT 102.730 188.075 103.050 188.090 ;
        RECT 102.730 187.845 103.215 188.075 ;
        RECT 102.730 187.830 103.050 187.845 ;
        RECT 103.650 187.830 103.970 188.090 ;
        RECT 115.700 188.075 115.840 188.230 ;
        RECT 117.910 188.170 118.230 188.230 ;
        RECT 106.425 188.030 106.715 188.075 ;
        RECT 115.625 188.030 115.915 188.075 ;
        RECT 106.425 187.890 115.915 188.030 ;
        RECT 106.425 187.845 106.715 187.890 ;
        RECT 115.625 187.845 115.915 187.890 ;
        RECT 91.245 187.690 91.535 187.735 ;
        RECT 98.590 187.690 98.910 187.750 ;
        RECT 91.245 187.550 98.910 187.690 ;
        RECT 91.245 187.505 91.535 187.550 ;
        RECT 98.590 187.490 98.910 187.550 ;
        RECT 93.545 187.350 93.835 187.395 ;
        RECT 114.705 187.350 114.995 187.395 ;
        RECT 116.990 187.350 117.310 187.410 ;
        RECT 78.350 187.210 79.575 187.350 ;
        RECT 78.350 187.150 78.670 187.210 ;
        RECT 79.285 187.165 79.575 187.210 ;
        RECT 83.500 187.210 92.840 187.350 ;
        RECT 72.845 186.870 76.280 187.010 ;
        RECT 66.390 186.810 66.710 186.870 ;
        RECT 72.845 186.825 73.135 186.870 ;
        RECT 76.510 186.810 76.830 187.070 ;
        RECT 76.970 186.810 77.290 187.070 ;
        RECT 80.650 187.010 80.970 187.070 ;
        RECT 82.045 187.010 82.335 187.055 ;
        RECT 83.500 187.010 83.640 187.210 ;
        RECT 92.700 187.070 92.840 187.210 ;
        RECT 93.545 187.210 103.420 187.350 ;
        RECT 93.545 187.165 93.835 187.210 ;
        RECT 103.280 187.070 103.420 187.210 ;
        RECT 104.200 187.210 117.310 187.350 ;
        RECT 104.200 187.070 104.340 187.210 ;
        RECT 114.705 187.165 114.995 187.210 ;
        RECT 116.990 187.150 117.310 187.210 ;
        RECT 80.650 186.870 83.640 187.010 ;
        RECT 80.650 186.810 80.970 186.870 ;
        RECT 82.045 186.825 82.335 186.870 ;
        RECT 83.870 186.810 84.190 187.070 ;
        RECT 87.550 186.810 87.870 187.070 ;
        RECT 92.610 186.810 92.930 187.070 ;
        RECT 96.290 186.810 96.610 187.070 ;
        RECT 98.605 187.010 98.895 187.055 ;
        RECT 99.050 187.010 99.370 187.070 ;
        RECT 98.605 186.870 99.370 187.010 ;
        RECT 98.605 186.825 98.895 186.870 ;
        RECT 99.050 186.810 99.370 186.870 ;
        RECT 103.190 186.810 103.510 187.070 ;
        RECT 104.110 186.810 104.430 187.070 ;
        RECT 117.450 186.810 117.770 187.070 ;
        RECT 11.120 186.190 150.500 186.670 ;
        RECT 17.170 185.790 17.490 186.050 ;
        RECT 19.010 185.790 19.330 186.050 ;
        RECT 24.530 185.790 24.850 186.050 ;
        RECT 26.830 185.790 27.150 186.050 ;
        RECT 27.290 185.790 27.610 186.050 ;
        RECT 30.970 185.790 31.290 186.050 ;
        RECT 38.330 185.990 38.650 186.050 ;
        RECT 39.250 185.990 39.570 186.050 ;
        RECT 40.185 185.990 40.475 186.035 ;
        RECT 35.200 185.850 38.100 185.990 ;
        RECT 17.260 185.650 17.400 185.790 ;
        RECT 19.945 185.650 20.235 185.695 ;
        RECT 17.260 185.510 20.235 185.650 ;
        RECT 19.945 185.465 20.235 185.510 ;
        RECT 26.920 185.310 27.060 185.790 ;
        RECT 17.260 185.170 20.620 185.310 ;
        RECT 17.260 185.015 17.400 185.170 ;
        RECT 20.480 185.030 20.620 185.170 ;
        RECT 22.320 185.170 27.980 185.310 ;
        RECT 17.185 184.785 17.475 185.015 ;
        RECT 18.105 184.970 18.395 185.015 ;
        RECT 19.485 184.970 19.775 185.015 ;
        RECT 18.105 184.830 19.775 184.970 ;
        RECT 18.105 184.785 18.395 184.830 ;
        RECT 19.485 184.785 19.775 184.830 ;
        RECT 20.390 184.970 20.710 185.030 ;
        RECT 22.320 184.970 22.460 185.170 ;
        RECT 20.390 184.830 22.460 184.970 ;
        RECT 19.560 184.630 19.700 184.785 ;
        RECT 20.390 184.770 20.710 184.830 ;
        RECT 25.450 184.770 25.770 185.030 ;
        RECT 26.920 185.015 27.060 185.170 ;
        RECT 27.840 185.015 27.980 185.170 ;
        RECT 26.845 184.785 27.135 185.015 ;
        RECT 27.305 184.785 27.595 185.015 ;
        RECT 27.765 184.785 28.055 185.015 ;
        RECT 31.060 184.970 31.200 185.790 ;
        RECT 35.200 185.695 35.340 185.850 ;
        RECT 35.125 185.465 35.415 185.695 ;
        RECT 37.960 185.650 38.100 185.850 ;
        RECT 38.330 185.850 40.475 185.990 ;
        RECT 38.330 185.790 38.650 185.850 ;
        RECT 39.250 185.790 39.570 185.850 ;
        RECT 40.185 185.805 40.475 185.850 ;
        RECT 42.930 185.990 43.250 186.050 ;
        RECT 48.005 185.990 48.295 186.035 ;
        RECT 42.930 185.850 48.295 185.990 ;
        RECT 42.930 185.790 43.250 185.850 ;
        RECT 48.005 185.805 48.295 185.850 ;
        RECT 53.050 185.990 53.370 186.050 ;
        RECT 57.650 185.990 57.970 186.050 ;
        RECT 60.410 185.990 60.730 186.050 ;
        RECT 53.050 185.850 60.730 185.990 ;
        RECT 53.050 185.790 53.370 185.850 ;
        RECT 57.650 185.790 57.970 185.850 ;
        RECT 60.410 185.790 60.730 185.850 ;
        RECT 64.565 185.990 64.855 186.035 ;
        RECT 65.470 185.990 65.790 186.050 ;
        RECT 64.565 185.850 65.790 185.990 ;
        RECT 64.565 185.805 64.855 185.850 ;
        RECT 65.470 185.790 65.790 185.850 ;
        RECT 67.310 185.790 67.630 186.050 ;
        RECT 67.770 185.790 68.090 186.050 ;
        RECT 69.150 185.790 69.470 186.050 ;
        RECT 71.005 185.990 71.295 186.035 ;
        RECT 71.450 185.990 71.770 186.050 ;
        RECT 71.005 185.850 71.770 185.990 ;
        RECT 71.005 185.805 71.295 185.850 ;
        RECT 71.450 185.790 71.770 185.850 ;
        RECT 72.845 185.990 73.135 186.035 ;
        RECT 77.445 185.990 77.735 186.035 ;
        RECT 72.845 185.850 76.280 185.990 ;
        RECT 72.845 185.805 73.135 185.850 ;
        RECT 41.090 185.650 41.410 185.710 ;
        RECT 37.960 185.510 41.410 185.650 ;
        RECT 41.090 185.450 41.410 185.510 ;
        RECT 42.485 185.650 42.775 185.695 ;
        RECT 47.085 185.650 47.375 185.695 ;
        RECT 66.390 185.650 66.710 185.710 ;
        RECT 42.485 185.510 47.375 185.650 ;
        RECT 42.485 185.465 42.775 185.510 ;
        RECT 47.085 185.465 47.375 185.510 ;
        RECT 51.760 185.510 66.710 185.650 ;
        RECT 31.905 185.310 32.195 185.355 ;
        RECT 36.045 185.310 36.335 185.355 ;
        RECT 40.170 185.310 40.490 185.370 ;
        RECT 31.905 185.170 33.960 185.310 ;
        RECT 31.905 185.125 32.195 185.170 ;
        RECT 32.365 184.970 32.655 185.015 ;
        RECT 28.300 184.830 30.695 184.970 ;
        RECT 31.060 184.830 32.655 184.970 ;
        RECT 26.370 184.630 26.690 184.690 ;
        RECT 27.380 184.630 27.520 184.785 ;
        RECT 28.300 184.630 28.440 184.830 ;
        RECT 19.560 184.490 28.440 184.630 ;
        RECT 26.370 184.430 26.690 184.490 ;
        RECT 28.685 184.445 28.975 184.675 ;
        RECT 25.450 184.290 25.770 184.350 ;
        RECT 28.760 184.290 28.900 184.445 ;
        RECT 30.050 184.430 30.370 184.690 ;
        RECT 30.555 184.630 30.695 184.830 ;
        RECT 32.365 184.785 32.655 184.830 ;
        RECT 32.810 184.970 33.130 185.030 ;
        RECT 33.820 185.015 33.960 185.170 ;
        RECT 34.740 185.170 36.335 185.310 ;
        RECT 33.285 184.970 33.575 185.015 ;
        RECT 32.810 184.830 33.575 184.970 ;
        RECT 32.810 184.770 33.130 184.830 ;
        RECT 33.285 184.785 33.575 184.830 ;
        RECT 33.745 184.785 34.035 185.015 ;
        RECT 34.205 184.980 34.495 185.015 ;
        RECT 34.740 184.980 34.880 185.170 ;
        RECT 36.045 185.125 36.335 185.170 ;
        RECT 36.580 185.170 40.490 185.310 ;
        RECT 34.205 184.840 34.880 184.980 ;
        RECT 35.110 184.970 35.430 185.030 ;
        RECT 36.580 185.015 36.720 185.170 ;
        RECT 40.170 185.110 40.490 185.170 ;
        RECT 40.630 185.110 40.950 185.370 ;
        RECT 47.160 185.310 47.300 185.465 ;
        RECT 51.760 185.355 51.900 185.510 ;
        RECT 66.390 185.450 66.710 185.510 ;
        RECT 47.160 185.170 51.440 185.310 ;
        RECT 35.585 184.970 35.875 185.015 ;
        RECT 34.205 184.785 34.495 184.840 ;
        RECT 35.110 184.830 35.875 184.970 ;
        RECT 35.110 184.770 35.430 184.830 ;
        RECT 35.585 184.785 35.875 184.830 ;
        RECT 36.505 184.785 36.795 185.015 ;
        RECT 37.425 184.785 37.715 185.015 ;
        RECT 39.265 184.970 39.555 185.015 ;
        RECT 40.260 184.970 40.400 185.110 ;
        RECT 41.565 184.970 41.855 185.015 ;
        RECT 39.265 184.830 41.855 184.970 ;
        RECT 39.265 184.785 39.555 184.830 ;
        RECT 41.565 184.785 41.855 184.830 ;
        RECT 46.625 184.970 46.915 185.015 ;
        RECT 48.450 184.970 48.770 185.030 ;
        RECT 51.300 185.015 51.440 185.170 ;
        RECT 51.685 185.125 51.975 185.355 ;
        RECT 52.130 185.110 52.450 185.370 ;
        RECT 67.400 185.310 67.540 185.790 ;
        RECT 64.180 185.170 67.540 185.310 ;
        RECT 67.860 185.650 68.000 185.790 ;
        RECT 72.920 185.650 73.060 185.805 ;
        RECT 67.860 185.510 73.060 185.650 ;
        RECT 50.765 184.980 51.055 185.015 ;
        RECT 46.625 184.830 48.770 184.970 ;
        RECT 46.625 184.785 46.915 184.830 ;
        RECT 30.985 184.630 31.275 184.675 ;
        RECT 36.580 184.630 36.720 184.785 ;
        RECT 30.555 184.490 36.720 184.630 ;
        RECT 37.500 184.630 37.640 184.785 ;
        RECT 48.450 184.770 48.770 184.830 ;
        RECT 50.380 184.840 51.055 184.980 ;
        RECT 40.185 184.630 40.475 184.675 ;
        RECT 42.010 184.630 42.330 184.690 ;
        RECT 37.500 184.490 42.330 184.630 ;
        RECT 30.985 184.445 31.275 184.490 ;
        RECT 40.185 184.445 40.475 184.490 ;
        RECT 42.010 184.430 42.330 184.490 ;
        RECT 46.165 184.630 46.455 184.675 ;
        RECT 47.070 184.630 47.390 184.690 ;
        RECT 46.165 184.490 47.390 184.630 ;
        RECT 46.165 184.445 46.455 184.490 ;
        RECT 47.070 184.430 47.390 184.490 ;
        RECT 48.005 184.630 48.295 184.675 ;
        RECT 49.830 184.630 50.150 184.690 ;
        RECT 48.005 184.490 50.150 184.630 ;
        RECT 50.380 184.630 50.520 184.840 ;
        RECT 50.765 184.785 51.055 184.840 ;
        RECT 51.225 184.785 51.515 185.015 ;
        RECT 56.730 184.970 57.050 185.030 ;
        RECT 53.140 184.860 57.050 184.970 ;
        RECT 51.760 184.830 57.050 184.860 ;
        RECT 51.760 184.720 53.280 184.830 ;
        RECT 56.730 184.770 57.050 184.830 ;
        RECT 61.790 184.970 62.110 185.030 ;
        RECT 64.180 185.015 64.320 185.170 ;
        RECT 63.185 184.970 63.475 185.015 ;
        RECT 61.790 184.830 63.475 184.970 ;
        RECT 61.790 184.770 62.110 184.830 ;
        RECT 63.185 184.785 63.475 184.830 ;
        RECT 64.105 184.785 64.395 185.015 ;
        RECT 64.565 184.785 64.855 185.015 ;
        RECT 67.325 184.970 67.615 185.015 ;
        RECT 67.860 184.970 68.000 185.510 ;
        RECT 71.910 185.310 72.230 185.370 ;
        RECT 76.140 185.310 76.280 185.850 ;
        RECT 77.445 185.850 79.960 185.990 ;
        RECT 77.445 185.805 77.735 185.850 ;
        RECT 76.510 185.650 76.830 185.710 ;
        RECT 77.905 185.650 78.195 185.695 ;
        RECT 76.510 185.510 78.195 185.650 ;
        RECT 76.510 185.450 76.830 185.510 ;
        RECT 77.905 185.465 78.195 185.510 ;
        RECT 78.350 185.450 78.670 185.710 ;
        RECT 79.820 185.650 79.960 185.850 ;
        RECT 90.310 185.790 90.630 186.050 ;
        RECT 101.825 185.990 102.115 186.035 ;
        RECT 103.650 185.990 103.970 186.050 ;
        RECT 109.185 185.990 109.475 186.035 ;
        RECT 112.390 185.990 112.710 186.050 ;
        RECT 101.825 185.850 103.970 185.990 ;
        RECT 101.825 185.805 102.115 185.850 ;
        RECT 103.650 185.790 103.970 185.850 ;
        RECT 104.200 185.850 112.710 185.990 ;
        RECT 84.790 185.650 85.110 185.710 ;
        RECT 89.405 185.650 89.695 185.695 ;
        RECT 79.820 185.510 85.110 185.650 ;
        RECT 84.790 185.450 85.110 185.510 ;
        RECT 86.260 185.510 89.695 185.650 ;
        RECT 71.910 185.170 73.060 185.310 ;
        RECT 76.140 185.170 77.660 185.310 ;
        RECT 71.910 185.110 72.230 185.170 ;
        RECT 67.325 184.830 68.000 184.970 ;
        RECT 68.245 184.970 68.535 185.015 ;
        RECT 72.370 184.970 72.690 185.030 ;
        RECT 72.920 185.015 73.060 185.170 ;
        RECT 68.245 184.830 72.690 184.970 ;
        RECT 67.325 184.785 67.615 184.830 ;
        RECT 68.245 184.785 68.535 184.830 ;
        RECT 51.760 184.630 51.900 184.720 ;
        RECT 50.380 184.490 51.900 184.630 ;
        RECT 48.005 184.445 48.295 184.490 ;
        RECT 49.830 184.430 50.150 184.490 ;
        RECT 31.430 184.290 31.750 184.350 ;
        RECT 37.410 184.290 37.730 184.350 ;
        RECT 37.885 184.290 38.175 184.335 ;
        RECT 25.450 184.150 38.175 184.290 ;
        RECT 25.450 184.090 25.770 184.150 ;
        RECT 31.430 184.090 31.750 184.150 ;
        RECT 37.410 184.090 37.730 184.150 ;
        RECT 37.885 184.105 38.175 184.150 ;
        RECT 38.330 184.090 38.650 184.350 ;
        RECT 39.265 184.290 39.555 184.335 ;
        RECT 52.130 184.290 52.450 184.350 ;
        RECT 39.265 184.150 52.450 184.290 ;
        RECT 39.265 184.105 39.555 184.150 ;
        RECT 52.130 184.090 52.450 184.150 ;
        RECT 53.050 184.090 53.370 184.350 ;
        RECT 64.640 184.290 64.780 184.785 ;
        RECT 72.370 184.770 72.690 184.830 ;
        RECT 72.845 184.785 73.135 185.015 ;
        RECT 66.850 184.630 67.170 184.690 ;
        RECT 75.130 184.630 75.450 184.690 ;
        RECT 76.985 184.630 77.275 184.675 ;
        RECT 66.850 184.490 71.625 184.630 ;
        RECT 66.850 184.430 67.170 184.490 ;
        RECT 70.990 184.290 71.310 184.350 ;
        RECT 64.640 184.150 71.310 184.290 ;
        RECT 71.485 184.290 71.625 184.490 ;
        RECT 75.130 184.490 77.275 184.630 ;
        RECT 77.520 184.630 77.660 185.170 ;
        RECT 78.440 185.015 78.580 185.450 ;
        RECT 86.260 185.355 86.400 185.510 ;
        RECT 89.405 185.465 89.695 185.510 ;
        RECT 103.190 185.650 103.510 185.710 ;
        RECT 104.200 185.650 104.340 185.850 ;
        RECT 109.185 185.805 109.475 185.850 ;
        RECT 112.390 185.790 112.710 185.850 ;
        RECT 120.210 185.790 120.530 186.050 ;
        RECT 103.190 185.510 104.340 185.650 ;
        RECT 105.030 185.650 105.350 185.710 ;
        RECT 108.725 185.650 109.015 185.695 ;
        RECT 105.030 185.510 109.015 185.650 ;
        RECT 103.190 185.450 103.510 185.510 ;
        RECT 105.030 185.450 105.350 185.510 ;
        RECT 108.725 185.465 109.015 185.510 ;
        RECT 109.630 185.450 109.950 185.710 ;
        RECT 111.930 185.650 112.250 185.710 ;
        RECT 110.180 185.510 112.250 185.650 ;
        RECT 86.185 185.125 86.475 185.355 ;
        RECT 87.550 185.110 87.870 185.370 ;
        RECT 99.510 185.310 99.830 185.370 ;
        RECT 99.510 185.170 103.880 185.310 ;
        RECT 99.510 185.110 99.830 185.170 ;
        RECT 103.740 185.030 103.880 185.170 ;
        RECT 104.110 185.110 104.430 185.370 ;
        RECT 110.180 185.310 110.320 185.510 ;
        RECT 111.930 185.450 112.250 185.510 ;
        RECT 114.230 185.650 114.550 185.710 ;
        RECT 120.300 185.650 120.440 185.790 ;
        RECT 128.070 185.650 128.360 185.695 ;
        RECT 130.170 185.650 130.460 185.695 ;
        RECT 131.740 185.650 132.030 185.695 ;
        RECT 114.230 185.510 120.900 185.650 ;
        RECT 114.230 185.450 114.550 185.510 ;
        RECT 109.720 185.170 110.320 185.310 ;
        RECT 111.485 185.310 111.775 185.355 ;
        RECT 119.290 185.310 119.610 185.370 ;
        RECT 120.760 185.355 120.900 185.510 ;
        RECT 128.070 185.510 132.030 185.650 ;
        RECT 128.070 185.465 128.360 185.510 ;
        RECT 130.170 185.465 130.460 185.510 ;
        RECT 131.740 185.465 132.030 185.510 ;
        RECT 120.225 185.310 120.515 185.355 ;
        RECT 111.485 185.170 120.515 185.310 ;
        RECT 78.365 184.785 78.655 185.015 ;
        RECT 78.825 184.970 79.115 185.015 ;
        RECT 79.270 184.970 79.590 185.030 ;
        RECT 82.490 184.970 82.810 185.030 ;
        RECT 78.825 184.830 82.810 184.970 ;
        RECT 78.825 184.785 79.115 184.830 ;
        RECT 79.270 184.770 79.590 184.830 ;
        RECT 82.490 184.770 82.810 184.830 ;
        RECT 85.725 184.785 86.015 185.015 ;
        RECT 80.650 184.630 80.970 184.690 ;
        RECT 77.520 184.490 80.970 184.630 ;
        RECT 75.130 184.430 75.450 184.490 ;
        RECT 76.985 184.445 77.275 184.490 ;
        RECT 80.650 184.430 80.970 184.490 ;
        RECT 72.830 184.290 73.150 184.350 ;
        RECT 79.745 184.290 80.035 184.335 ;
        RECT 85.800 184.290 85.940 184.785 ;
        RECT 103.650 184.770 103.970 185.030 ;
        RECT 108.145 184.970 108.435 185.015 ;
        RECT 109.720 184.980 109.860 185.170 ;
        RECT 111.485 185.125 111.775 185.170 ;
        RECT 110.230 184.980 110.520 185.015 ;
        RECT 104.890 184.830 109.400 184.970 ;
        RECT 109.720 184.840 110.520 184.980 ;
        RECT 110.180 184.830 110.520 184.840 ;
        RECT 91.245 184.630 91.535 184.675 ;
        RECT 99.050 184.630 99.370 184.690 ;
        RECT 104.890 184.630 105.030 184.830 ;
        RECT 108.145 184.785 108.435 184.830 ;
        RECT 91.245 184.490 105.030 184.630 ;
        RECT 91.245 184.445 91.535 184.490 ;
        RECT 99.050 184.430 99.370 184.490 ;
        RECT 71.485 184.150 85.940 184.290 ;
        RECT 90.245 184.290 90.535 184.335 ;
        RECT 90.770 184.290 91.090 184.350 ;
        RECT 90.245 184.150 91.090 184.290 ;
        RECT 109.260 184.290 109.400 184.830 ;
        RECT 110.230 184.785 110.520 184.830 ;
        RECT 111.010 184.970 111.330 185.030 ;
        RECT 111.010 184.830 113.080 184.970 ;
        RECT 111.010 184.770 111.330 184.830 ;
        RECT 109.630 184.630 109.950 184.690 ;
        RECT 111.945 184.630 112.235 184.675 ;
        RECT 109.630 184.490 112.235 184.630 ;
        RECT 112.940 184.630 113.080 184.830 ;
        RECT 113.310 184.770 113.630 185.030 ;
        RECT 116.160 185.015 116.300 185.170 ;
        RECT 119.290 185.110 119.610 185.170 ;
        RECT 120.225 185.125 120.515 185.170 ;
        RECT 120.685 185.310 120.975 185.355 ;
        RECT 121.590 185.310 121.910 185.370 ;
        RECT 120.685 185.170 121.910 185.310 ;
        RECT 120.685 185.125 120.975 185.170 ;
        RECT 121.590 185.110 121.910 185.170 ;
        RECT 124.810 185.110 125.130 185.370 ;
        RECT 127.570 185.110 127.890 185.370 ;
        RECT 128.465 185.310 128.755 185.355 ;
        RECT 129.655 185.310 129.945 185.355 ;
        RECT 132.175 185.310 132.465 185.355 ;
        RECT 128.465 185.170 132.465 185.310 ;
        RECT 128.465 185.125 128.755 185.170 ;
        RECT 129.655 185.125 129.945 185.170 ;
        RECT 132.175 185.125 132.465 185.170 ;
        RECT 115.165 184.785 115.455 185.015 ;
        RECT 116.085 184.785 116.375 185.015 ;
        RECT 119.765 184.785 120.055 185.015 ;
        RECT 115.240 184.630 115.380 184.785 ;
        RECT 112.940 184.490 115.380 184.630 ;
        RECT 109.630 184.430 109.950 184.490 ;
        RECT 111.945 184.445 112.235 184.490 ;
        RECT 119.840 184.350 119.980 184.785 ;
        RECT 121.130 184.770 121.450 185.030 ;
        RECT 125.730 184.770 126.050 185.030 ;
        RECT 123.890 184.430 124.210 184.690 ;
        RECT 128.920 184.630 129.210 184.675 ;
        RECT 129.870 184.630 130.190 184.690 ;
        RECT 128.920 184.490 130.190 184.630 ;
        RECT 128.920 184.445 129.210 184.490 ;
        RECT 129.870 184.430 130.190 184.490 ;
        RECT 111.010 184.290 111.330 184.350 ;
        RECT 112.405 184.290 112.695 184.335 ;
        RECT 109.260 184.150 112.695 184.290 ;
        RECT 70.990 184.090 71.310 184.150 ;
        RECT 72.830 184.090 73.150 184.150 ;
        RECT 79.745 184.105 80.035 184.150 ;
        RECT 90.245 184.105 90.535 184.150 ;
        RECT 90.770 184.090 91.090 184.150 ;
        RECT 111.010 184.090 111.330 184.150 ;
        RECT 112.405 184.105 112.695 184.150 ;
        RECT 115.625 184.290 115.915 184.335 ;
        RECT 116.530 184.290 116.850 184.350 ;
        RECT 115.625 184.150 116.850 184.290 ;
        RECT 115.625 184.105 115.915 184.150 ;
        RECT 116.530 184.090 116.850 184.150 ;
        RECT 118.830 184.090 119.150 184.350 ;
        RECT 119.750 184.290 120.070 184.350 ;
        RECT 123.980 184.290 124.120 184.430 ;
        RECT 119.750 184.150 124.120 184.290 ;
        RECT 119.750 184.090 120.070 184.150 ;
        RECT 126.650 184.090 126.970 184.350 ;
        RECT 134.470 184.090 134.790 184.350 ;
        RECT 11.120 183.470 151.295 183.950 ;
        RECT 32.365 183.270 32.655 183.315 ;
        RECT 32.810 183.270 33.130 183.330 ;
        RECT 32.365 183.130 33.130 183.270 ;
        RECT 32.365 183.085 32.655 183.130 ;
        RECT 32.810 183.070 33.130 183.130 ;
        RECT 37.410 183.270 37.730 183.330 ;
        RECT 40.630 183.270 40.950 183.330 ;
        RECT 37.410 183.130 40.950 183.270 ;
        RECT 37.410 183.070 37.730 183.130 ;
        RECT 40.630 183.070 40.950 183.130 ;
        RECT 53.050 183.070 53.370 183.330 ;
        RECT 56.360 183.130 62.480 183.270 ;
        RECT 30.510 182.930 30.830 182.990 ;
        RECT 35.110 182.930 35.430 182.990 ;
        RECT 30.510 182.790 35.430 182.930 ;
        RECT 30.510 182.730 30.830 182.790 ;
        RECT 35.110 182.730 35.430 182.790 ;
        RECT 15.790 182.390 16.110 182.650 ;
        RECT 16.265 182.405 16.555 182.635 ;
        RECT 17.185 182.590 17.475 182.635 ;
        RECT 17.630 182.590 17.950 182.650 ;
        RECT 17.185 182.450 17.950 182.590 ;
        RECT 17.185 182.405 17.475 182.450 ;
        RECT 16.340 182.250 16.480 182.405 ;
        RECT 17.630 182.390 17.950 182.450 ;
        RECT 31.445 182.405 31.735 182.635 ;
        RECT 42.010 182.590 42.330 182.650 ;
        RECT 43.865 182.590 44.155 182.635 ;
        RECT 42.010 182.450 44.155 182.590 ;
        RECT 21.325 182.250 21.615 182.295 ;
        RECT 25.450 182.250 25.770 182.310 ;
        RECT 31.520 182.250 31.660 182.405 ;
        RECT 42.010 182.390 42.330 182.450 ;
        RECT 43.865 182.405 44.155 182.450 ;
        RECT 50.750 182.390 51.070 182.650 ;
        RECT 51.685 182.405 51.975 182.635 ;
        RECT 53.140 182.590 53.280 183.070 ;
        RECT 56.360 182.650 56.500 183.130 ;
        RECT 56.730 182.930 57.050 182.990 ;
        RECT 61.330 182.930 61.650 182.990 ;
        RECT 62.340 182.975 62.480 183.130 ;
        RECT 73.380 183.130 76.280 183.270 ;
        RECT 56.730 182.790 61.650 182.930 ;
        RECT 56.730 182.730 57.050 182.790 ;
        RECT 61.330 182.730 61.650 182.790 ;
        RECT 62.265 182.930 62.555 182.975 ;
        RECT 69.610 182.930 69.930 182.990 ;
        RECT 73.380 182.930 73.520 183.130 ;
        RECT 62.265 182.790 65.240 182.930 ;
        RECT 62.265 182.745 62.555 182.790 ;
        RECT 54.905 182.590 55.195 182.635 ;
        RECT 53.140 182.450 55.195 182.590 ;
        RECT 54.905 182.405 55.195 182.450 ;
        RECT 55.365 182.405 55.655 182.635 ;
        RECT 56.270 182.590 56.590 182.650 ;
        RECT 56.075 182.450 56.590 182.590 ;
        RECT 16.340 182.110 18.780 182.250 ;
        RECT 18.640 181.630 18.780 182.110 ;
        RECT 20.480 182.110 22.230 182.250 ;
        RECT 20.480 181.630 20.620 182.110 ;
        RECT 21.325 182.065 21.615 182.110 ;
        RECT 22.090 181.910 22.230 182.110 ;
        RECT 25.450 182.110 31.660 182.250 ;
        RECT 51.760 182.250 51.900 182.405 ;
        RECT 55.440 182.250 55.580 182.405 ;
        RECT 56.270 182.390 56.590 182.450 ;
        RECT 60.870 182.590 61.190 182.650 ;
        RECT 63.185 182.590 63.475 182.635 ;
        RECT 60.870 182.450 63.475 182.590 ;
        RECT 60.870 182.390 61.190 182.450 ;
        RECT 63.185 182.405 63.475 182.450 ;
        RECT 63.630 182.590 63.950 182.650 ;
        RECT 65.100 182.635 65.240 182.790 ;
        RECT 69.610 182.790 73.520 182.930 ;
        RECT 69.610 182.730 69.930 182.790 ;
        RECT 75.130 182.730 75.450 182.990 ;
        RECT 76.140 182.975 76.280 183.130 ;
        RECT 95.000 183.130 105.030 183.270 ;
        RECT 76.065 182.745 76.355 182.975 ;
        RECT 76.510 182.930 76.830 182.990 ;
        RECT 76.985 182.930 77.275 182.975 ;
        RECT 76.510 182.790 77.275 182.930 ;
        RECT 76.510 182.730 76.830 182.790 ;
        RECT 76.985 182.745 77.275 182.790 ;
        RECT 88.930 182.930 89.250 182.990 ;
        RECT 94.450 182.930 94.770 182.990 ;
        RECT 88.930 182.790 94.770 182.930 ;
        RECT 88.930 182.730 89.250 182.790 ;
        RECT 94.450 182.730 94.770 182.790 ;
        RECT 64.105 182.590 64.395 182.635 ;
        RECT 63.630 182.450 64.395 182.590 ;
        RECT 63.630 182.390 63.950 182.450 ;
        RECT 64.105 182.405 64.395 182.450 ;
        RECT 64.565 182.405 64.855 182.635 ;
        RECT 65.025 182.590 65.315 182.635 ;
        RECT 82.030 182.590 82.350 182.650 ;
        RECT 90.325 182.590 90.615 182.635 ;
        RECT 65.025 182.450 65.425 182.590 ;
        RECT 82.030 182.450 90.615 182.590 ;
        RECT 65.025 182.405 65.315 182.450 ;
        RECT 64.640 182.250 64.780 182.405 ;
        RECT 82.030 182.390 82.350 182.450 ;
        RECT 90.325 182.405 90.615 182.450 ;
        RECT 51.760 182.110 53.740 182.250 ;
        RECT 25.450 182.050 25.770 182.110 ;
        RECT 40.630 181.910 40.950 181.970 ;
        RECT 22.090 181.770 50.980 181.910 ;
        RECT 40.630 181.710 40.950 181.770 ;
        RECT 17.170 181.370 17.490 181.630 ;
        RECT 18.550 181.370 18.870 181.630 ;
        RECT 20.390 181.370 20.710 181.630 ;
        RECT 41.550 181.570 41.870 181.630 ;
        RECT 42.945 181.570 43.235 181.615 ;
        RECT 41.550 181.430 43.235 181.570 ;
        RECT 41.550 181.370 41.870 181.430 ;
        RECT 42.945 181.385 43.235 181.430 ;
        RECT 49.830 181.370 50.150 181.630 ;
        RECT 50.840 181.615 50.980 181.770 ;
        RECT 53.600 181.630 53.740 182.110 ;
        RECT 54.980 182.110 64.780 182.250 ;
        RECT 66.405 182.250 66.695 182.295 ;
        RECT 70.530 182.250 70.850 182.310 ;
        RECT 66.405 182.110 70.850 182.250 ;
        RECT 54.980 181.630 55.120 182.110 ;
        RECT 66.405 182.065 66.695 182.110 ;
        RECT 70.530 182.050 70.850 182.110 ;
        RECT 71.450 182.250 71.770 182.310 ;
        RECT 83.870 182.250 84.190 182.310 ;
        RECT 71.450 182.110 84.190 182.250 ;
        RECT 71.450 182.050 71.770 182.110 ;
        RECT 83.870 182.050 84.190 182.110 ;
        RECT 90.770 182.050 91.090 182.310 ;
        RECT 56.285 181.910 56.575 181.955 ;
        RECT 58.110 181.910 58.430 181.970 ;
        RECT 56.285 181.770 58.430 181.910 ;
        RECT 56.285 181.725 56.575 181.770 ;
        RECT 58.110 181.710 58.430 181.770 ;
        RECT 62.265 181.910 62.555 181.955 ;
        RECT 64.090 181.910 64.410 181.970 ;
        RECT 62.265 181.770 64.410 181.910 ;
        RECT 62.265 181.725 62.555 181.770 ;
        RECT 64.090 181.710 64.410 181.770 ;
        RECT 68.230 181.910 68.550 181.970 ;
        RECT 95.000 181.910 95.140 183.130 ;
        RECT 102.730 182.930 103.050 182.990 ;
        RECT 103.510 182.930 103.800 182.975 ;
        RECT 102.730 182.790 103.800 182.930 ;
        RECT 102.730 182.730 103.050 182.790 ;
        RECT 103.510 182.745 103.800 182.790 ;
        RECT 104.890 182.590 105.030 183.130 ;
        RECT 106.870 183.070 107.190 183.330 ;
        RECT 113.310 183.270 113.630 183.330 ;
        RECT 111.560 183.130 113.630 183.270 ;
        RECT 106.960 182.930 107.100 183.070 ;
        RECT 111.560 182.975 111.700 183.130 ;
        RECT 113.310 183.070 113.630 183.130 ;
        RECT 121.130 183.270 121.450 183.330 ;
        RECT 121.130 183.130 122.280 183.270 ;
        RECT 121.130 183.070 121.450 183.130 ;
        RECT 111.485 182.930 111.775 182.975 ;
        RECT 106.960 182.790 111.775 182.930 ;
        RECT 111.485 182.745 111.775 182.790 ;
        RECT 116.990 182.730 117.310 182.990 ;
        RECT 118.830 182.930 119.150 182.990 ;
        RECT 118.000 182.790 119.150 182.930 ;
        RECT 105.490 182.590 105.810 182.650 ;
        RECT 109.630 182.590 109.950 182.650 ;
        RECT 110.105 182.590 110.395 182.635 ;
        RECT 104.890 182.450 109.400 182.590 ;
        RECT 105.490 182.390 105.810 182.450 ;
        RECT 102.270 182.050 102.590 182.310 ;
        RECT 103.165 182.250 103.455 182.295 ;
        RECT 104.355 182.250 104.645 182.295 ;
        RECT 106.875 182.250 107.165 182.295 ;
        RECT 103.165 182.110 107.165 182.250 ;
        RECT 109.260 182.250 109.400 182.450 ;
        RECT 109.630 182.450 110.395 182.590 ;
        RECT 109.630 182.390 109.950 182.450 ;
        RECT 110.105 182.405 110.395 182.450 ;
        RECT 110.565 182.590 110.855 182.635 ;
        RECT 111.010 182.590 111.330 182.650 ;
        RECT 110.565 182.450 111.330 182.590 ;
        RECT 110.565 182.405 110.855 182.450 ;
        RECT 111.010 182.390 111.330 182.450 ;
        RECT 116.545 182.590 116.835 182.635 ;
        RECT 118.000 182.590 118.140 182.790 ;
        RECT 118.830 182.730 119.150 182.790 ;
        RECT 119.750 182.930 120.070 182.990 ;
        RECT 119.750 182.790 120.900 182.930 ;
        RECT 119.750 182.730 120.070 182.790 ;
        RECT 116.545 182.450 118.140 182.590 ;
        RECT 118.385 182.590 118.675 182.635 ;
        RECT 120.225 182.590 120.515 182.635 ;
        RECT 118.385 182.450 120.515 182.590 ;
        RECT 120.760 182.590 120.900 182.790 ;
        RECT 122.140 182.660 122.280 183.130 ;
        RECT 126.650 183.070 126.970 183.330 ;
        RECT 129.870 183.070 130.190 183.330 ;
        RECT 123.060 182.790 125.500 182.930 ;
        RECT 121.145 182.590 121.435 182.635 ;
        RECT 120.760 182.450 121.435 182.590 ;
        RECT 116.545 182.405 116.835 182.450 ;
        RECT 118.385 182.405 118.675 182.450 ;
        RECT 120.225 182.405 120.515 182.450 ;
        RECT 121.145 182.405 121.435 182.450 ;
        RECT 121.590 182.390 121.910 182.650 ;
        RECT 122.140 182.635 122.740 182.660 ;
        RECT 123.060 182.650 123.200 182.790 ;
        RECT 122.140 182.520 122.815 182.635 ;
        RECT 122.525 182.405 122.815 182.520 ;
        RECT 122.970 182.390 123.290 182.650 ;
        RECT 125.360 182.635 125.500 182.790 ;
        RECT 123.905 182.405 124.195 182.635 ;
        RECT 124.825 182.405 125.115 182.635 ;
        RECT 125.265 182.405 125.555 182.635 ;
        RECT 113.310 182.250 113.630 182.310 ;
        RECT 109.260 182.110 113.630 182.250 ;
        RECT 103.165 182.065 103.455 182.110 ;
        RECT 104.355 182.065 104.645 182.110 ;
        RECT 106.875 182.065 107.165 182.110 ;
        RECT 113.310 182.050 113.630 182.110 ;
        RECT 118.845 182.065 119.135 182.295 ;
        RECT 120.670 182.250 120.990 182.310 ;
        RECT 123.980 182.250 124.120 182.405 ;
        RECT 120.670 182.110 124.120 182.250 ;
        RECT 68.230 181.770 95.140 181.910 ;
        RECT 102.770 181.910 103.060 181.955 ;
        RECT 104.870 181.910 105.160 181.955 ;
        RECT 106.440 181.910 106.730 181.955 ;
        RECT 102.770 181.770 106.730 181.910 ;
        RECT 68.230 181.710 68.550 181.770 ;
        RECT 102.770 181.725 103.060 181.770 ;
        RECT 104.870 181.725 105.160 181.770 ;
        RECT 106.440 181.725 106.730 181.770 ;
        RECT 110.090 181.910 110.410 181.970 ;
        RECT 111.485 181.910 111.775 181.955 ;
        RECT 110.090 181.770 111.775 181.910 ;
        RECT 110.090 181.710 110.410 181.770 ;
        RECT 111.485 181.725 111.775 181.770 ;
        RECT 116.530 181.910 116.850 181.970 ;
        RECT 118.920 181.910 119.060 182.065 ;
        RECT 120.670 182.050 120.990 182.110 ;
        RECT 116.530 181.770 119.060 181.910 ;
        RECT 119.765 181.910 120.055 181.955 ;
        RECT 124.900 181.910 125.040 182.405 ;
        RECT 125.730 182.390 126.050 182.650 ;
        RECT 126.740 182.590 126.880 183.070 ;
        RECT 130.805 182.590 131.095 182.635 ;
        RECT 126.740 182.450 131.095 182.590 ;
        RECT 130.805 182.405 131.095 182.450 ;
        RECT 119.765 181.770 125.040 181.910 ;
        RECT 126.190 181.910 126.510 181.970 ;
        RECT 126.665 181.910 126.955 181.955 ;
        RECT 126.190 181.770 126.955 181.910 ;
        RECT 116.530 181.710 116.850 181.770 ;
        RECT 119.765 181.725 120.055 181.770 ;
        RECT 126.190 181.710 126.510 181.770 ;
        RECT 126.665 181.725 126.955 181.770 ;
        RECT 50.765 181.570 51.055 181.615 ;
        RECT 51.670 181.570 51.990 181.630 ;
        RECT 50.765 181.430 51.990 181.570 ;
        RECT 50.765 181.385 51.055 181.430 ;
        RECT 51.670 181.370 51.990 181.430 ;
        RECT 53.510 181.370 53.830 181.630 ;
        RECT 54.890 181.370 55.210 181.630 ;
        RECT 57.650 181.570 57.970 181.630 ;
        RECT 65.470 181.570 65.790 181.630 ;
        RECT 57.650 181.430 65.790 181.570 ;
        RECT 57.650 181.370 57.970 181.430 ;
        RECT 65.470 181.370 65.790 181.430 ;
        RECT 83.870 181.570 84.190 181.630 ;
        RECT 91.690 181.570 92.010 181.630 ;
        RECT 83.870 181.430 92.010 181.570 ;
        RECT 83.870 181.370 84.190 181.430 ;
        RECT 91.690 181.370 92.010 181.430 ;
        RECT 92.165 181.570 92.455 181.615 ;
        RECT 96.750 181.570 97.070 181.630 ;
        RECT 92.165 181.430 97.070 181.570 ;
        RECT 92.165 181.385 92.455 181.430 ;
        RECT 96.750 181.370 97.070 181.430 ;
        RECT 109.185 181.570 109.475 181.615 ;
        RECT 109.630 181.570 109.950 181.630 ;
        RECT 109.185 181.430 109.950 181.570 ;
        RECT 109.185 181.385 109.475 181.430 ;
        RECT 109.630 181.370 109.950 181.430 ;
        RECT 116.990 181.570 117.310 181.630 ;
        RECT 122.970 181.570 123.290 181.630 ;
        RECT 116.990 181.430 123.290 181.570 ;
        RECT 116.990 181.370 117.310 181.430 ;
        RECT 122.970 181.370 123.290 181.430 ;
        RECT 11.120 180.750 150.500 181.230 ;
        RECT 20.390 180.350 20.710 180.610 ;
        RECT 35.585 180.550 35.875 180.595 ;
        RECT 42.930 180.550 43.250 180.610 ;
        RECT 49.830 180.550 50.150 180.610 ;
        RECT 51.225 180.550 51.515 180.595 ;
        RECT 54.890 180.550 55.210 180.610 ;
        RECT 35.585 180.410 45.920 180.550 ;
        RECT 35.585 180.365 35.875 180.410 ;
        RECT 42.930 180.350 43.250 180.410 ;
        RECT 13.990 180.210 14.280 180.255 ;
        RECT 16.090 180.210 16.380 180.255 ;
        RECT 17.660 180.210 17.950 180.255 ;
        RECT 13.990 180.070 17.950 180.210 ;
        RECT 13.990 180.025 14.280 180.070 ;
        RECT 16.090 180.025 16.380 180.070 ;
        RECT 17.660 180.025 17.950 180.070 ;
        RECT 23.625 180.025 23.915 180.255 ;
        RECT 25.030 180.210 25.320 180.255 ;
        RECT 27.130 180.210 27.420 180.255 ;
        RECT 28.700 180.210 28.990 180.255 ;
        RECT 25.030 180.070 28.990 180.210 ;
        RECT 25.030 180.025 25.320 180.070 ;
        RECT 27.130 180.025 27.420 180.070 ;
        RECT 28.700 180.025 28.990 180.070 ;
        RECT 34.190 180.210 34.510 180.270 ;
        RECT 35.110 180.210 35.430 180.270 ;
        RECT 34.190 180.070 35.430 180.210 ;
        RECT 14.385 179.870 14.675 179.915 ;
        RECT 15.575 179.870 15.865 179.915 ;
        RECT 18.095 179.870 18.385 179.915 ;
        RECT 14.385 179.730 18.385 179.870 ;
        RECT 14.385 179.685 14.675 179.730 ;
        RECT 15.575 179.685 15.865 179.730 ;
        RECT 18.095 179.685 18.385 179.730 ;
        RECT 13.505 179.530 13.795 179.575 ;
        RECT 13.950 179.530 14.270 179.590 ;
        RECT 13.505 179.390 14.270 179.530 ;
        RECT 13.505 179.345 13.795 179.390 ;
        RECT 13.950 179.330 14.270 179.390 ;
        RECT 14.840 179.530 15.130 179.575 ;
        RECT 17.170 179.530 17.490 179.590 ;
        RECT 14.840 179.390 17.490 179.530 ;
        RECT 14.840 179.345 15.130 179.390 ;
        RECT 17.170 179.330 17.490 179.390 ;
        RECT 22.245 179.530 22.535 179.575 ;
        RECT 23.700 179.530 23.840 180.025 ;
        RECT 34.190 180.010 34.510 180.070 ;
        RECT 35.110 180.010 35.430 180.070 ;
        RECT 36.530 180.210 36.820 180.255 ;
        RECT 38.630 180.210 38.920 180.255 ;
        RECT 40.200 180.210 40.490 180.255 ;
        RECT 36.530 180.070 40.490 180.210 ;
        RECT 36.530 180.025 36.820 180.070 ;
        RECT 38.630 180.025 38.920 180.070 ;
        RECT 40.200 180.025 40.490 180.070 ;
        RECT 25.425 179.870 25.715 179.915 ;
        RECT 26.615 179.870 26.905 179.915 ;
        RECT 29.135 179.870 29.425 179.915 ;
        RECT 36.030 179.870 36.350 179.930 ;
        RECT 25.425 179.730 29.425 179.870 ;
        RECT 25.425 179.685 25.715 179.730 ;
        RECT 26.615 179.685 26.905 179.730 ;
        RECT 29.135 179.685 29.425 179.730 ;
        RECT 32.900 179.730 36.350 179.870 ;
        RECT 24.545 179.530 24.835 179.575 ;
        RECT 32.900 179.530 33.040 179.730 ;
        RECT 36.030 179.670 36.350 179.730 ;
        RECT 36.925 179.870 37.215 179.915 ;
        RECT 38.115 179.870 38.405 179.915 ;
        RECT 40.635 179.870 40.925 179.915 ;
        RECT 36.925 179.730 40.925 179.870 ;
        RECT 36.925 179.685 37.215 179.730 ;
        RECT 38.115 179.685 38.405 179.730 ;
        RECT 40.635 179.685 40.925 179.730 ;
        RECT 43.480 179.730 44.540 179.870 ;
        RECT 43.480 179.590 43.620 179.730 ;
        RECT 22.245 179.390 23.380 179.530 ;
        RECT 23.700 179.390 24.300 179.530 ;
        RECT 22.245 179.345 22.535 179.390 ;
        RECT 22.690 178.650 23.010 178.910 ;
        RECT 23.240 178.850 23.380 179.390 ;
        RECT 23.610 178.990 23.930 179.250 ;
        RECT 24.160 179.190 24.300 179.390 ;
        RECT 24.545 179.390 33.040 179.530 ;
        RECT 33.285 179.530 33.575 179.575 ;
        RECT 34.665 179.530 34.955 179.575 ;
        RECT 33.285 179.390 34.955 179.530 ;
        RECT 24.545 179.345 24.835 179.390 ;
        RECT 33.285 179.345 33.575 179.390 ;
        RECT 34.665 179.345 34.955 179.390 ;
        RECT 35.110 179.530 35.430 179.590 ;
        RECT 35.585 179.530 35.875 179.575 ;
        RECT 35.110 179.390 35.875 179.530 ;
        RECT 25.770 179.190 26.060 179.235 ;
        RECT 33.360 179.190 33.500 179.345 ;
        RECT 35.110 179.330 35.430 179.390 ;
        RECT 35.585 179.345 35.875 179.390 ;
        RECT 43.390 179.330 43.710 179.590 ;
        RECT 43.850 179.330 44.170 179.590 ;
        RECT 44.400 179.575 44.540 179.730 ;
        RECT 45.780 179.575 45.920 180.410 ;
        RECT 49.830 180.410 51.515 180.550 ;
        RECT 49.830 180.350 50.150 180.410 ;
        RECT 51.225 180.365 51.515 180.410 ;
        RECT 52.680 180.410 55.210 180.550 ;
        RECT 50.305 180.210 50.595 180.255 ;
        RECT 52.680 180.210 52.820 180.410 ;
        RECT 54.890 180.350 55.210 180.410 ;
        RECT 55.365 180.550 55.655 180.595 ;
        RECT 56.270 180.550 56.590 180.610 ;
        RECT 55.365 180.410 56.590 180.550 ;
        RECT 55.365 180.365 55.655 180.410 ;
        RECT 56.270 180.350 56.590 180.410 ;
        RECT 78.350 180.550 78.670 180.610 ;
        RECT 79.285 180.550 79.575 180.595 ;
        RECT 86.630 180.550 86.950 180.610 ;
        RECT 78.350 180.410 79.575 180.550 ;
        RECT 78.350 180.350 78.670 180.410 ;
        RECT 79.285 180.365 79.575 180.410 ;
        RECT 80.280 180.410 86.950 180.550 ;
        RECT 50.305 180.070 52.820 180.210 ;
        RECT 53.140 180.070 67.080 180.210 ;
        RECT 50.305 180.025 50.595 180.070 ;
        RECT 48.450 179.670 48.770 179.930 ;
        RECT 44.325 179.345 44.615 179.575 ;
        RECT 45.705 179.345 45.995 179.575 ;
        RECT 47.070 179.330 47.390 179.590 ;
        RECT 47.545 179.345 47.835 179.575 ;
        RECT 48.540 179.530 48.680 179.670 ;
        RECT 50.290 179.530 50.610 179.590 ;
        RECT 51.225 179.530 51.515 179.575 ;
        RECT 48.540 179.390 51.515 179.530 ;
        RECT 37.410 179.235 37.730 179.250 ;
        RECT 24.160 179.050 26.060 179.190 ;
        RECT 25.770 179.005 26.060 179.050 ;
        RECT 31.520 179.050 33.500 179.190 ;
        RECT 24.990 178.850 25.310 178.910 ;
        RECT 31.520 178.895 31.660 179.050 ;
        RECT 37.380 179.005 37.730 179.235 ;
        RECT 37.410 178.990 37.730 179.005 ;
        RECT 23.240 178.710 25.310 178.850 ;
        RECT 24.990 178.650 25.310 178.710 ;
        RECT 31.445 178.665 31.735 178.895 ;
        RECT 32.350 178.650 32.670 178.910 ;
        RECT 42.010 178.850 42.330 178.910 ;
        RECT 42.945 178.850 43.235 178.895 ;
        RECT 47.620 178.850 47.760 179.345 ;
        RECT 50.290 179.330 50.610 179.390 ;
        RECT 51.225 179.345 51.515 179.390 ;
        RECT 51.670 179.330 51.990 179.590 ;
        RECT 53.140 179.575 53.280 180.070 ;
        RECT 54.890 179.870 55.210 179.930 ;
        RECT 57.650 179.870 57.970 179.930 ;
        RECT 54.890 179.730 57.420 179.870 ;
        RECT 54.890 179.670 55.210 179.730 ;
        RECT 53.065 179.345 53.355 179.575 ;
        RECT 53.510 179.530 53.830 179.590 ;
        RECT 56.055 179.530 56.345 179.575 ;
        RECT 53.510 179.390 56.345 179.530 ;
        RECT 57.280 179.530 57.420 179.730 ;
        RECT 57.650 179.730 58.340 179.870 ;
        RECT 57.650 179.670 57.970 179.730 ;
        RECT 58.200 179.575 58.340 179.730 ;
        RECT 57.280 179.390 57.880 179.530 ;
        RECT 53.510 179.330 53.830 179.390 ;
        RECT 56.055 179.345 56.345 179.390 ;
        RECT 51.760 179.190 51.900 179.330 ;
        RECT 56.745 179.190 57.035 179.235 ;
        RECT 51.760 179.050 57.035 179.190 ;
        RECT 56.360 178.910 56.500 179.050 ;
        RECT 56.745 179.005 57.035 179.050 ;
        RECT 57.205 179.005 57.495 179.235 ;
        RECT 57.740 179.190 57.880 179.390 ;
        RECT 58.120 179.345 58.410 179.575 ;
        RECT 58.570 179.330 58.890 179.590 ;
        RECT 59.965 179.530 60.255 179.575 ;
        RECT 59.120 179.390 60.255 179.530 ;
        RECT 59.120 179.190 59.260 179.390 ;
        RECT 59.965 179.345 60.255 179.390 ;
        RECT 60.870 179.330 61.190 179.590 ;
        RECT 57.740 179.050 59.260 179.190 ;
        RECT 59.490 179.190 59.810 179.250 ;
        RECT 60.425 179.190 60.715 179.235 ;
        RECT 59.490 179.050 60.715 179.190 ;
        RECT 42.010 178.710 47.760 178.850 ;
        RECT 42.010 178.650 42.330 178.710 ;
        RECT 42.945 178.665 43.235 178.710 ;
        RECT 56.270 178.650 56.590 178.910 ;
        RECT 57.280 178.850 57.420 179.005 ;
        RECT 59.490 178.990 59.810 179.050 ;
        RECT 60.425 179.005 60.715 179.050 ;
        RECT 59.950 178.850 60.270 178.910 ;
        RECT 57.280 178.710 60.270 178.850 ;
        RECT 60.960 178.850 61.100 179.330 ;
        RECT 66.940 179.190 67.080 180.070 ;
        RECT 67.770 180.010 68.090 180.270 ;
        RECT 68.690 179.870 69.010 179.930 ;
        RECT 80.280 179.915 80.420 180.410 ;
        RECT 86.630 180.350 86.950 180.410 ;
        RECT 87.550 180.550 87.870 180.610 ;
        RECT 89.405 180.550 89.695 180.595 ;
        RECT 94.450 180.550 94.770 180.610 ;
        RECT 87.550 180.410 89.695 180.550 ;
        RECT 87.550 180.350 87.870 180.410 ;
        RECT 89.405 180.365 89.695 180.410 ;
        RECT 89.940 180.410 94.770 180.550 ;
        RECT 80.690 180.210 80.980 180.255 ;
        RECT 82.790 180.210 83.080 180.255 ;
        RECT 84.360 180.210 84.650 180.255 ;
        RECT 89.940 180.210 90.080 180.410 ;
        RECT 94.450 180.350 94.770 180.410 ;
        RECT 102.730 180.550 103.050 180.610 ;
        RECT 104.125 180.550 104.415 180.595 ;
        RECT 102.730 180.410 104.415 180.550 ;
        RECT 102.730 180.350 103.050 180.410 ;
        RECT 104.125 180.365 104.415 180.410 ;
        RECT 113.770 180.550 114.090 180.610 ;
        RECT 114.705 180.550 114.995 180.595 ;
        RECT 113.770 180.410 114.995 180.550 ;
        RECT 113.770 180.350 114.090 180.410 ;
        RECT 114.705 180.365 114.995 180.410 ;
        RECT 118.385 180.550 118.675 180.595 ;
        RECT 122.050 180.550 122.370 180.610 ;
        RECT 118.385 180.410 122.370 180.550 ;
        RECT 118.385 180.365 118.675 180.410 ;
        RECT 122.050 180.350 122.370 180.410 ;
        RECT 122.510 180.550 122.830 180.610 ;
        RECT 124.365 180.550 124.655 180.595 ;
        RECT 122.510 180.410 129.135 180.550 ;
        RECT 122.510 180.350 122.830 180.410 ;
        RECT 124.365 180.365 124.655 180.410 ;
        RECT 80.690 180.070 84.650 180.210 ;
        RECT 80.690 180.025 80.980 180.070 ;
        RECT 82.790 180.025 83.080 180.070 ;
        RECT 84.360 180.025 84.650 180.070 ;
        RECT 87.180 180.070 90.080 180.210 ;
        RECT 90.325 180.210 90.615 180.255 ;
        RECT 95.385 180.210 95.675 180.255 ;
        RECT 90.325 180.070 95.675 180.210 ;
        RECT 67.400 179.730 79.960 179.870 ;
        RECT 67.400 179.575 67.540 179.730 ;
        RECT 68.690 179.670 69.010 179.730 ;
        RECT 67.325 179.345 67.615 179.575 ;
        RECT 68.245 179.530 68.535 179.575 ;
        RECT 71.910 179.530 72.230 179.590 ;
        RECT 78.365 179.530 78.655 179.575 ;
        RECT 68.245 179.390 70.530 179.530 ;
        RECT 68.245 179.345 68.535 179.390 ;
        RECT 70.390 179.190 70.530 179.390 ;
        RECT 71.910 179.390 78.655 179.530 ;
        RECT 71.910 179.330 72.230 179.390 ;
        RECT 78.365 179.345 78.655 179.390 ;
        RECT 79.285 179.345 79.575 179.575 ;
        RECT 79.820 179.530 79.960 179.730 ;
        RECT 80.205 179.685 80.495 179.915 ;
        RECT 81.085 179.870 81.375 179.915 ;
        RECT 82.275 179.870 82.565 179.915 ;
        RECT 84.795 179.870 85.085 179.915 ;
        RECT 81.085 179.730 85.085 179.870 ;
        RECT 81.085 179.685 81.375 179.730 ;
        RECT 82.275 179.685 82.565 179.730 ;
        RECT 84.795 179.685 85.085 179.730 ;
        RECT 83.410 179.530 83.730 179.590 ;
        RECT 79.820 179.390 83.730 179.530 ;
        RECT 78.810 179.190 79.130 179.250 ;
        RECT 79.360 179.190 79.500 179.345 ;
        RECT 83.410 179.330 83.730 179.390 ;
        RECT 66.940 179.050 69.840 179.190 ;
        RECT 70.390 179.050 79.500 179.190 ;
        RECT 81.540 179.190 81.830 179.235 ;
        RECT 82.490 179.190 82.810 179.250 ;
        RECT 81.540 179.050 82.810 179.190 ;
        RECT 67.310 178.850 67.630 178.910 ;
        RECT 60.960 178.710 67.630 178.850 ;
        RECT 69.700 178.850 69.840 179.050 ;
        RECT 78.810 178.990 79.130 179.050 ;
        RECT 81.540 179.005 81.830 179.050 ;
        RECT 82.490 178.990 82.810 179.050 ;
        RECT 87.180 178.895 87.320 180.070 ;
        RECT 90.325 180.025 90.615 180.070 ;
        RECT 95.385 180.025 95.675 180.070 ;
        RECT 119.750 180.210 120.070 180.270 ;
        RECT 128.505 180.210 128.795 180.255 ;
        RECT 119.750 180.070 128.795 180.210 ;
        RECT 119.750 180.010 120.070 180.070 ;
        RECT 96.750 179.670 97.070 179.930 ;
        RECT 111.930 179.870 112.250 179.930 ;
        RECT 112.865 179.870 113.155 179.915 ;
        RECT 120.225 179.870 120.515 179.915 ;
        RECT 121.590 179.870 121.910 179.930 ;
        RECT 99.600 179.730 105.260 179.870 ;
        RECT 88.945 179.345 89.235 179.575 ;
        RECT 89.020 179.190 89.160 179.345 ;
        RECT 89.850 179.330 90.170 179.590 ;
        RECT 91.320 179.575 92.255 179.610 ;
        RECT 91.245 179.510 92.255 179.575 ;
        RECT 91.245 179.470 92.380 179.510 ;
        RECT 91.245 179.345 91.535 179.470 ;
        RECT 92.115 179.370 92.380 179.470 ;
        RECT 89.020 179.050 91.120 179.190 ;
        RECT 87.105 178.850 87.395 178.895 ;
        RECT 69.700 178.710 87.395 178.850 ;
        RECT 59.950 178.650 60.270 178.710 ;
        RECT 67.310 178.650 67.630 178.710 ;
        RECT 87.105 178.665 87.395 178.710 ;
        RECT 87.550 178.650 87.870 178.910 ;
        RECT 90.980 178.850 91.120 179.050 ;
        RECT 91.705 179.005 91.995 179.235 ;
        RECT 92.240 179.190 92.380 179.370 ;
        RECT 94.450 179.330 94.770 179.590 ;
        RECT 96.290 179.330 96.610 179.590 ;
        RECT 97.225 179.345 97.515 179.575 ;
        RECT 96.380 179.190 96.520 179.330 ;
        RECT 92.240 179.050 96.520 179.190 ;
        RECT 97.300 179.190 97.440 179.345 ;
        RECT 98.590 179.330 98.910 179.590 ;
        RECT 99.600 179.575 99.740 179.730 ;
        RECT 105.120 179.590 105.260 179.730 ;
        RECT 111.930 179.730 115.840 179.870 ;
        RECT 111.930 179.670 112.250 179.730 ;
        RECT 112.865 179.685 113.155 179.730 ;
        RECT 99.525 179.345 99.815 179.575 ;
        RECT 103.190 179.330 103.510 179.590 ;
        RECT 105.030 179.330 105.350 179.590 ;
        RECT 110.090 179.530 110.410 179.590 ;
        RECT 112.405 179.530 112.695 179.575 ;
        RECT 105.580 179.390 112.695 179.530 ;
        RECT 99.065 179.190 99.355 179.235 ;
        RECT 97.300 179.050 99.355 179.190 ;
        RECT 99.065 179.005 99.355 179.050 ;
        RECT 91.780 178.850 91.920 179.005 ;
        RECT 90.980 178.710 91.920 178.850 ;
        RECT 92.150 178.850 92.470 178.910 ;
        RECT 105.580 178.850 105.720 179.390 ;
        RECT 110.090 179.330 110.410 179.390 ;
        RECT 112.405 179.345 112.695 179.390 ;
        RECT 113.310 179.530 113.630 179.590 ;
        RECT 113.785 179.530 114.075 179.575 ;
        RECT 113.310 179.390 114.075 179.530 ;
        RECT 106.870 179.190 107.190 179.250 ;
        RECT 108.250 179.190 108.570 179.250 ;
        RECT 112.480 179.190 112.620 179.345 ;
        RECT 113.310 179.330 113.630 179.390 ;
        RECT 113.785 179.345 114.075 179.390 ;
        RECT 115.165 179.345 115.455 179.575 ;
        RECT 115.700 179.530 115.840 179.730 ;
        RECT 120.225 179.730 121.910 179.870 ;
        RECT 120.225 179.685 120.515 179.730 ;
        RECT 121.590 179.670 121.910 179.730 ;
        RECT 122.970 179.870 123.290 179.930 ;
        RECT 124.825 179.870 125.115 179.915 ;
        RECT 122.970 179.730 125.115 179.870 ;
        RECT 122.970 179.670 123.290 179.730 ;
        RECT 124.825 179.685 125.115 179.730 ;
        RECT 116.085 179.530 116.375 179.575 ;
        RECT 116.530 179.530 116.850 179.590 ;
        RECT 115.700 179.390 116.850 179.530 ;
        RECT 116.085 179.345 116.375 179.390 ;
        RECT 115.240 179.190 115.380 179.345 ;
        RECT 116.530 179.330 116.850 179.390 ;
        RECT 119.290 179.330 119.610 179.590 ;
        RECT 106.870 179.050 110.320 179.190 ;
        RECT 112.480 179.050 115.380 179.190 ;
        RECT 124.900 179.190 125.040 179.685 ;
        RECT 125.360 179.575 125.500 180.070 ;
        RECT 128.505 180.025 128.795 180.070 ;
        RECT 127.585 179.870 127.875 179.915 ;
        RECT 128.995 179.870 129.135 180.410 ;
        RECT 129.870 179.870 130.190 179.930 ;
        RECT 127.585 179.730 130.190 179.870 ;
        RECT 127.585 179.685 127.875 179.730 ;
        RECT 129.870 179.670 130.190 179.730 ;
        RECT 125.285 179.345 125.575 179.575 ;
        RECT 128.965 179.530 129.255 179.575 ;
        RECT 134.470 179.530 134.790 179.590 ;
        RECT 128.965 179.390 134.790 179.530 ;
        RECT 128.965 179.345 129.255 179.390 ;
        RECT 129.040 179.190 129.180 179.345 ;
        RECT 134.470 179.330 134.790 179.390 ;
        RECT 124.900 179.050 129.180 179.190 ;
        RECT 106.870 178.990 107.190 179.050 ;
        RECT 108.250 178.990 108.570 179.050 ;
        RECT 92.150 178.710 105.720 178.850 ;
        RECT 105.950 178.850 106.270 178.910 ;
        RECT 109.630 178.850 109.950 178.910 ;
        RECT 105.950 178.710 109.950 178.850 ;
        RECT 110.180 178.850 110.320 179.050 ;
        RECT 116.545 178.850 116.835 178.895 ;
        RECT 117.910 178.850 118.230 178.910 ;
        RECT 110.180 178.710 118.230 178.850 ;
        RECT 92.150 178.650 92.470 178.710 ;
        RECT 105.950 178.650 106.270 178.710 ;
        RECT 109.630 178.650 109.950 178.710 ;
        RECT 116.545 178.665 116.835 178.710 ;
        RECT 117.910 178.650 118.230 178.710 ;
        RECT 123.430 178.650 123.750 178.910 ;
        RECT 127.570 178.650 127.890 178.910 ;
        RECT 11.120 178.030 151.295 178.510 ;
        RECT 17.185 177.830 17.475 177.875 ;
        RECT 17.630 177.830 17.950 177.890 ;
        RECT 17.185 177.690 17.950 177.830 ;
        RECT 17.185 177.645 17.475 177.690 ;
        RECT 17.630 177.630 17.950 177.690 ;
        RECT 23.610 177.830 23.930 177.890 ;
        RECT 24.545 177.830 24.835 177.875 ;
        RECT 23.610 177.690 24.835 177.830 ;
        RECT 23.610 177.630 23.930 177.690 ;
        RECT 24.545 177.645 24.835 177.690 ;
        RECT 34.650 177.830 34.970 177.890 ;
        RECT 36.030 177.830 36.350 177.890 ;
        RECT 53.985 177.830 54.275 177.875 ;
        RECT 55.810 177.830 56.130 177.890 ;
        RECT 57.190 177.830 57.510 177.890 ;
        RECT 34.650 177.690 35.340 177.830 ;
        RECT 34.650 177.630 34.970 177.690 ;
        RECT 35.200 177.490 35.340 177.690 ;
        RECT 36.030 177.690 57.510 177.830 ;
        RECT 36.030 177.630 36.350 177.690 ;
        RECT 53.985 177.645 54.275 177.690 ;
        RECT 55.810 177.630 56.130 177.690 ;
        RECT 57.190 177.630 57.510 177.690 ;
        RECT 59.950 177.830 60.270 177.890 ;
        RECT 70.990 177.830 71.310 177.890 ;
        RECT 59.950 177.690 71.310 177.830 ;
        RECT 59.950 177.630 60.270 177.690 ;
        RECT 33.360 177.350 35.340 177.490 ;
        RECT 33.360 177.210 33.500 177.350 ;
        RECT 16.710 177.150 17.030 177.210 ;
        RECT 16.710 177.010 17.400 177.150 ;
        RECT 16.710 176.950 17.030 177.010 ;
        RECT 17.260 176.855 17.400 177.010 ;
        RECT 18.550 176.950 18.870 177.210 ;
        RECT 22.690 177.150 23.010 177.210 ;
        RECT 25.925 177.150 26.215 177.195 ;
        RECT 32.350 177.150 32.670 177.210 ;
        RECT 22.690 177.010 32.670 177.150 ;
        RECT 22.690 176.950 23.010 177.010 ;
        RECT 25.925 176.965 26.215 177.010 ;
        RECT 32.350 176.950 32.670 177.010 ;
        RECT 33.270 176.950 33.590 177.210 ;
        RECT 35.200 177.195 35.340 177.350 ;
        RECT 56.730 177.290 57.050 177.550 ;
        RECT 60.500 177.535 60.640 177.690 ;
        RECT 70.990 177.630 71.310 177.690 ;
        RECT 76.050 177.830 76.370 177.890 ;
        RECT 76.050 177.690 80.420 177.830 ;
        RECT 76.050 177.630 76.370 177.690 ;
        RECT 60.425 177.305 60.715 177.535 ;
        RECT 64.105 177.490 64.395 177.535 ;
        RECT 65.930 177.490 66.250 177.550 ;
        RECT 64.105 177.350 66.250 177.490 ;
        RECT 64.105 177.305 64.395 177.350 ;
        RECT 65.930 177.290 66.250 177.350 ;
        RECT 68.230 177.290 68.550 177.550 ;
        RECT 77.890 177.490 78.210 177.550 ;
        RECT 71.080 177.350 78.210 177.490 ;
        RECT 34.665 176.965 34.955 177.195 ;
        RECT 35.125 176.965 35.415 177.195 ;
        RECT 35.570 177.150 35.890 177.210 ;
        RECT 37.425 177.150 37.715 177.195 ;
        RECT 39.710 177.150 40.030 177.210 ;
        RECT 35.570 177.010 40.030 177.150 ;
        RECT 17.185 176.810 17.475 176.855 ;
        RECT 24.545 176.810 24.835 176.855 ;
        RECT 17.185 176.670 24.835 176.810 ;
        RECT 17.185 176.625 17.475 176.670 ;
        RECT 24.545 176.625 24.835 176.670 ;
        RECT 33.730 176.810 34.050 176.870 ;
        RECT 34.205 176.810 34.495 176.855 ;
        RECT 34.740 176.810 34.880 176.965 ;
        RECT 35.570 176.950 35.890 177.010 ;
        RECT 37.425 176.965 37.715 177.010 ;
        RECT 39.710 176.950 40.030 177.010 ;
        RECT 46.165 177.150 46.455 177.195 ;
        RECT 47.545 177.150 47.835 177.195 ;
        RECT 49.370 177.150 49.690 177.210 ;
        RECT 46.165 177.010 49.690 177.150 ;
        RECT 46.165 176.965 46.455 177.010 ;
        RECT 47.545 176.965 47.835 177.010 ;
        RECT 49.370 176.950 49.690 177.010 ;
        RECT 59.490 177.150 59.810 177.210 ;
        RECT 71.080 177.195 71.220 177.350 ;
        RECT 77.890 177.290 78.210 177.350 ;
        RECT 78.900 177.350 79.960 177.490 ;
        RECT 72.370 177.195 72.690 177.210 ;
        RECT 67.325 177.150 67.615 177.195 ;
        RECT 59.490 177.010 67.615 177.150 ;
        RECT 59.490 176.950 59.810 177.010 ;
        RECT 67.325 176.965 67.615 177.010 ;
        RECT 68.705 176.965 68.995 177.195 ;
        RECT 71.005 176.965 71.295 177.195 ;
        RECT 72.340 177.150 72.690 177.195 ;
        RECT 78.900 177.150 79.040 177.350 ;
        RECT 72.175 177.010 72.690 177.150 ;
        RECT 72.340 176.965 72.690 177.010 ;
        RECT 33.730 176.670 34.880 176.810 ;
        RECT 36.030 176.810 36.350 176.870 ;
        RECT 36.030 176.670 39.020 176.810 ;
        RECT 15.790 176.130 16.110 176.190 ;
        RECT 18.105 176.130 18.395 176.175 ;
        RECT 15.790 175.990 18.395 176.130 ;
        RECT 24.620 176.130 24.760 176.625 ;
        RECT 33.730 176.610 34.050 176.670 ;
        RECT 34.205 176.625 34.495 176.670 ;
        RECT 36.030 176.610 36.350 176.670 ;
        RECT 38.880 176.530 39.020 176.670 ;
        RECT 57.650 176.610 57.970 176.870 ;
        RECT 58.110 176.610 58.430 176.870 ;
        RECT 58.570 176.810 58.890 176.870 ;
        RECT 66.850 176.810 67.170 176.870 ;
        RECT 58.570 176.670 67.170 176.810 ;
        RECT 58.570 176.610 58.890 176.670 ;
        RECT 24.990 176.470 25.310 176.530 ;
        RECT 25.465 176.470 25.755 176.515 ;
        RECT 32.365 176.470 32.655 176.515 ;
        RECT 24.990 176.330 38.560 176.470 ;
        RECT 24.990 176.270 25.310 176.330 ;
        RECT 25.465 176.285 25.755 176.330 ;
        RECT 32.365 176.285 32.655 176.330 ;
        RECT 38.420 176.190 38.560 176.330 ;
        RECT 38.790 176.270 39.110 176.530 ;
        RECT 60.500 176.515 60.640 176.670 ;
        RECT 66.850 176.610 67.170 176.670 ;
        RECT 68.230 176.810 68.550 176.870 ;
        RECT 68.780 176.810 68.920 176.965 ;
        RECT 72.370 176.950 72.690 176.965 ;
        RECT 77.520 177.010 79.040 177.150 ;
        RECT 68.230 176.670 68.920 176.810 ;
        RECT 71.885 176.810 72.175 176.855 ;
        RECT 73.075 176.810 73.365 176.855 ;
        RECT 75.595 176.810 75.885 176.855 ;
        RECT 71.885 176.670 75.885 176.810 ;
        RECT 68.230 176.610 68.550 176.670 ;
        RECT 71.885 176.625 72.175 176.670 ;
        RECT 73.075 176.625 73.365 176.670 ;
        RECT 75.595 176.625 75.885 176.670 ;
        RECT 60.425 176.285 60.715 176.515 ;
        RECT 63.185 176.470 63.475 176.515 ;
        RECT 64.550 176.470 64.870 176.530 ;
        RECT 63.185 176.330 64.870 176.470 ;
        RECT 63.185 176.285 63.475 176.330 ;
        RECT 64.550 176.270 64.870 176.330 ;
        RECT 65.945 176.470 66.235 176.515 ;
        RECT 71.490 176.470 71.780 176.515 ;
        RECT 73.590 176.470 73.880 176.515 ;
        RECT 75.160 176.470 75.450 176.515 ;
        RECT 65.945 176.330 70.530 176.470 ;
        RECT 65.945 176.285 66.235 176.330 ;
        RECT 26.830 176.130 27.150 176.190 ;
        RECT 24.620 175.990 27.150 176.130 ;
        RECT 15.790 175.930 16.110 175.990 ;
        RECT 18.105 175.945 18.395 175.990 ;
        RECT 26.830 175.930 27.150 175.990 ;
        RECT 35.585 176.130 35.875 176.175 ;
        RECT 36.490 176.130 36.810 176.190 ;
        RECT 35.585 175.990 36.810 176.130 ;
        RECT 35.585 175.945 35.875 175.990 ;
        RECT 36.490 175.930 36.810 175.990 ;
        RECT 38.330 175.930 38.650 176.190 ;
        RECT 64.105 176.130 64.395 176.175 ;
        RECT 66.405 176.130 66.695 176.175 ;
        RECT 64.105 175.990 66.695 176.130 ;
        RECT 70.390 176.130 70.530 176.330 ;
        RECT 71.490 176.330 75.450 176.470 ;
        RECT 71.490 176.285 71.780 176.330 ;
        RECT 73.590 176.285 73.880 176.330 ;
        RECT 75.160 176.285 75.450 176.330 ;
        RECT 77.520 176.130 77.660 177.010 ;
        RECT 79.270 176.950 79.590 177.210 ;
        RECT 77.905 176.470 78.195 176.515 ;
        RECT 79.360 176.470 79.500 176.950 ;
        RECT 79.820 176.810 79.960 177.350 ;
        RECT 80.280 177.195 80.420 177.690 ;
        RECT 82.490 177.630 82.810 177.890 ;
        RECT 87.550 177.630 87.870 177.890 ;
        RECT 90.770 177.830 91.090 177.890 ;
        RECT 102.285 177.830 102.575 177.875 ;
        RECT 103.190 177.830 103.510 177.890 ;
        RECT 90.770 177.690 102.040 177.830 ;
        RECT 90.770 177.630 91.090 177.690 ;
        RECT 80.205 176.965 80.495 177.195 ;
        RECT 83.410 176.950 83.730 177.210 ;
        RECT 84.345 177.150 84.635 177.195 ;
        RECT 87.640 177.150 87.780 177.630 ;
        RECT 92.040 177.490 92.330 177.535 ;
        RECT 95.385 177.490 95.675 177.535 ;
        RECT 92.040 177.350 95.675 177.490 ;
        RECT 92.040 177.305 92.330 177.350 ;
        RECT 95.385 177.305 95.675 177.350 ;
        RECT 95.920 177.350 96.980 177.490 ;
        RECT 84.345 177.010 87.780 177.150 ;
        RECT 93.990 177.150 94.310 177.210 ;
        RECT 95.920 177.195 96.060 177.350 ;
        RECT 96.840 177.210 96.980 177.350 ;
        RECT 94.925 177.150 95.215 177.195 ;
        RECT 93.990 177.010 95.215 177.150 ;
        RECT 84.345 176.965 84.635 177.010 ;
        RECT 93.990 176.950 94.310 177.010 ;
        RECT 94.925 176.965 95.215 177.010 ;
        RECT 95.845 176.965 96.135 177.195 ;
        RECT 96.290 176.950 96.610 177.210 ;
        RECT 96.750 176.950 97.070 177.210 ;
        RECT 101.900 177.150 102.040 177.690 ;
        RECT 102.285 177.690 103.510 177.830 ;
        RECT 102.285 177.645 102.575 177.690 ;
        RECT 103.190 177.630 103.510 177.690 ;
        RECT 104.585 177.645 104.875 177.875 ;
        RECT 104.660 177.490 104.800 177.645 ;
        RECT 112.390 177.630 112.710 177.890 ;
        RECT 122.050 177.630 122.370 177.890 ;
        RECT 127.570 177.630 127.890 177.890 ;
        RECT 105.505 177.490 105.795 177.535 ;
        RECT 105.950 177.490 106.270 177.550 ;
        RECT 107.805 177.490 108.095 177.535 ;
        RECT 104.660 177.350 105.260 177.490 ;
        RECT 104.125 177.150 104.415 177.195 ;
        RECT 101.900 177.010 104.415 177.150 ;
        RECT 105.120 177.150 105.260 177.350 ;
        RECT 105.505 177.350 108.095 177.490 ;
        RECT 105.505 177.305 105.795 177.350 ;
        RECT 105.950 177.290 106.270 177.350 ;
        RECT 107.805 177.305 108.095 177.350 ;
        RECT 108.250 177.490 108.570 177.550 ;
        RECT 112.480 177.490 112.620 177.630 ;
        RECT 116.990 177.490 117.310 177.550 ;
        RECT 122.510 177.490 122.830 177.550 ;
        RECT 108.250 177.350 108.765 177.490 ;
        RECT 112.480 177.350 122.830 177.490 ;
        RECT 108.250 177.290 108.570 177.350 ;
        RECT 116.990 177.290 117.310 177.350 ;
        RECT 106.870 177.180 107.190 177.210 ;
        RECT 108.710 177.195 109.030 177.210 ;
        RECT 106.500 177.150 107.190 177.180 ;
        RECT 105.120 177.040 107.190 177.150 ;
        RECT 105.120 177.010 106.640 177.040 ;
        RECT 104.125 176.965 104.415 177.010 ;
        RECT 84.805 176.810 85.095 176.855 ;
        RECT 92.150 176.810 92.470 176.870 ;
        RECT 92.625 176.810 92.915 176.855 ;
        RECT 79.820 176.670 91.460 176.810 ;
        RECT 84.805 176.625 85.095 176.670 ;
        RECT 91.320 176.515 91.460 176.670 ;
        RECT 92.150 176.670 92.915 176.810 ;
        RECT 92.150 176.610 92.470 176.670 ;
        RECT 92.625 176.625 92.915 176.670 ;
        RECT 93.085 176.625 93.375 176.855 ;
        RECT 94.465 176.810 94.755 176.855 ;
        RECT 96.380 176.810 96.520 176.950 ;
        RECT 94.465 176.670 96.520 176.810 ;
        RECT 99.985 176.810 100.275 176.855 ;
        RECT 102.745 176.810 103.035 176.855 ;
        RECT 99.985 176.670 103.035 176.810 ;
        RECT 94.465 176.625 94.755 176.670 ;
        RECT 99.985 176.625 100.275 176.670 ;
        RECT 102.745 176.625 103.035 176.670 ;
        RECT 103.190 176.810 103.510 176.870 ;
        RECT 103.665 176.810 103.955 176.855 ;
        RECT 103.190 176.670 103.955 176.810 ;
        RECT 104.200 176.810 104.340 176.965 ;
        RECT 106.870 176.950 107.190 177.040 ;
        RECT 107.345 176.965 107.635 177.195 ;
        RECT 108.710 176.965 109.145 177.195 ;
        RECT 105.490 176.810 105.810 176.870 ;
        RECT 104.200 176.670 105.810 176.810 ;
        RECT 77.905 176.330 79.500 176.470 ;
        RECT 77.905 176.285 78.195 176.330 ;
        RECT 91.245 176.285 91.535 176.515 ;
        RECT 93.160 176.470 93.300 176.625 ;
        RECT 103.190 176.610 103.510 176.670 ;
        RECT 103.665 176.625 103.955 176.670 ;
        RECT 105.490 176.610 105.810 176.670 ;
        RECT 105.965 176.810 106.255 176.855 ;
        RECT 107.420 176.810 107.560 176.965 ;
        RECT 108.710 176.950 109.030 176.965 ;
        RECT 109.630 176.950 109.950 177.210 ;
        RECT 117.450 176.950 117.770 177.210 ;
        RECT 118.460 177.195 118.600 177.350 ;
        RECT 122.510 177.290 122.830 177.350 ;
        RECT 118.385 176.965 118.675 177.195 ;
        RECT 123.430 177.150 123.750 177.210 ;
        RECT 123.905 177.150 124.195 177.195 ;
        RECT 123.430 177.010 124.195 177.150 ;
        RECT 123.430 176.950 123.750 177.010 ;
        RECT 123.905 176.965 124.195 177.010 ;
        RECT 124.365 177.150 124.655 177.195 ;
        RECT 127.660 177.150 127.800 177.630 ;
        RECT 124.365 177.010 127.800 177.150 ;
        RECT 124.365 176.965 124.655 177.010 ;
        RECT 105.965 176.670 107.100 176.810 ;
        RECT 107.420 176.670 107.605 176.810 ;
        RECT 105.965 176.625 106.255 176.670 ;
        RECT 101.825 176.470 102.115 176.515 ;
        RECT 106.425 176.470 106.715 176.515 ;
        RECT 93.160 176.330 94.680 176.470 ;
        RECT 94.540 176.190 94.680 176.330 ;
        RECT 101.825 176.330 106.715 176.470 ;
        RECT 106.960 176.470 107.100 176.670 ;
        RECT 107.465 176.470 107.605 176.670 ;
        RECT 120.670 176.470 120.990 176.530 ;
        RECT 130.330 176.470 130.650 176.530 ;
        RECT 106.960 176.330 113.080 176.470 ;
        RECT 101.825 176.285 102.115 176.330 ;
        RECT 106.425 176.285 106.715 176.330 ;
        RECT 112.940 176.190 113.080 176.330 ;
        RECT 120.670 176.330 130.650 176.470 ;
        RECT 120.670 176.270 120.990 176.330 ;
        RECT 130.330 176.270 130.650 176.330 ;
        RECT 70.390 175.990 77.660 176.130 ;
        RECT 78.365 176.130 78.655 176.175 ;
        RECT 78.810 176.130 79.130 176.190 ;
        RECT 78.365 175.990 79.130 176.130 ;
        RECT 64.105 175.945 64.395 175.990 ;
        RECT 66.405 175.945 66.695 175.990 ;
        RECT 78.365 175.945 78.655 175.990 ;
        RECT 78.810 175.930 79.130 175.990 ;
        RECT 80.205 176.130 80.495 176.175 ;
        RECT 82.030 176.130 82.350 176.190 ;
        RECT 80.205 175.990 82.350 176.130 ;
        RECT 80.205 175.945 80.495 175.990 ;
        RECT 82.030 175.930 82.350 175.990 ;
        RECT 94.450 175.930 94.770 176.190 ;
        RECT 104.570 176.130 104.890 176.190 ;
        RECT 108.710 176.130 109.030 176.190 ;
        RECT 104.570 175.990 109.030 176.130 ;
        RECT 104.570 175.930 104.890 175.990 ;
        RECT 108.710 175.930 109.030 175.990 ;
        RECT 112.850 175.930 113.170 176.190 ;
        RECT 117.465 176.130 117.755 176.175 ;
        RECT 119.290 176.130 119.610 176.190 ;
        RECT 117.465 175.990 119.610 176.130 ;
        RECT 117.465 175.945 117.755 175.990 ;
        RECT 119.290 175.930 119.610 175.990 ;
        RECT 125.270 175.930 125.590 176.190 ;
        RECT 11.120 175.310 150.500 175.790 ;
        RECT 37.410 174.910 37.730 175.170 ;
        RECT 42.470 175.110 42.790 175.170 ;
        RECT 52.145 175.110 52.435 175.155 ;
        RECT 55.365 175.110 55.655 175.155 ;
        RECT 42.470 174.970 55.655 175.110 ;
        RECT 42.470 174.910 42.790 174.970 ;
        RECT 52.145 174.925 52.435 174.970 ;
        RECT 55.365 174.925 55.655 174.970 ;
        RECT 55.825 175.110 56.115 175.155 ;
        RECT 58.110 175.110 58.430 175.170 ;
        RECT 55.825 174.970 58.430 175.110 ;
        RECT 55.825 174.925 56.115 174.970 ;
        RECT 58.110 174.910 58.430 174.970 ;
        RECT 63.630 175.110 63.950 175.170 ;
        RECT 67.325 175.110 67.615 175.155 ;
        RECT 63.630 174.970 67.615 175.110 ;
        RECT 63.630 174.910 63.950 174.970 ;
        RECT 67.325 174.925 67.615 174.970 ;
        RECT 72.370 174.910 72.690 175.170 ;
        RECT 89.850 174.910 90.170 175.170 ;
        RECT 90.310 175.110 90.630 175.170 ;
        RECT 105.030 175.110 105.350 175.170 ;
        RECT 90.310 174.970 105.350 175.110 ;
        RECT 90.310 174.910 90.630 174.970 ;
        RECT 105.030 174.910 105.350 174.970 ;
        RECT 105.950 175.110 106.270 175.170 ;
        RECT 109.185 175.110 109.475 175.155 ;
        RECT 105.950 174.970 109.475 175.110 ;
        RECT 105.950 174.910 106.270 174.970 ;
        RECT 109.185 174.925 109.475 174.970 ;
        RECT 112.850 174.910 113.170 175.170 ;
        RECT 114.230 174.910 114.550 175.170 ;
        RECT 117.450 174.910 117.770 175.170 ;
        RECT 119.290 174.910 119.610 175.170 ;
        RECT 125.270 174.910 125.590 175.170 ;
        RECT 42.010 174.570 42.330 174.830 ;
        RECT 71.910 174.770 72.230 174.830 ;
        RECT 54.980 174.630 88.240 174.770 ;
        RECT 38.790 174.430 39.110 174.490 ;
        RECT 44.310 174.430 44.630 174.490 ;
        RECT 38.790 174.290 44.630 174.430 ;
        RECT 38.790 174.230 39.110 174.290 ;
        RECT 44.310 174.230 44.630 174.290 ;
        RECT 44.770 174.430 45.090 174.490 ;
        RECT 50.290 174.430 50.610 174.490 ;
        RECT 44.770 174.290 50.610 174.430 ;
        RECT 44.770 174.230 45.090 174.290 ;
        RECT 50.290 174.230 50.610 174.290 ;
        RECT 50.750 174.230 51.070 174.490 ;
        RECT 54.980 174.430 55.120 174.630 ;
        RECT 71.910 174.570 72.230 174.630 ;
        RECT 54.520 174.290 55.120 174.430 ;
        RECT 17.185 174.090 17.475 174.135 ;
        RECT 18.090 174.090 18.410 174.150 ;
        RECT 17.185 173.950 18.410 174.090 ;
        RECT 17.185 173.905 17.475 173.950 ;
        RECT 18.090 173.890 18.410 173.950 ;
        RECT 36.490 174.090 36.810 174.150 ;
        RECT 37.425 174.090 37.715 174.135 ;
        RECT 36.490 173.950 37.715 174.090 ;
        RECT 36.490 173.890 36.810 173.950 ;
        RECT 37.425 173.905 37.715 173.950 ;
        RECT 38.330 173.890 38.650 174.150 ;
        RECT 42.930 173.890 43.250 174.150 ;
        RECT 43.850 173.890 44.170 174.150 ;
        RECT 50.840 174.090 50.980 174.230 ;
        RECT 54.520 174.135 54.660 174.290 ;
        RECT 56.270 174.230 56.590 174.490 ;
        RECT 71.450 174.430 71.770 174.490 ;
        RECT 77.445 174.430 77.735 174.475 ;
        RECT 78.350 174.430 78.670 174.490 ;
        RECT 65.100 174.290 71.770 174.430 ;
        RECT 51.225 174.090 51.515 174.135 ;
        RECT 44.400 174.070 50.100 174.090 ;
        RECT 50.840 174.070 51.515 174.090 ;
        RECT 44.400 173.950 51.515 174.070 ;
        RECT 35.110 173.750 35.430 173.810 ;
        RECT 36.950 173.750 37.270 173.810 ;
        RECT 42.010 173.750 42.330 173.810 ;
        RECT 44.400 173.750 44.540 173.950 ;
        RECT 49.960 173.930 50.980 173.950 ;
        RECT 51.225 173.905 51.515 173.950 ;
        RECT 53.525 173.905 53.815 174.135 ;
        RECT 54.445 173.905 54.735 174.135 ;
        RECT 35.110 173.610 44.540 173.750 ;
        RECT 44.785 173.750 45.075 173.795 ;
        RECT 53.600 173.750 53.740 173.905 ;
        RECT 54.890 173.890 55.210 174.150 ;
        RECT 64.105 174.090 64.395 174.135 ;
        RECT 64.550 174.090 64.870 174.150 ;
        RECT 64.105 173.950 64.870 174.090 ;
        RECT 64.105 173.905 64.395 173.950 ;
        RECT 64.550 173.890 64.870 173.950 ;
        RECT 65.100 173.750 65.240 174.290 ;
        RECT 71.450 174.230 71.770 174.290 ;
        RECT 73.840 174.290 76.740 174.430 ;
        RECT 68.230 173.890 68.550 174.150 ;
        RECT 70.085 174.090 70.375 174.135 ;
        RECT 73.290 174.090 73.610 174.150 ;
        RECT 73.840 174.135 73.980 174.290 ;
        RECT 76.600 174.150 76.740 174.290 ;
        RECT 77.445 174.290 78.670 174.430 ;
        RECT 77.445 174.245 77.735 174.290 ;
        RECT 78.350 174.230 78.670 174.290 ;
        RECT 82.030 174.430 82.350 174.490 ;
        RECT 85.250 174.430 85.570 174.490 ;
        RECT 82.030 174.290 85.570 174.430 ;
        RECT 82.030 174.230 82.350 174.290 ;
        RECT 85.250 174.230 85.570 174.290 ;
        RECT 70.085 173.950 73.610 174.090 ;
        RECT 70.085 173.905 70.375 173.950 ;
        RECT 73.290 173.890 73.610 173.950 ;
        RECT 73.765 173.905 74.055 174.135 ;
        RECT 74.210 174.090 74.530 174.150 ;
        RECT 76.065 174.090 76.355 174.135 ;
        RECT 74.210 173.950 76.355 174.090 ;
        RECT 74.210 173.890 74.530 173.950 ;
        RECT 76.065 173.905 76.355 173.950 ;
        RECT 76.510 173.890 76.830 174.150 ;
        RECT 44.785 173.610 65.240 173.750 ;
        RECT 65.470 173.750 65.790 173.810 ;
        RECT 68.705 173.750 68.995 173.795 ;
        RECT 65.470 173.610 68.995 173.750 ;
        RECT 35.110 173.550 35.430 173.610 ;
        RECT 36.950 173.550 37.270 173.610 ;
        RECT 42.010 173.550 42.330 173.610 ;
        RECT 44.785 173.565 45.075 173.610 ;
        RECT 65.470 173.550 65.790 173.610 ;
        RECT 68.705 173.565 68.995 173.610 ;
        RECT 16.250 173.210 16.570 173.470 ;
        RECT 33.270 173.410 33.590 173.470 ;
        RECT 38.790 173.410 39.110 173.470 ;
        RECT 43.390 173.410 43.710 173.470 ;
        RECT 33.270 173.270 43.710 173.410 ;
        RECT 33.270 173.210 33.590 173.270 ;
        RECT 38.790 173.210 39.110 173.270 ;
        RECT 43.390 173.210 43.710 173.270 ;
        RECT 44.310 173.410 44.630 173.470 ;
        RECT 53.065 173.410 53.355 173.455 ;
        RECT 44.310 173.270 53.355 173.410 ;
        RECT 44.310 173.210 44.630 173.270 ;
        RECT 53.065 173.225 53.355 173.270 ;
        RECT 65.010 173.210 65.330 173.470 ;
        RECT 68.780 173.410 68.920 173.565 ;
        RECT 69.150 173.550 69.470 173.810 ;
        RECT 72.385 173.750 72.675 173.795 ;
        RECT 77.445 173.750 77.735 173.795 ;
        RECT 72.385 173.610 77.735 173.750 ;
        RECT 88.100 173.750 88.240 174.630 ;
        RECT 92.150 174.230 92.470 174.490 ;
        RECT 93.070 174.430 93.390 174.490 ;
        RECT 93.990 174.430 94.310 174.490 ;
        RECT 93.070 174.290 94.310 174.430 ;
        RECT 105.120 174.430 105.260 174.910 ;
        RECT 114.320 174.770 114.460 174.910 ;
        RECT 112.480 174.630 114.460 174.770 ;
        RECT 112.480 174.475 112.620 174.630 ;
        RECT 110.565 174.430 110.855 174.475 ;
        RECT 105.120 174.290 110.855 174.430 ;
        RECT 93.070 174.230 93.390 174.290 ;
        RECT 93.990 174.230 94.310 174.290 ;
        RECT 110.565 174.245 110.855 174.290 ;
        RECT 111.485 174.430 111.775 174.475 ;
        RECT 112.405 174.430 112.695 174.475 ;
        RECT 117.540 174.430 117.680 174.910 ;
        RECT 111.485 174.290 112.695 174.430 ;
        RECT 111.485 174.245 111.775 174.290 ;
        RECT 112.405 174.245 112.695 174.290 ;
        RECT 112.940 174.290 114.000 174.430 ;
        RECT 91.230 174.090 91.550 174.150 ;
        RECT 101.825 174.090 102.115 174.135 ;
        RECT 91.230 173.950 102.115 174.090 ;
        RECT 91.230 173.890 91.550 173.950 ;
        RECT 101.825 173.905 102.115 173.950 ;
        RECT 110.105 173.905 110.395 174.135 ;
        RECT 111.010 174.090 111.330 174.150 ;
        RECT 112.940 174.090 113.080 174.290 ;
        RECT 111.010 173.950 113.080 174.090 ;
        RECT 99.985 173.750 100.275 173.795 ;
        RECT 102.285 173.750 102.575 173.795 ;
        RECT 103.190 173.750 103.510 173.810 ;
        RECT 88.100 173.610 103.510 173.750 ;
        RECT 110.180 173.750 110.320 173.905 ;
        RECT 111.010 173.890 111.330 173.950 ;
        RECT 113.310 173.890 113.630 174.150 ;
        RECT 113.860 174.135 114.000 174.290 ;
        RECT 116.620 174.290 117.680 174.430 ;
        RECT 120.225 174.430 120.515 174.475 ;
        RECT 125.360 174.430 125.500 174.910 ;
        RECT 120.225 174.290 125.500 174.430 ;
        RECT 116.620 174.135 116.760 174.290 ;
        RECT 120.225 174.245 120.515 174.290 ;
        RECT 113.785 173.905 114.075 174.135 ;
        RECT 116.545 173.905 116.835 174.135 ;
        RECT 116.990 173.890 117.310 174.150 ;
        RECT 118.830 173.890 119.150 174.150 ;
        RECT 120.670 173.890 120.990 174.150 ;
        RECT 122.525 174.090 122.815 174.135 ;
        RECT 125.730 174.090 126.050 174.150 ;
        RECT 122.525 173.950 126.050 174.090 ;
        RECT 122.525 173.905 122.815 173.950 ;
        RECT 125.730 173.890 126.050 173.950 ;
        RECT 115.625 173.750 115.915 173.795 ;
        RECT 110.180 173.610 115.915 173.750 ;
        RECT 72.385 173.565 72.675 173.610 ;
        RECT 77.445 173.565 77.735 173.610 ;
        RECT 99.985 173.565 100.275 173.610 ;
        RECT 102.285 173.565 102.575 173.610 ;
        RECT 103.190 173.550 103.510 173.610 ;
        RECT 115.625 173.565 115.915 173.610 ;
        RECT 70.070 173.410 70.390 173.470 ;
        RECT 68.780 173.270 70.390 173.410 ;
        RECT 70.070 173.210 70.390 173.270 ;
        RECT 72.830 173.410 73.150 173.470 ;
        RECT 73.305 173.410 73.595 173.455 ;
        RECT 74.210 173.410 74.530 173.470 ;
        RECT 72.830 173.270 74.530 173.410 ;
        RECT 72.830 173.210 73.150 173.270 ;
        RECT 73.305 173.225 73.595 173.270 ;
        RECT 74.210 173.210 74.530 173.270 ;
        RECT 82.490 173.210 82.810 173.470 ;
        RECT 91.705 173.410 91.995 173.455 ;
        RECT 94.450 173.410 94.770 173.470 ;
        RECT 91.705 173.270 94.770 173.410 ;
        RECT 91.705 173.225 91.995 173.270 ;
        RECT 94.450 173.210 94.770 173.270 ;
        RECT 98.605 173.410 98.895 173.455 ;
        RECT 99.050 173.410 99.370 173.470 ;
        RECT 98.605 173.270 99.370 173.410 ;
        RECT 115.700 173.410 115.840 173.565 ;
        RECT 116.530 173.410 116.850 173.470 ;
        RECT 115.700 173.270 116.850 173.410 ;
        RECT 117.080 173.410 117.220 173.890 ;
        RECT 120.225 173.750 120.515 173.795 ;
        RECT 121.605 173.750 121.895 173.795 ;
        RECT 120.225 173.610 121.895 173.750 ;
        RECT 120.225 173.565 120.515 173.610 ;
        RECT 121.605 173.565 121.895 173.610 ;
        RECT 122.065 173.565 122.355 173.795 ;
        RECT 122.140 173.410 122.280 173.565 ;
        RECT 117.080 173.270 122.280 173.410 ;
        RECT 122.510 173.410 122.830 173.470 ;
        RECT 123.445 173.410 123.735 173.455 ;
        RECT 122.510 173.270 123.735 173.410 ;
        RECT 98.605 173.225 98.895 173.270 ;
        RECT 99.050 173.210 99.370 173.270 ;
        RECT 116.530 173.210 116.850 173.270 ;
        RECT 122.510 173.210 122.830 173.270 ;
        RECT 123.445 173.225 123.735 173.270 ;
        RECT 11.120 172.590 151.295 173.070 ;
        RECT 30.065 172.390 30.355 172.435 ;
        RECT 32.365 172.390 32.655 172.435 ;
        RECT 23.700 172.250 29.820 172.390 ;
        RECT 16.250 172.095 16.570 172.110 ;
        RECT 16.220 172.050 16.570 172.095 ;
        RECT 16.055 171.910 16.570 172.050 ;
        RECT 16.220 171.865 16.570 171.910 ;
        RECT 16.250 171.850 16.570 171.865 ;
        RECT 13.950 171.710 14.270 171.770 ;
        RECT 14.885 171.710 15.175 171.755 ;
        RECT 13.950 171.570 15.175 171.710 ;
        RECT 13.950 171.510 14.270 171.570 ;
        RECT 14.885 171.525 15.175 171.570 ;
        RECT 15.765 171.370 16.055 171.415 ;
        RECT 16.955 171.370 17.245 171.415 ;
        RECT 19.475 171.370 19.765 171.415 ;
        RECT 15.765 171.230 19.765 171.370 ;
        RECT 15.765 171.185 16.055 171.230 ;
        RECT 16.955 171.185 17.245 171.230 ;
        RECT 19.475 171.185 19.765 171.230 ;
        RECT 15.370 171.030 15.660 171.075 ;
        RECT 17.470 171.030 17.760 171.075 ;
        RECT 19.040 171.030 19.330 171.075 ;
        RECT 23.165 171.030 23.455 171.075 ;
        RECT 15.370 170.890 19.330 171.030 ;
        RECT 15.370 170.845 15.660 170.890 ;
        RECT 17.470 170.845 17.760 170.890 ;
        RECT 19.040 170.845 19.330 170.890 ;
        RECT 19.560 170.890 23.455 171.030 ;
        RECT 15.790 170.690 16.110 170.750 ;
        RECT 19.560 170.690 19.700 170.890 ;
        RECT 23.165 170.845 23.455 170.890 ;
        RECT 15.790 170.550 19.700 170.690 ;
        RECT 21.785 170.690 22.075 170.735 ;
        RECT 22.690 170.690 23.010 170.750 ;
        RECT 23.700 170.690 23.840 172.250 ;
        RECT 24.005 172.050 24.295 172.095 ;
        RECT 25.005 172.050 25.295 172.095 ;
        RECT 26.370 172.050 26.690 172.110 ;
        RECT 24.005 171.910 24.760 172.050 ;
        RECT 24.005 171.865 24.295 171.910 ;
        RECT 24.620 171.710 24.760 171.910 ;
        RECT 25.005 171.910 26.690 172.050 ;
        RECT 29.680 172.050 29.820 172.250 ;
        RECT 30.065 172.250 32.655 172.390 ;
        RECT 30.065 172.205 30.355 172.250 ;
        RECT 32.365 172.205 32.655 172.250 ;
        RECT 41.565 172.390 41.855 172.435 ;
        RECT 43.390 172.390 43.710 172.450 ;
        RECT 41.565 172.250 43.710 172.390 ;
        RECT 41.565 172.205 41.855 172.250 ;
        RECT 43.390 172.190 43.710 172.250 ;
        RECT 43.865 172.390 44.155 172.435 ;
        RECT 44.785 172.390 45.075 172.435 ;
        RECT 43.865 172.250 45.075 172.390 ;
        RECT 43.865 172.205 44.155 172.250 ;
        RECT 44.785 172.205 45.075 172.250 ;
        RECT 46.165 172.205 46.455 172.435 ;
        RECT 50.305 172.390 50.595 172.435 ;
        RECT 53.510 172.390 53.830 172.450 ;
        RECT 54.890 172.390 55.210 172.450 ;
        RECT 50.305 172.250 55.210 172.390 ;
        RECT 50.305 172.205 50.595 172.250 ;
        RECT 45.230 172.095 45.550 172.110 ;
        RECT 40.645 172.050 40.935 172.095 ;
        RECT 29.680 171.910 45.000 172.050 ;
        RECT 25.005 171.865 25.295 171.910 ;
        RECT 26.370 171.850 26.690 171.910 ;
        RECT 40.645 171.865 40.935 171.910 ;
        RECT 32.350 171.710 32.670 171.770 ;
        RECT 34.205 171.710 34.495 171.755 ;
        RECT 38.805 171.710 39.095 171.755 ;
        RECT 39.250 171.710 39.570 171.770 ;
        RECT 24.620 171.570 27.520 171.710 ;
        RECT 27.380 171.090 27.520 171.570 ;
        RECT 32.350 171.570 37.640 171.710 ;
        RECT 32.350 171.510 32.670 171.570 ;
        RECT 34.205 171.525 34.495 171.570 ;
        RECT 33.270 171.170 33.590 171.430 ;
        RECT 33.730 171.170 34.050 171.430 ;
        RECT 34.665 171.370 34.955 171.415 ;
        RECT 36.950 171.370 37.270 171.430 ;
        RECT 34.665 171.230 37.270 171.370 ;
        RECT 37.500 171.370 37.640 171.570 ;
        RECT 38.805 171.570 39.570 171.710 ;
        RECT 38.805 171.525 39.095 171.570 ;
        RECT 39.250 171.510 39.570 171.570 ;
        RECT 42.010 171.510 42.330 171.770 ;
        RECT 42.930 171.710 43.250 171.770 ;
        RECT 44.325 171.710 44.615 171.755 ;
        RECT 42.930 171.570 44.615 171.710 ;
        RECT 44.860 171.710 45.000 171.910 ;
        RECT 45.230 171.865 45.630 172.095 ;
        RECT 46.240 172.050 46.380 172.205 ;
        RECT 53.510 172.190 53.830 172.250 ;
        RECT 54.890 172.190 55.210 172.250 ;
        RECT 65.010 172.190 65.330 172.450 ;
        RECT 68.230 172.390 68.550 172.450 ;
        RECT 70.085 172.390 70.375 172.435 ;
        RECT 68.230 172.250 70.375 172.390 ;
        RECT 68.230 172.190 68.550 172.250 ;
        RECT 70.085 172.205 70.375 172.250 ;
        RECT 73.290 172.390 73.610 172.450 ;
        RECT 74.670 172.390 74.990 172.450 ;
        RECT 73.290 172.250 74.990 172.390 ;
        RECT 73.290 172.190 73.610 172.250 ;
        RECT 74.670 172.190 74.990 172.250 ;
        RECT 76.050 172.190 76.370 172.450 ;
        RECT 76.510 172.190 76.830 172.450 ;
        RECT 77.365 172.390 77.655 172.435 ;
        RECT 82.030 172.390 82.350 172.450 ;
        RECT 82.950 172.390 83.270 172.450 ;
        RECT 77.365 172.250 83.270 172.390 ;
        RECT 77.365 172.205 77.655 172.250 ;
        RECT 82.030 172.190 82.350 172.250 ;
        RECT 82.950 172.190 83.270 172.250 ;
        RECT 85.250 172.390 85.570 172.450 ;
        RECT 85.725 172.390 86.015 172.435 ;
        RECT 85.250 172.250 86.015 172.390 ;
        RECT 85.250 172.190 85.570 172.250 ;
        RECT 85.725 172.205 86.015 172.250 ;
        RECT 90.310 172.190 90.630 172.450 ;
        RECT 91.705 172.390 91.995 172.435 ;
        RECT 92.150 172.390 92.470 172.450 ;
        RECT 91.705 172.250 92.470 172.390 ;
        RECT 91.705 172.205 91.995 172.250 ;
        RECT 92.150 172.190 92.470 172.250 ;
        RECT 94.450 172.190 94.770 172.450 ;
        RECT 111.945 172.390 112.235 172.435 ;
        RECT 113.310 172.390 113.630 172.450 ;
        RECT 111.945 172.250 113.630 172.390 ;
        RECT 111.945 172.205 112.235 172.250 ;
        RECT 113.310 172.190 113.630 172.250 ;
        RECT 115.625 172.205 115.915 172.435 ;
        RECT 51.210 172.050 51.530 172.110 ;
        RECT 46.240 171.910 51.530 172.050 ;
        RECT 45.230 171.850 45.550 171.865 ;
        RECT 51.210 171.850 51.530 171.910 ;
        RECT 64.520 172.050 64.810 172.095 ;
        RECT 65.100 172.050 65.240 172.190 ;
        RECT 76.600 172.050 76.740 172.190 ;
        RECT 78.365 172.050 78.655 172.095 ;
        RECT 88.930 172.050 89.250 172.110 ;
        RECT 64.520 171.910 65.240 172.050 ;
        RECT 73.840 171.910 76.740 172.050 ;
        RECT 77.520 171.910 89.250 172.050 ;
        RECT 64.520 171.865 64.810 171.910 ;
        RECT 48.465 171.710 48.755 171.755 ;
        RECT 48.910 171.710 49.230 171.770 ;
        RECT 44.860 171.570 49.230 171.710 ;
        RECT 42.930 171.510 43.250 171.570 ;
        RECT 44.325 171.525 44.615 171.570 ;
        RECT 48.465 171.525 48.755 171.570 ;
        RECT 48.910 171.510 49.230 171.570 ;
        RECT 49.385 171.525 49.675 171.755 ;
        RECT 42.485 171.370 42.775 171.415 ;
        RECT 44.770 171.370 45.090 171.430 ;
        RECT 37.500 171.230 45.090 171.370 ;
        RECT 34.665 171.185 34.955 171.230 ;
        RECT 36.950 171.170 37.270 171.230 ;
        RECT 42.485 171.185 42.775 171.230 ;
        RECT 44.770 171.170 45.090 171.230 ;
        RECT 46.165 171.370 46.455 171.415 ;
        RECT 49.460 171.370 49.600 171.525 ;
        RECT 57.190 171.510 57.510 171.770 ;
        RECT 58.110 171.510 58.430 171.770 ;
        RECT 58.585 171.710 58.875 171.755 ;
        RECT 72.370 171.710 72.690 171.770 ;
        RECT 73.840 171.755 73.980 171.910 ;
        RECT 77.520 171.770 77.660 171.910 ;
        RECT 78.365 171.865 78.655 171.910 ;
        RECT 88.930 171.850 89.250 171.910 ;
        RECT 90.400 172.050 90.540 172.190 ;
        RECT 115.700 172.050 115.840 172.205 ;
        RECT 118.830 172.190 119.150 172.450 ;
        RECT 123.430 172.190 123.750 172.450 ;
        RECT 129.870 172.190 130.190 172.450 ;
        RECT 117.910 172.050 118.230 172.110 ;
        RECT 90.400 171.910 92.840 172.050 ;
        RECT 58.585 171.570 72.690 171.710 ;
        RECT 58.585 171.525 58.875 171.570 ;
        RECT 72.370 171.510 72.690 171.570 ;
        RECT 73.765 171.525 74.055 171.755 ;
        RECT 74.210 171.510 74.530 171.770 ;
        RECT 77.430 171.510 77.750 171.770 ;
        RECT 77.890 171.710 78.210 171.770 ;
        RECT 78.825 171.710 79.115 171.755 ;
        RECT 77.890 171.570 79.115 171.710 ;
        RECT 77.890 171.510 78.210 171.570 ;
        RECT 78.825 171.525 79.115 171.570 ;
        RECT 79.270 171.710 79.590 171.770 ;
        RECT 80.105 171.710 80.395 171.755 ;
        RECT 79.270 171.570 80.395 171.710 ;
        RECT 79.270 171.510 79.590 171.570 ;
        RECT 80.105 171.525 80.395 171.570 ;
        RECT 89.405 171.710 89.695 171.755 ;
        RECT 90.400 171.710 90.540 171.910 ;
        RECT 89.405 171.570 90.540 171.710 ;
        RECT 89.405 171.525 89.695 171.570 ;
        RECT 92.165 171.525 92.455 171.755 ;
        RECT 46.165 171.230 49.600 171.370 ;
        RECT 57.280 171.370 57.420 171.510 ;
        RECT 63.185 171.370 63.475 171.415 ;
        RECT 57.280 171.230 63.475 171.370 ;
        RECT 46.165 171.185 46.455 171.230 ;
        RECT 27.290 171.030 27.610 171.090 ;
        RECT 28.225 171.030 28.515 171.075 ;
        RECT 27.290 170.890 28.515 171.030 ;
        RECT 27.290 170.830 27.610 170.890 ;
        RECT 28.225 170.845 28.515 170.890 ;
        RECT 30.140 170.890 31.660 171.030 ;
        RECT 30.140 170.735 30.280 170.890 ;
        RECT 24.085 170.690 24.375 170.735 ;
        RECT 21.785 170.550 24.375 170.690 ;
        RECT 15.790 170.490 16.110 170.550 ;
        RECT 21.785 170.505 22.075 170.550 ;
        RECT 22.690 170.490 23.010 170.550 ;
        RECT 24.085 170.505 24.375 170.550 ;
        RECT 30.065 170.690 30.355 170.735 ;
        RECT 30.510 170.690 30.830 170.750 ;
        RECT 30.065 170.550 30.830 170.690 ;
        RECT 30.065 170.505 30.355 170.550 ;
        RECT 30.510 170.490 30.830 170.550 ;
        RECT 30.970 170.490 31.290 170.750 ;
        RECT 31.520 170.690 31.660 170.890 ;
        RECT 41.640 170.890 42.700 171.030 ;
        RECT 41.640 170.750 41.780 170.890 ;
        RECT 36.030 170.690 36.350 170.750 ;
        RECT 31.520 170.550 36.350 170.690 ;
        RECT 36.030 170.490 36.350 170.550 ;
        RECT 40.630 170.490 40.950 170.750 ;
        RECT 41.550 170.490 41.870 170.750 ;
        RECT 42.560 170.735 42.700 170.890 ;
        RECT 48.540 170.750 48.680 171.230 ;
        RECT 63.185 171.185 63.475 171.230 ;
        RECT 64.065 171.370 64.355 171.415 ;
        RECT 65.255 171.370 65.545 171.415 ;
        RECT 67.775 171.370 68.065 171.415 ;
        RECT 64.065 171.230 68.065 171.370 ;
        RECT 64.065 171.185 64.355 171.230 ;
        RECT 65.255 171.185 65.545 171.230 ;
        RECT 67.775 171.185 68.065 171.230 ;
        RECT 72.830 171.370 73.150 171.430 ;
        RECT 74.685 171.370 74.975 171.415 ;
        RECT 72.830 171.230 74.975 171.370 ;
        RECT 42.485 170.505 42.775 170.735 ;
        RECT 48.450 170.490 48.770 170.750 ;
        RECT 59.045 170.690 59.335 170.735 ;
        RECT 59.490 170.690 59.810 170.750 ;
        RECT 59.045 170.550 59.810 170.690 ;
        RECT 59.045 170.505 59.335 170.550 ;
        RECT 59.490 170.490 59.810 170.550 ;
        RECT 59.950 170.490 60.270 170.750 ;
        RECT 63.260 170.690 63.400 171.185 ;
        RECT 72.830 171.170 73.150 171.230 ;
        RECT 74.685 171.185 74.975 171.230 ;
        RECT 76.510 171.370 76.830 171.430 ;
        RECT 79.705 171.370 79.995 171.415 ;
        RECT 80.895 171.370 81.185 171.415 ;
        RECT 83.415 171.370 83.705 171.415 ;
        RECT 92.240 171.370 92.380 171.525 ;
        RECT 76.510 171.230 79.040 171.370 ;
        RECT 76.510 171.170 76.830 171.230 ;
        RECT 63.670 171.030 63.960 171.075 ;
        RECT 65.770 171.030 66.060 171.075 ;
        RECT 67.340 171.030 67.630 171.075 ;
        RECT 75.590 171.030 75.910 171.090 ;
        RECT 63.670 170.890 67.630 171.030 ;
        RECT 63.670 170.845 63.960 170.890 ;
        RECT 65.770 170.845 66.060 170.890 ;
        RECT 67.340 170.845 67.630 170.890 ;
        RECT 71.080 170.890 77.660 171.030 ;
        RECT 71.080 170.750 71.220 170.890 ;
        RECT 75.590 170.830 75.910 170.890 ;
        RECT 64.550 170.690 64.870 170.750 ;
        RECT 63.260 170.550 64.870 170.690 ;
        RECT 64.550 170.490 64.870 170.550 ;
        RECT 70.990 170.490 71.310 170.750 ;
        RECT 73.290 170.490 73.610 170.750 ;
        RECT 74.670 170.690 74.990 170.750 ;
        RECT 76.510 170.690 76.830 170.750 ;
        RECT 77.520 170.735 77.660 170.890 ;
        RECT 74.670 170.550 76.830 170.690 ;
        RECT 74.670 170.490 74.990 170.550 ;
        RECT 76.510 170.490 76.830 170.550 ;
        RECT 77.445 170.505 77.735 170.735 ;
        RECT 78.900 170.690 79.040 171.230 ;
        RECT 79.705 171.230 83.705 171.370 ;
        RECT 79.705 171.185 79.995 171.230 ;
        RECT 80.895 171.185 81.185 171.230 ;
        RECT 83.415 171.185 83.705 171.230 ;
        RECT 89.940 171.230 92.380 171.370 ;
        RECT 79.310 171.030 79.600 171.075 ;
        RECT 81.410 171.030 81.700 171.075 ;
        RECT 82.980 171.030 83.270 171.075 ;
        RECT 79.310 170.890 83.270 171.030 ;
        RECT 79.310 170.845 79.600 170.890 ;
        RECT 81.410 170.845 81.700 170.890 ;
        RECT 82.980 170.845 83.270 170.890 ;
        RECT 89.940 170.735 90.080 171.230 ;
        RECT 92.700 170.735 92.840 171.910 ;
        RECT 112.940 171.910 115.840 172.050 ;
        RECT 117.540 171.910 118.230 172.050 ;
        RECT 112.940 171.755 113.080 171.910 ;
        RECT 102.745 171.710 103.035 171.755 ;
        RECT 105.965 171.710 106.255 171.755 ;
        RECT 102.745 171.570 106.255 171.710 ;
        RECT 102.745 171.525 103.035 171.570 ;
        RECT 105.965 171.525 106.255 171.570 ;
        RECT 112.865 171.525 113.155 171.755 ;
        RECT 113.785 171.525 114.075 171.755 ;
        RECT 114.230 171.710 114.550 171.770 ;
        RECT 114.705 171.710 114.995 171.755 ;
        RECT 114.230 171.570 114.995 171.710 ;
        RECT 105.030 171.370 105.350 171.430 ;
        RECT 108.710 171.370 109.030 171.430 ;
        RECT 112.940 171.370 113.080 171.525 ;
        RECT 105.030 171.230 113.080 171.370 ;
        RECT 105.030 171.170 105.350 171.230 ;
        RECT 108.710 171.170 109.030 171.230 ;
        RECT 113.860 171.030 114.000 171.525 ;
        RECT 114.230 171.510 114.550 171.570 ;
        RECT 114.705 171.525 114.995 171.570 ;
        RECT 116.085 171.710 116.375 171.755 ;
        RECT 116.530 171.710 116.850 171.770 ;
        RECT 117.005 171.710 117.295 171.755 ;
        RECT 116.085 171.570 117.295 171.710 ;
        RECT 116.085 171.525 116.375 171.570 ;
        RECT 114.780 171.370 114.920 171.525 ;
        RECT 116.530 171.510 116.850 171.570 ;
        RECT 117.005 171.525 117.295 171.570 ;
        RECT 117.540 171.370 117.680 171.910 ;
        RECT 117.910 171.850 118.230 171.910 ;
        RECT 119.750 171.710 120.070 171.770 ;
        RECT 123.520 171.710 123.660 172.190 ;
        RECT 124.350 171.755 124.670 171.770 ;
        RECT 114.780 171.230 117.680 171.370 ;
        RECT 118.690 171.570 123.660 171.710 ;
        RECT 118.690 171.030 118.830 171.570 ;
        RECT 119.750 171.510 120.070 171.570 ;
        RECT 124.320 171.525 124.670 171.755 ;
        RECT 124.350 171.510 124.670 171.525 ;
        RECT 122.970 171.170 123.290 171.430 ;
        RECT 123.865 171.370 124.155 171.415 ;
        RECT 125.055 171.370 125.345 171.415 ;
        RECT 127.575 171.370 127.865 171.415 ;
        RECT 123.865 171.230 127.865 171.370 ;
        RECT 123.865 171.185 124.155 171.230 ;
        RECT 125.055 171.185 125.345 171.230 ;
        RECT 127.575 171.185 127.865 171.230 ;
        RECT 113.860 170.890 118.830 171.030 ;
        RECT 123.470 171.030 123.760 171.075 ;
        RECT 125.570 171.030 125.860 171.075 ;
        RECT 127.140 171.030 127.430 171.075 ;
        RECT 123.470 170.890 127.430 171.030 ;
        RECT 123.470 170.845 123.760 170.890 ;
        RECT 125.570 170.845 125.860 170.890 ;
        RECT 127.140 170.845 127.430 170.890 ;
        RECT 89.865 170.690 90.155 170.735 ;
        RECT 78.900 170.550 90.155 170.690 ;
        RECT 89.865 170.505 90.155 170.550 ;
        RECT 92.625 170.505 92.915 170.735 ;
        RECT 99.510 170.690 99.830 170.750 ;
        RECT 102.285 170.690 102.575 170.735 ;
        RECT 102.730 170.690 103.050 170.750 ;
        RECT 99.510 170.550 103.050 170.690 ;
        RECT 99.510 170.490 99.830 170.550 ;
        RECT 102.285 170.505 102.575 170.550 ;
        RECT 102.730 170.490 103.050 170.550 ;
        RECT 114.690 170.490 115.010 170.750 ;
        RECT 11.120 169.870 150.500 170.350 ;
        RECT 16.710 169.670 17.030 169.730 ;
        RECT 17.185 169.670 17.475 169.715 ;
        RECT 16.710 169.530 17.475 169.670 ;
        RECT 16.710 169.470 17.030 169.530 ;
        RECT 17.185 169.485 17.475 169.530 ;
        RECT 18.090 169.470 18.410 169.730 ;
        RECT 26.830 169.670 27.150 169.730 ;
        RECT 30.510 169.670 30.830 169.730 ;
        RECT 26.830 169.530 30.830 169.670 ;
        RECT 26.830 169.470 27.150 169.530 ;
        RECT 30.510 169.470 30.830 169.530 ;
        RECT 36.045 169.670 36.335 169.715 ;
        RECT 36.950 169.670 37.270 169.730 ;
        RECT 36.045 169.530 37.270 169.670 ;
        RECT 36.045 169.485 36.335 169.530 ;
        RECT 36.950 169.470 37.270 169.530 ;
        RECT 38.805 169.485 39.095 169.715 ;
        RECT 15.345 169.330 15.635 169.375 ;
        RECT 15.790 169.330 16.110 169.390 ;
        RECT 15.345 169.190 16.110 169.330 ;
        RECT 15.345 169.145 15.635 169.190 ;
        RECT 15.790 169.130 16.110 169.190 ;
        RECT 20.940 168.850 24.300 168.990 ;
        RECT 20.405 168.650 20.695 168.695 ;
        RECT 20.940 168.650 21.080 168.850 ;
        RECT 20.405 168.510 21.080 168.650 ;
        RECT 21.325 168.650 21.615 168.695 ;
        RECT 24.160 168.650 24.300 168.850 ;
        RECT 26.370 168.790 26.690 169.050 ;
        RECT 26.920 169.035 27.060 169.470 ;
        RECT 29.630 169.330 29.920 169.375 ;
        RECT 31.730 169.330 32.020 169.375 ;
        RECT 33.300 169.330 33.590 169.375 ;
        RECT 29.630 169.190 33.590 169.330 ;
        RECT 29.630 169.145 29.920 169.190 ;
        RECT 31.730 169.145 32.020 169.190 ;
        RECT 33.300 169.145 33.590 169.190 ;
        RECT 26.845 168.805 27.135 169.035 ;
        RECT 30.025 168.990 30.315 169.035 ;
        RECT 31.215 168.990 31.505 169.035 ;
        RECT 33.735 168.990 34.025 169.035 ;
        RECT 30.025 168.850 34.025 168.990 ;
        RECT 30.025 168.805 30.315 168.850 ;
        RECT 31.215 168.805 31.505 168.850 ;
        RECT 33.735 168.805 34.025 168.850 ;
        RECT 25.465 168.650 25.755 168.695 ;
        RECT 27.290 168.650 27.610 168.710 ;
        RECT 27.765 168.650 28.055 168.695 ;
        RECT 21.325 168.510 23.840 168.650 ;
        RECT 24.160 168.510 25.220 168.650 ;
        RECT 20.405 168.465 20.695 168.510 ;
        RECT 21.325 168.465 21.615 168.510 ;
        RECT 17.185 168.310 17.475 168.355 ;
        RECT 21.785 168.310 22.075 168.355 ;
        RECT 17.185 168.170 22.075 168.310 ;
        RECT 17.185 168.125 17.475 168.170 ;
        RECT 21.785 168.125 22.075 168.170 ;
        RECT 22.690 168.110 23.010 168.370 ;
        RECT 23.700 168.355 23.840 168.510 ;
        RECT 23.625 168.310 23.915 168.355 ;
        RECT 24.545 168.310 24.835 168.355 ;
        RECT 23.625 168.170 24.835 168.310 ;
        RECT 25.080 168.310 25.220 168.510 ;
        RECT 25.465 168.510 28.055 168.650 ;
        RECT 25.465 168.465 25.755 168.510 ;
        RECT 27.290 168.450 27.610 168.510 ;
        RECT 27.765 168.465 28.055 168.510 ;
        RECT 26.845 168.310 27.135 168.355 ;
        RECT 25.080 168.170 27.135 168.310 ;
        RECT 23.625 168.125 23.915 168.170 ;
        RECT 24.545 168.125 24.835 168.170 ;
        RECT 26.845 168.125 27.135 168.170 ;
        RECT 19.010 167.970 19.330 168.030 ;
        RECT 20.865 167.970 21.155 168.015 ;
        RECT 19.010 167.830 21.155 167.970 ;
        RECT 27.840 167.970 27.980 168.465 ;
        RECT 28.210 168.450 28.530 168.710 ;
        RECT 29.145 168.650 29.435 168.695 ;
        RECT 35.570 168.650 35.890 168.710 ;
        RECT 29.145 168.510 35.890 168.650 ;
        RECT 38.880 168.650 39.020 169.485 ;
        RECT 40.630 169.470 40.950 169.730 ;
        RECT 42.930 169.470 43.250 169.730 ;
        RECT 48.910 169.470 49.230 169.730 ;
        RECT 49.370 169.670 49.690 169.730 ;
        RECT 88.485 169.670 88.775 169.715 ;
        RECT 93.070 169.670 93.390 169.730 ;
        RECT 49.370 169.530 77.200 169.670 ;
        RECT 49.370 169.470 49.690 169.530 ;
        RECT 40.720 169.330 40.860 169.470 ;
        RECT 45.230 169.330 45.550 169.390 ;
        RECT 40.720 169.190 45.550 169.330 ;
        RECT 45.230 169.130 45.550 169.190 ;
        RECT 49.000 169.330 49.140 169.470 ;
        RECT 77.060 169.390 77.200 169.530 ;
        RECT 88.485 169.530 93.390 169.670 ;
        RECT 88.485 169.485 88.775 169.530 ;
        RECT 93.070 169.470 93.390 169.530 ;
        RECT 108.710 169.470 109.030 169.730 ;
        RECT 111.025 169.670 111.315 169.715 ;
        RECT 114.690 169.670 115.010 169.730 ;
        RECT 111.025 169.530 115.010 169.670 ;
        RECT 111.025 169.485 111.315 169.530 ;
        RECT 114.690 169.470 115.010 169.530 ;
        RECT 117.465 169.670 117.755 169.715 ;
        RECT 118.830 169.670 119.150 169.730 ;
        RECT 117.465 169.530 119.150 169.670 ;
        RECT 117.465 169.485 117.755 169.530 ;
        RECT 118.830 169.470 119.150 169.530 ;
        RECT 124.350 169.470 124.670 169.730 ;
        RECT 56.270 169.330 56.590 169.390 ;
        RECT 49.000 169.190 52.360 169.330 ;
        RECT 39.250 168.990 39.570 169.050 ;
        RECT 48.450 168.990 48.770 169.050 ;
        RECT 39.250 168.850 48.770 168.990 ;
        RECT 39.250 168.790 39.570 168.850 ;
        RECT 48.450 168.790 48.770 168.850 ;
        RECT 41.565 168.650 41.855 168.695 ;
        RECT 42.470 168.650 42.790 168.710 ;
        RECT 38.880 168.510 42.790 168.650 ;
        RECT 29.145 168.465 29.435 168.510 ;
        RECT 35.570 168.450 35.890 168.510 ;
        RECT 41.565 168.465 41.855 168.510 ;
        RECT 42.470 168.450 42.790 168.510 ;
        RECT 42.945 168.650 43.235 168.695 ;
        RECT 49.000 168.650 49.140 169.190 ;
        RECT 51.685 168.805 51.975 169.035 ;
        RECT 42.945 168.510 49.140 168.650 ;
        RECT 42.945 168.465 43.235 168.510 ;
        RECT 30.480 168.310 30.770 168.355 ;
        RECT 32.810 168.310 33.130 168.370 ;
        RECT 30.480 168.170 33.130 168.310 ;
        RECT 30.480 168.125 30.770 168.170 ;
        RECT 32.810 168.110 33.130 168.170 ;
        RECT 33.730 168.310 34.050 168.370 ;
        RECT 39.725 168.310 40.015 168.355 ;
        RECT 42.025 168.310 42.315 168.355 ;
        RECT 33.730 168.170 42.315 168.310 ;
        RECT 33.730 168.110 34.050 168.170 ;
        RECT 39.725 168.125 40.015 168.170 ;
        RECT 41.640 168.030 41.780 168.170 ;
        RECT 42.025 168.125 42.315 168.170 ;
        RECT 51.760 168.030 51.900 168.805 ;
        RECT 52.220 168.695 52.360 169.190 ;
        RECT 55.440 169.190 56.590 169.330 ;
        RECT 55.440 168.695 55.580 169.190 ;
        RECT 56.270 169.130 56.590 169.190 ;
        RECT 56.745 169.330 57.035 169.375 ;
        RECT 58.110 169.330 58.430 169.390 ;
        RECT 56.745 169.190 58.430 169.330 ;
        RECT 56.745 169.145 57.035 169.190 ;
        RECT 58.110 169.130 58.430 169.190 ;
        RECT 58.570 169.130 58.890 169.390 ;
        RECT 67.350 169.330 67.640 169.375 ;
        RECT 69.450 169.330 69.740 169.375 ;
        RECT 71.020 169.330 71.310 169.375 ;
        RECT 67.350 169.190 71.310 169.330 ;
        RECT 67.350 169.145 67.640 169.190 ;
        RECT 69.450 169.145 69.740 169.190 ;
        RECT 71.020 169.145 71.310 169.190 ;
        RECT 73.765 169.330 74.055 169.375 ;
        RECT 74.210 169.330 74.530 169.390 ;
        RECT 73.765 169.190 74.530 169.330 ;
        RECT 73.765 169.145 74.055 169.190 ;
        RECT 74.210 169.130 74.530 169.190 ;
        RECT 76.970 169.330 77.290 169.390 ;
        RECT 78.365 169.330 78.655 169.375 ;
        RECT 95.370 169.330 95.690 169.390 ;
        RECT 102.310 169.330 102.600 169.375 ;
        RECT 104.410 169.330 104.700 169.375 ;
        RECT 105.980 169.330 106.270 169.375 ;
        RECT 76.970 169.190 101.120 169.330 ;
        RECT 76.970 169.130 77.290 169.190 ;
        RECT 78.365 169.145 78.655 169.190 ;
        RECT 95.370 169.130 95.690 169.190 ;
        RECT 100.980 169.050 101.120 169.190 ;
        RECT 102.310 169.190 106.270 169.330 ;
        RECT 102.310 169.145 102.600 169.190 ;
        RECT 104.410 169.145 104.700 169.190 ;
        RECT 105.980 169.145 106.270 169.190 ;
        RECT 111.930 169.130 112.250 169.390 ;
        RECT 55.825 168.805 56.115 169.035 ;
        RECT 64.550 168.990 64.870 169.050 ;
        RECT 67.745 168.990 68.035 169.035 ;
        RECT 68.935 168.990 69.225 169.035 ;
        RECT 71.455 168.990 71.745 169.035 ;
        RECT 64.550 168.850 67.080 168.990 ;
        RECT 52.145 168.465 52.435 168.695 ;
        RECT 55.365 168.465 55.655 168.695 ;
        RECT 55.900 168.650 56.040 168.805 ;
        RECT 64.550 168.790 64.870 168.850 ;
        RECT 57.190 168.650 57.510 168.710 ;
        RECT 55.900 168.510 57.510 168.650 ;
        RECT 57.190 168.450 57.510 168.510 ;
        RECT 57.665 168.650 57.955 168.695 ;
        RECT 58.110 168.650 58.430 168.710 ;
        RECT 66.940 168.695 67.080 168.850 ;
        RECT 67.745 168.850 71.745 168.990 ;
        RECT 67.745 168.805 68.035 168.850 ;
        RECT 68.935 168.805 69.225 168.850 ;
        RECT 71.455 168.805 71.745 168.850 ;
        RECT 72.370 168.990 72.690 169.050 ;
        RECT 76.050 168.990 76.370 169.050 ;
        RECT 72.370 168.850 76.370 168.990 ;
        RECT 72.370 168.790 72.690 168.850 ;
        RECT 76.050 168.790 76.370 168.850 ;
        RECT 87.105 168.805 87.395 169.035 ;
        RECT 97.760 168.850 100.660 168.990 ;
        RECT 57.665 168.510 58.430 168.650 ;
        RECT 57.665 168.465 57.955 168.510 ;
        RECT 58.110 168.450 58.430 168.510 ;
        RECT 59.045 168.650 59.335 168.695 ;
        RECT 59.965 168.650 60.255 168.695 ;
        RECT 59.045 168.510 60.255 168.650 ;
        RECT 59.045 168.465 59.335 168.510 ;
        RECT 59.965 168.465 60.255 168.510 ;
        RECT 60.425 168.650 60.715 168.695 ;
        RECT 60.425 168.510 63.400 168.650 ;
        RECT 60.425 168.465 60.715 168.510 ;
        RECT 63.260 168.030 63.400 168.510 ;
        RECT 66.865 168.465 67.155 168.695 ;
        RECT 85.250 168.650 85.570 168.710 ;
        RECT 86.645 168.650 86.935 168.695 ;
        RECT 85.250 168.510 86.935 168.650 ;
        RECT 87.180 168.650 87.320 168.805 ;
        RECT 95.370 168.650 95.690 168.710 ;
        RECT 87.180 168.510 95.690 168.650 ;
        RECT 85.250 168.450 85.570 168.510 ;
        RECT 86.645 168.465 86.935 168.510 ;
        RECT 95.370 168.450 95.690 168.510 ;
        RECT 96.750 168.650 97.070 168.710 ;
        RECT 97.760 168.650 97.900 168.850 ;
        RECT 96.750 168.510 97.900 168.650 ;
        RECT 96.750 168.450 97.070 168.510 ;
        RECT 98.130 168.450 98.450 168.710 ;
        RECT 98.590 168.450 98.910 168.710 ;
        RECT 99.510 168.450 99.830 168.710 ;
        RECT 99.970 168.450 100.290 168.710 ;
        RECT 100.520 168.650 100.660 168.850 ;
        RECT 100.890 168.790 101.210 169.050 ;
        RECT 102.705 168.990 102.995 169.035 ;
        RECT 103.895 168.990 104.185 169.035 ;
        RECT 106.415 168.990 106.705 169.035 ;
        RECT 102.705 168.850 106.705 168.990 ;
        RECT 102.705 168.805 102.995 168.850 ;
        RECT 103.895 168.805 104.185 168.850 ;
        RECT 106.415 168.805 106.705 168.850 ;
        RECT 109.170 168.990 109.490 169.050 ;
        RECT 111.485 168.990 111.775 169.035 ;
        RECT 119.305 168.990 119.595 169.035 ;
        RECT 109.170 168.850 111.775 168.990 ;
        RECT 109.170 168.790 109.490 168.850 ;
        RECT 111.485 168.805 111.775 168.850 ;
        RECT 118.460 168.850 119.595 168.990 ;
        RECT 101.825 168.650 102.115 168.695 ;
        RECT 100.520 168.510 102.115 168.650 ;
        RECT 101.825 168.465 102.115 168.510 ;
        RECT 102.820 168.510 105.030 168.650 ;
        RECT 68.230 168.355 68.550 168.370 ;
        RECT 68.200 168.125 68.550 168.355 ;
        RECT 83.410 168.310 83.730 168.370 ;
        RECT 68.230 168.110 68.550 168.125 ;
        RECT 75.220 168.170 83.730 168.310 ;
        RECT 75.220 168.030 75.360 168.170 ;
        RECT 83.410 168.110 83.730 168.170 ;
        RECT 84.805 168.310 85.095 168.355 ;
        RECT 102.820 168.310 102.960 168.510 ;
        RECT 84.805 168.170 102.960 168.310 ;
        RECT 84.805 168.125 85.095 168.170 ;
        RECT 103.160 168.125 103.450 168.355 ;
        RECT 104.890 168.310 105.030 168.510 ;
        RECT 113.310 168.450 113.630 168.710 ;
        RECT 116.070 168.450 116.390 168.710 ;
        RECT 117.310 168.650 118.140 168.660 ;
        RECT 118.460 168.650 118.600 168.850 ;
        RECT 119.305 168.805 119.595 168.850 ;
        RECT 117.310 168.520 118.600 168.650 ;
        RECT 116.160 168.310 116.300 168.450 ;
        RECT 104.890 168.170 116.300 168.310 ;
        RECT 117.310 168.355 117.450 168.520 ;
        RECT 118.000 168.510 118.600 168.520 ;
        RECT 118.830 168.450 119.150 168.710 ;
        RECT 119.750 168.450 120.070 168.710 ;
        RECT 121.130 168.450 121.450 168.710 ;
        RECT 122.065 168.650 122.355 168.695 ;
        RECT 122.510 168.650 122.830 168.710 ;
        RECT 122.065 168.510 122.830 168.650 ;
        RECT 122.065 168.465 122.355 168.510 ;
        RECT 122.510 168.450 122.830 168.510 ;
        RECT 122.985 168.650 123.275 168.695 ;
        RECT 125.285 168.650 125.575 168.695 ;
        RECT 122.985 168.510 125.575 168.650 ;
        RECT 122.985 168.465 123.275 168.510 ;
        RECT 125.285 168.465 125.575 168.510 ;
        RECT 117.310 168.170 117.675 168.355 ;
        RECT 117.385 168.125 117.675 168.170 ;
        RECT 117.910 168.310 118.230 168.370 ;
        RECT 118.385 168.310 118.675 168.355 ;
        RECT 117.910 168.170 118.675 168.310 ;
        RECT 38.790 168.015 39.110 168.030 ;
        RECT 37.885 167.970 38.175 168.015 ;
        RECT 27.840 167.830 38.175 167.970 ;
        RECT 19.010 167.770 19.330 167.830 ;
        RECT 20.865 167.785 21.155 167.830 ;
        RECT 37.885 167.785 38.175 167.830 ;
        RECT 38.725 167.785 39.110 168.015 ;
        RECT 38.790 167.770 39.110 167.785 ;
        RECT 41.550 167.770 41.870 168.030 ;
        RECT 50.290 167.770 50.610 168.030 ;
        RECT 51.670 167.770 51.990 168.030 ;
        RECT 53.510 167.770 53.830 168.030 ;
        RECT 63.170 167.770 63.490 168.030 ;
        RECT 75.130 167.770 75.450 168.030 ;
        RECT 78.350 167.970 78.670 168.030 ;
        RECT 91.230 167.970 91.550 168.030 ;
        RECT 78.350 167.830 91.550 167.970 ;
        RECT 78.350 167.770 78.670 167.830 ;
        RECT 91.230 167.770 91.550 167.830 ;
        RECT 100.905 167.970 101.195 168.015 ;
        RECT 103.280 167.970 103.420 168.125 ;
        RECT 117.910 168.110 118.230 168.170 ;
        RECT 118.385 168.125 118.675 168.170 ;
        RECT 100.905 167.830 103.420 167.970 ;
        RECT 109.645 167.970 109.935 168.015 ;
        RECT 110.550 167.970 110.870 168.030 ;
        RECT 109.645 167.830 110.870 167.970 ;
        RECT 100.905 167.785 101.195 167.830 ;
        RECT 109.645 167.785 109.935 167.830 ;
        RECT 110.550 167.770 110.870 167.830 ;
        RECT 112.865 167.970 113.155 168.015 ;
        RECT 114.230 167.970 114.550 168.030 ;
        RECT 112.865 167.830 114.550 167.970 ;
        RECT 112.865 167.785 113.155 167.830 ;
        RECT 114.230 167.770 114.550 167.830 ;
        RECT 116.530 167.770 116.850 168.030 ;
        RECT 11.120 167.150 151.295 167.630 ;
        RECT 28.210 166.950 28.530 167.010 ;
        RECT 29.145 166.950 29.435 166.995 ;
        RECT 28.210 166.810 29.435 166.950 ;
        RECT 28.210 166.750 28.530 166.810 ;
        RECT 29.145 166.765 29.435 166.810 ;
        RECT 30.970 166.750 31.290 167.010 ;
        RECT 32.810 166.750 33.130 167.010 ;
        RECT 35.570 166.950 35.890 167.010 ;
        RECT 52.130 166.950 52.450 167.010 ;
        RECT 35.570 166.810 52.450 166.950 ;
        RECT 35.570 166.750 35.890 166.810 ;
        RECT 52.130 166.750 52.450 166.810 ;
        RECT 67.310 166.750 67.630 167.010 ;
        RECT 68.230 166.750 68.550 167.010 ;
        RECT 73.290 166.950 73.610 167.010 ;
        RECT 79.270 166.950 79.590 167.010 ;
        RECT 79.745 166.950 80.035 166.995 ;
        RECT 98.130 166.950 98.450 167.010 ;
        RECT 73.290 166.810 77.200 166.950 ;
        RECT 73.290 166.750 73.610 166.810 ;
        RECT 26.370 166.070 26.690 166.330 ;
        RECT 30.525 166.085 30.815 166.315 ;
        RECT 31.060 166.270 31.200 166.750 ;
        RECT 52.605 166.610 52.895 166.655 ;
        RECT 51.760 166.470 52.895 166.610 ;
        RECT 51.760 166.330 51.900 166.470 ;
        RECT 52.605 166.425 52.895 166.470 ;
        RECT 53.510 166.410 53.830 166.670 ;
        RECT 74.210 166.410 74.530 166.670 ;
        RECT 75.130 166.410 75.450 166.670 ;
        RECT 33.745 166.270 34.035 166.315 ;
        RECT 31.060 166.130 34.035 166.270 ;
        RECT 33.745 166.085 34.035 166.130 ;
        RECT 30.600 165.590 30.740 166.085 ;
        RECT 42.010 166.070 42.330 166.330 ;
        RECT 51.670 166.070 51.990 166.330 ;
        RECT 52.145 166.085 52.435 166.315 ;
        RECT 56.270 166.270 56.590 166.330 ;
        RECT 63.170 166.270 63.490 166.330 ;
        RECT 56.270 166.130 63.490 166.270 ;
        RECT 42.485 165.930 42.775 165.975 ;
        RECT 43.850 165.930 44.170 165.990 ;
        RECT 42.485 165.790 44.170 165.930 ;
        RECT 52.220 165.930 52.360 166.085 ;
        RECT 56.270 166.070 56.590 166.130 ;
        RECT 63.170 166.070 63.490 166.130 ;
        RECT 66.405 166.270 66.695 166.315 ;
        RECT 66.865 166.270 67.155 166.315 ;
        RECT 66.405 166.130 67.155 166.270 ;
        RECT 66.405 166.085 66.695 166.130 ;
        RECT 66.865 166.085 67.155 166.130 ;
        RECT 67.785 166.085 68.075 166.315 ;
        RECT 67.860 165.930 68.000 166.085 ;
        RECT 69.150 166.070 69.470 166.330 ;
        RECT 73.290 166.270 73.610 166.330 ;
        RECT 75.220 166.270 75.360 166.410 ;
        RECT 76.525 166.270 76.815 166.315 ;
        RECT 73.290 166.130 76.815 166.270 ;
        RECT 77.060 166.270 77.200 166.810 ;
        RECT 79.270 166.810 80.035 166.950 ;
        RECT 79.270 166.750 79.590 166.810 ;
        RECT 79.745 166.765 80.035 166.810 ;
        RECT 92.240 166.810 98.450 166.950 ;
        RECT 77.445 166.270 77.735 166.315 ;
        RECT 77.060 166.130 77.735 166.270 ;
        RECT 73.290 166.070 73.610 166.130 ;
        RECT 76.525 166.085 76.815 166.130 ;
        RECT 77.445 166.085 77.735 166.130 ;
        RECT 77.905 166.085 78.195 166.315 ;
        RECT 78.365 166.270 78.655 166.315 ;
        RECT 82.490 166.270 82.810 166.330 ;
        RECT 78.365 166.130 82.810 166.270 ;
        RECT 78.365 166.085 78.655 166.130 ;
        RECT 74.670 165.930 74.990 165.990 ;
        RECT 52.220 165.790 53.280 165.930 ;
        RECT 67.860 165.790 74.990 165.930 ;
        RECT 42.485 165.745 42.775 165.790 ;
        RECT 43.850 165.730 44.170 165.790 ;
        RECT 53.140 165.650 53.280 165.790 ;
        RECT 74.670 165.730 74.990 165.790 ;
        RECT 75.130 165.930 75.450 165.990 ;
        RECT 77.980 165.930 78.120 166.085 ;
        RECT 82.490 166.070 82.810 166.130 ;
        RECT 75.130 165.790 78.120 165.930 ;
        RECT 75.130 165.730 75.450 165.790 ;
        RECT 31.890 165.590 32.210 165.650 ;
        RECT 52.590 165.590 52.910 165.650 ;
        RECT 30.600 165.450 52.910 165.590 ;
        RECT 31.890 165.390 32.210 165.450 ;
        RECT 52.590 165.390 52.910 165.450 ;
        RECT 53.050 165.390 53.370 165.650 ;
        RECT 76.050 165.590 76.370 165.650 ;
        RECT 92.240 165.590 92.380 166.810 ;
        RECT 98.130 166.750 98.450 166.810 ;
        RECT 98.590 166.950 98.910 167.010 ;
        RECT 101.855 166.950 102.145 166.995 ;
        RECT 98.590 166.810 102.145 166.950 ;
        RECT 98.590 166.750 98.910 166.810 ;
        RECT 101.855 166.765 102.145 166.810 ;
        RECT 102.285 166.950 102.575 166.995 ;
        RECT 102.730 166.950 103.050 167.010 ;
        RECT 116.530 166.950 116.850 167.010 ;
        RECT 102.285 166.810 103.050 166.950 ;
        RECT 102.285 166.765 102.575 166.810 ;
        RECT 102.730 166.750 103.050 166.810 ;
        RECT 103.280 166.810 116.850 166.950 ;
        RECT 95.370 166.410 95.690 166.670 ;
        RECT 99.970 166.610 100.290 166.670 ;
        RECT 101.365 166.610 101.655 166.655 ;
        RECT 103.280 166.610 103.420 166.810 ;
        RECT 116.530 166.750 116.850 166.810 ;
        RECT 99.970 166.470 103.420 166.610 ;
        RECT 110.105 166.610 110.395 166.655 ;
        RECT 111.945 166.610 112.235 166.655 ;
        RECT 110.105 166.470 112.235 166.610 ;
        RECT 99.970 166.410 100.290 166.470 ;
        RECT 101.365 166.425 101.655 166.470 ;
        RECT 110.105 166.425 110.395 166.470 ;
        RECT 111.945 166.425 112.235 166.470 ;
        RECT 112.390 166.610 112.710 166.670 ;
        RECT 124.810 166.610 125.130 166.670 ;
        RECT 126.205 166.610 126.495 166.655 ;
        RECT 112.390 166.470 113.540 166.610 ;
        RECT 112.390 166.410 112.710 166.470 ;
        RECT 92.610 166.070 92.930 166.330 ;
        RECT 94.925 166.270 95.215 166.315 ;
        RECT 94.540 166.130 95.215 166.270 ;
        RECT 94.540 165.975 94.680 166.130 ;
        RECT 94.925 166.085 95.215 166.130 ;
        RECT 93.085 165.745 93.375 165.975 ;
        RECT 94.465 165.745 94.755 165.975 ;
        RECT 95.460 165.930 95.600 166.410 ;
        RECT 95.830 166.070 96.150 166.330 ;
        RECT 96.290 166.070 96.610 166.330 ;
        RECT 102.745 166.270 103.035 166.315 ;
        RECT 104.570 166.270 104.890 166.330 ;
        RECT 102.745 166.130 104.890 166.270 ;
        RECT 102.745 166.085 103.035 166.130 ;
        RECT 104.570 166.070 104.890 166.130 ;
        RECT 109.645 166.270 109.935 166.315 ;
        RECT 111.010 166.270 111.330 166.330 ;
        RECT 113.400 166.315 113.540 166.470 ;
        RECT 124.810 166.470 126.495 166.610 ;
        RECT 124.810 166.410 125.130 166.470 ;
        RECT 126.205 166.425 126.495 166.470 ;
        RECT 109.645 166.130 112.160 166.270 ;
        RECT 109.645 166.085 109.935 166.130 ;
        RECT 109.720 165.930 109.860 166.085 ;
        RECT 111.010 166.070 111.330 166.130 ;
        RECT 112.020 165.990 112.160 166.130 ;
        RECT 112.865 166.085 113.155 166.315 ;
        RECT 113.325 166.085 113.615 166.315 ;
        RECT 118.385 166.270 118.675 166.315 ;
        RECT 127.110 166.270 127.430 166.330 ;
        RECT 127.585 166.270 127.875 166.315 ;
        RECT 118.385 166.130 127.875 166.270 ;
        RECT 118.385 166.085 118.675 166.130 ;
        RECT 95.460 165.790 109.860 165.930 ;
        RECT 76.050 165.450 92.380 165.590 ;
        RECT 93.160 165.590 93.300 165.745 ;
        RECT 110.550 165.730 110.870 165.990 ;
        RECT 111.930 165.730 112.250 165.990 ;
        RECT 112.940 165.930 113.080 166.085 ;
        RECT 127.110 166.070 127.430 166.130 ;
        RECT 127.585 166.085 127.875 166.130 ;
        RECT 117.910 165.930 118.230 165.990 ;
        RECT 112.940 165.790 118.230 165.930 ;
        RECT 117.910 165.730 118.230 165.790 ;
        RECT 111.010 165.590 111.330 165.650 ;
        RECT 93.160 165.450 111.330 165.590 ;
        RECT 76.050 165.390 76.370 165.450 ;
        RECT 111.010 165.390 111.330 165.450 ;
        RECT 30.985 165.250 31.275 165.295 ;
        RECT 32.810 165.250 33.130 165.310 ;
        RECT 35.570 165.250 35.890 165.310 ;
        RECT 30.985 165.110 35.890 165.250 ;
        RECT 30.985 165.065 31.275 165.110 ;
        RECT 32.810 165.050 33.130 165.110 ;
        RECT 35.570 165.050 35.890 165.110 ;
        RECT 43.390 165.050 43.710 165.310 ;
        RECT 52.130 165.250 52.450 165.310 ;
        RECT 53.525 165.250 53.815 165.295 ;
        RECT 52.130 165.110 53.815 165.250 ;
        RECT 52.130 165.050 52.450 165.110 ;
        RECT 53.525 165.065 53.815 165.110 ;
        RECT 71.450 165.250 71.770 165.310 ;
        RECT 74.685 165.250 74.975 165.295 ;
        RECT 77.430 165.250 77.750 165.310 ;
        RECT 71.450 165.110 77.750 165.250 ;
        RECT 71.450 165.050 71.770 165.110 ;
        RECT 74.685 165.065 74.975 165.110 ;
        RECT 77.430 165.050 77.750 165.110 ;
        RECT 94.925 165.250 95.215 165.295 ;
        RECT 95.370 165.250 95.690 165.310 ;
        RECT 94.925 165.110 95.690 165.250 ;
        RECT 94.925 165.065 95.215 165.110 ;
        RECT 95.370 165.050 95.690 165.110 ;
        RECT 107.790 165.050 108.110 165.310 ;
        RECT 119.290 165.250 119.610 165.310 ;
        RECT 121.130 165.250 121.450 165.310 ;
        RECT 119.290 165.110 121.450 165.250 ;
        RECT 119.290 165.050 119.610 165.110 ;
        RECT 121.130 165.050 121.450 165.110 ;
        RECT 11.120 164.430 150.500 164.910 ;
        RECT 23.165 164.230 23.455 164.275 ;
        RECT 26.370 164.230 26.690 164.290 ;
        RECT 37.870 164.230 38.190 164.290 ;
        RECT 23.165 164.090 26.690 164.230 ;
        RECT 23.165 164.045 23.455 164.090 ;
        RECT 26.370 164.030 26.690 164.090 ;
        RECT 30.140 164.090 38.190 164.230 ;
        RECT 16.750 163.890 17.040 163.935 ;
        RECT 18.850 163.890 19.140 163.935 ;
        RECT 20.420 163.890 20.710 163.935 ;
        RECT 16.750 163.750 20.710 163.890 ;
        RECT 16.750 163.705 17.040 163.750 ;
        RECT 18.850 163.705 19.140 163.750 ;
        RECT 20.420 163.705 20.710 163.750 ;
        RECT 17.145 163.550 17.435 163.595 ;
        RECT 18.335 163.550 18.625 163.595 ;
        RECT 20.855 163.550 21.145 163.595 ;
        RECT 17.145 163.410 21.145 163.550 ;
        RECT 17.145 163.365 17.435 163.410 ;
        RECT 18.335 163.365 18.625 163.410 ;
        RECT 20.855 163.365 21.145 163.410 ;
        RECT 16.250 163.010 16.570 163.270 ;
        RECT 17.600 163.210 17.890 163.255 ;
        RECT 19.010 163.210 19.330 163.270 ;
        RECT 30.140 163.255 30.280 164.090 ;
        RECT 37.870 164.030 38.190 164.090 ;
        RECT 51.670 164.230 51.990 164.290 ;
        RECT 51.670 164.090 53.280 164.230 ;
        RECT 51.670 164.030 51.990 164.090 ;
        RECT 35.125 163.705 35.415 163.935 ;
        RECT 44.785 163.890 45.075 163.935 ;
        RECT 44.785 163.750 52.360 163.890 ;
        RECT 44.785 163.705 45.075 163.750 ;
        RECT 30.510 163.350 30.830 163.610 ;
        RECT 31.430 163.550 31.750 163.610 ;
        RECT 32.825 163.550 33.115 163.595 ;
        RECT 31.430 163.410 33.115 163.550 ;
        RECT 31.430 163.350 31.750 163.410 ;
        RECT 32.825 163.365 33.115 163.410 ;
        RECT 17.600 163.070 19.330 163.210 ;
        RECT 17.600 163.025 17.890 163.070 ;
        RECT 19.010 163.010 19.330 163.070 ;
        RECT 30.065 163.025 30.355 163.255 ;
        RECT 33.285 163.210 33.575 163.255 ;
        RECT 33.730 163.210 34.050 163.270 ;
        RECT 33.285 163.070 34.050 163.210 ;
        RECT 35.200 163.210 35.340 163.705 ;
        RECT 37.885 163.550 38.175 163.595 ;
        RECT 43.990 163.550 44.280 163.595 ;
        RECT 48.005 163.550 48.295 163.595 ;
        RECT 50.290 163.550 50.610 163.610 ;
        RECT 52.220 163.595 52.360 163.750 ;
        RECT 53.140 163.595 53.280 164.090 ;
        RECT 53.510 164.030 53.830 164.290 ;
        RECT 65.930 164.230 66.250 164.290 ;
        RECT 68.705 164.230 68.995 164.275 ;
        RECT 65.930 164.090 68.995 164.230 ;
        RECT 65.930 164.030 66.250 164.090 ;
        RECT 68.705 164.045 68.995 164.090 ;
        RECT 69.150 164.230 69.470 164.290 ;
        RECT 74.210 164.275 74.530 164.290 ;
        RECT 69.625 164.230 69.915 164.275 ;
        RECT 69.150 164.090 69.915 164.230 ;
        RECT 37.885 163.410 44.280 163.550 ;
        RECT 37.885 163.365 38.175 163.410 ;
        RECT 43.990 163.365 44.280 163.410 ;
        RECT 46.240 163.410 50.610 163.550 ;
        RECT 39.710 163.210 40.030 163.270 ;
        RECT 35.200 163.070 40.030 163.210 ;
        RECT 33.285 163.025 33.575 163.070 ;
        RECT 33.730 163.010 34.050 163.070 ;
        RECT 39.710 163.010 40.030 163.070 ;
        RECT 41.090 163.210 41.410 163.270 ;
        RECT 41.565 163.210 41.855 163.255 ;
        RECT 41.090 163.070 41.855 163.210 ;
        RECT 41.090 163.010 41.410 163.070 ;
        RECT 41.565 163.025 41.855 163.070 ;
        RECT 42.945 163.210 43.235 163.255 ;
        RECT 43.390 163.210 43.710 163.270 ;
        RECT 42.945 163.070 43.710 163.210 ;
        RECT 42.945 163.025 43.235 163.070 ;
        RECT 43.390 163.010 43.710 163.070 ;
        RECT 37.410 162.870 37.730 162.930 ;
        RECT 39.265 162.870 39.555 162.915 ;
        RECT 31.980 162.730 39.555 162.870 ;
        RECT 31.980 162.575 32.120 162.730 ;
        RECT 37.410 162.670 37.730 162.730 ;
        RECT 39.265 162.685 39.555 162.730 ;
        RECT 40.645 162.870 40.935 162.915 ;
        RECT 46.240 162.870 46.380 163.410 ;
        RECT 48.005 163.365 48.295 163.410 ;
        RECT 50.290 163.350 50.610 163.410 ;
        RECT 52.145 163.365 52.435 163.595 ;
        RECT 53.065 163.365 53.355 163.595 ;
        RECT 53.600 163.550 53.740 164.030 ;
        RECT 68.780 163.550 68.920 164.045 ;
        RECT 69.150 164.030 69.470 164.090 ;
        RECT 69.625 164.045 69.915 164.090 ;
        RECT 74.210 164.045 74.625 164.275 ;
        RECT 74.210 164.030 74.530 164.045 ;
        RECT 75.130 164.030 75.450 164.290 ;
        RECT 77.890 164.230 78.210 164.290 ;
        RECT 82.505 164.230 82.795 164.275 ;
        RECT 95.385 164.230 95.675 164.275 ;
        RECT 96.290 164.230 96.610 164.290 ;
        RECT 77.890 164.090 92.380 164.230 ;
        RECT 77.890 164.030 78.210 164.090 ;
        RECT 82.505 164.045 82.795 164.090 ;
        RECT 88.010 163.890 88.300 163.935 ;
        RECT 89.580 163.890 89.870 163.935 ;
        RECT 91.680 163.890 91.970 163.935 ;
        RECT 88.010 163.750 91.970 163.890 ;
        RECT 88.010 163.705 88.300 163.750 ;
        RECT 89.580 163.705 89.870 163.750 ;
        RECT 91.680 163.705 91.970 163.750 ;
        RECT 92.240 163.610 92.380 164.090 ;
        RECT 95.385 164.090 96.610 164.230 ;
        RECT 95.385 164.045 95.675 164.090 ;
        RECT 96.290 164.030 96.610 164.090 ;
        RECT 107.790 164.030 108.110 164.290 ;
        RECT 92.625 163.890 92.915 163.935 ;
        RECT 95.830 163.890 96.150 163.950 ;
        RECT 92.625 163.750 96.150 163.890 ;
        RECT 92.625 163.705 92.915 163.750 ;
        RECT 95.830 163.690 96.150 163.750 ;
        RECT 78.350 163.550 78.670 163.610 ;
        RECT 53.600 163.410 55.120 163.550 ;
        RECT 68.780 163.410 78.670 163.550 ;
        RECT 47.545 163.210 47.835 163.255 ;
        RECT 47.545 163.070 51.900 163.210 ;
        RECT 47.545 163.025 47.835 163.070 ;
        RECT 40.645 162.730 46.380 162.870 ;
        RECT 51.760 162.870 51.900 163.070 ;
        RECT 52.590 163.010 52.910 163.270 ;
        RECT 54.980 163.255 55.120 163.410 ;
        RECT 78.350 163.350 78.670 163.410 ;
        RECT 87.575 163.550 87.865 163.595 ;
        RECT 90.095 163.550 90.385 163.595 ;
        RECT 91.285 163.550 91.575 163.595 ;
        RECT 87.575 163.410 91.575 163.550 ;
        RECT 87.575 163.365 87.865 163.410 ;
        RECT 90.095 163.365 90.385 163.410 ;
        RECT 91.285 163.365 91.575 163.410 ;
        RECT 92.150 163.350 92.470 163.610 ;
        RECT 93.620 163.410 96.060 163.550 ;
        RECT 93.620 163.270 93.760 163.410 ;
        RECT 53.525 163.025 53.815 163.255 ;
        RECT 54.905 163.025 55.195 163.255 ;
        RECT 53.600 162.870 53.740 163.025 ;
        RECT 56.270 163.010 56.590 163.270 ;
        RECT 56.730 163.010 57.050 163.270 ;
        RECT 66.865 163.210 67.155 163.255 ;
        RECT 70.530 163.210 70.850 163.270 ;
        RECT 76.065 163.210 76.355 163.255 ;
        RECT 76.970 163.210 77.290 163.270 ;
        RECT 66.865 163.070 73.980 163.210 ;
        RECT 66.865 163.025 67.155 163.070 ;
        RECT 70.530 163.010 70.850 163.070 ;
        RECT 55.825 162.870 56.115 162.915 ;
        RECT 51.760 162.730 53.740 162.870 ;
        RECT 54.520 162.730 56.115 162.870 ;
        RECT 40.645 162.685 40.935 162.730 ;
        RECT 53.140 162.590 53.280 162.730 ;
        RECT 31.905 162.345 32.195 162.575 ;
        RECT 38.330 162.530 38.650 162.590 ;
        RECT 38.805 162.530 39.095 162.575 ;
        RECT 38.330 162.390 39.095 162.530 ;
        RECT 38.330 162.330 38.650 162.390 ;
        RECT 38.805 162.345 39.095 162.390 ;
        RECT 43.390 162.330 43.710 162.590 ;
        RECT 49.385 162.530 49.675 162.575 ;
        RECT 50.750 162.530 51.070 162.590 ;
        RECT 49.385 162.390 51.070 162.530 ;
        RECT 49.385 162.345 49.675 162.390 ;
        RECT 50.750 162.330 51.070 162.390 ;
        RECT 53.050 162.330 53.370 162.590 ;
        RECT 54.520 162.575 54.660 162.730 ;
        RECT 55.825 162.685 56.115 162.730 ;
        RECT 71.005 162.870 71.295 162.915 ;
        RECT 71.450 162.870 71.770 162.930 ;
        RECT 71.005 162.730 71.770 162.870 ;
        RECT 71.005 162.685 71.295 162.730 ;
        RECT 71.450 162.670 71.770 162.730 ;
        RECT 71.910 162.670 72.230 162.930 ;
        RECT 72.830 162.870 73.150 162.930 ;
        RECT 73.305 162.870 73.595 162.915 ;
        RECT 72.830 162.730 73.595 162.870 ;
        RECT 73.840 162.870 73.980 163.070 ;
        RECT 76.065 163.070 77.290 163.210 ;
        RECT 76.065 163.025 76.355 163.070 ;
        RECT 76.970 163.010 77.290 163.070 ;
        RECT 93.530 163.010 93.850 163.270 ;
        RECT 95.920 163.255 96.060 163.410 ;
        RECT 94.465 163.210 94.755 163.255 ;
        RECT 94.925 163.210 95.215 163.255 ;
        RECT 94.465 163.070 95.215 163.210 ;
        RECT 94.465 163.025 94.755 163.070 ;
        RECT 94.925 163.025 95.215 163.070 ;
        RECT 95.845 163.025 96.135 163.255 ;
        RECT 99.050 163.210 99.370 163.270 ;
        RECT 105.965 163.210 106.255 163.255 ;
        RECT 99.050 163.070 106.255 163.210 ;
        RECT 90.770 162.915 91.090 162.930 ;
        RECT 74.305 162.870 74.595 162.915 ;
        RECT 73.840 162.730 74.595 162.870 ;
        RECT 72.830 162.670 73.150 162.730 ;
        RECT 73.305 162.685 73.595 162.730 ;
        RECT 74.305 162.685 74.595 162.730 ;
        RECT 90.770 162.685 91.120 162.915 ;
        RECT 95.000 162.870 95.140 163.025 ;
        RECT 99.050 163.010 99.370 163.070 ;
        RECT 105.965 163.025 106.255 163.070 ;
        RECT 106.885 163.210 107.175 163.255 ;
        RECT 107.880 163.210 108.020 164.030 ;
        RECT 106.885 163.070 108.020 163.210 ;
        RECT 106.885 163.025 107.175 163.070 ;
        RECT 99.970 162.870 100.290 162.930 ;
        RECT 95.000 162.730 100.290 162.870 ;
        RECT 54.445 162.345 54.735 162.575 ;
        RECT 57.650 162.330 57.970 162.590 ;
        RECT 68.705 162.530 68.995 162.575 ;
        RECT 70.085 162.530 70.375 162.575 ;
        RECT 68.705 162.390 70.375 162.530 ;
        RECT 73.380 162.530 73.520 162.685 ;
        RECT 90.770 162.670 91.090 162.685 ;
        RECT 99.970 162.670 100.290 162.730 ;
        RECT 82.490 162.530 82.810 162.590 ;
        RECT 85.250 162.530 85.570 162.590 ;
        RECT 73.380 162.390 85.570 162.530 ;
        RECT 68.705 162.345 68.995 162.390 ;
        RECT 70.085 162.345 70.375 162.390 ;
        RECT 82.490 162.330 82.810 162.390 ;
        RECT 85.250 162.330 85.570 162.390 ;
        RECT 106.410 162.330 106.730 162.590 ;
        RECT 11.120 161.710 151.295 162.190 ;
        RECT 43.390 161.510 43.710 161.570 ;
        RECT 44.325 161.510 44.615 161.555 ;
        RECT 43.390 161.370 44.615 161.510 ;
        RECT 43.390 161.310 43.710 161.370 ;
        RECT 44.325 161.325 44.615 161.370 ;
        RECT 53.065 161.510 53.355 161.555 ;
        RECT 56.730 161.510 57.050 161.570 ;
        RECT 53.065 161.370 57.050 161.510 ;
        RECT 53.065 161.325 53.355 161.370 ;
        RECT 56.730 161.310 57.050 161.370 ;
        RECT 63.185 161.325 63.475 161.555 ;
        RECT 75.130 161.510 75.450 161.570 ;
        RECT 76.970 161.510 77.290 161.570 ;
        RECT 75.130 161.370 77.290 161.510 ;
        RECT 61.040 161.170 61.330 161.215 ;
        RECT 63.260 161.170 63.400 161.325 ;
        RECT 75.130 161.310 75.450 161.370 ;
        RECT 76.970 161.310 77.290 161.370 ;
        RECT 78.825 161.510 79.115 161.555 ;
        RECT 80.205 161.510 80.495 161.555 ;
        RECT 101.810 161.510 102.130 161.570 ;
        RECT 103.665 161.510 103.955 161.555 ;
        RECT 78.825 161.370 80.495 161.510 ;
        RECT 78.825 161.325 79.115 161.370 ;
        RECT 80.205 161.325 80.495 161.370 ;
        RECT 82.120 161.370 103.955 161.510 ;
        RECT 61.040 161.030 63.400 161.170 ;
        RECT 74.670 161.170 74.990 161.230 ;
        RECT 82.120 161.170 82.260 161.370 ;
        RECT 74.670 161.030 82.260 161.170 ;
        RECT 61.040 160.985 61.330 161.030 ;
        RECT 74.670 160.970 74.990 161.030 ;
        RECT 24.500 160.830 24.790 160.875 ;
        RECT 26.830 160.830 27.150 160.890 ;
        RECT 24.500 160.690 27.150 160.830 ;
        RECT 24.500 160.645 24.790 160.690 ;
        RECT 26.830 160.630 27.150 160.690 ;
        RECT 37.410 160.830 37.730 160.890 ;
        RECT 37.885 160.830 38.175 160.875 ;
        RECT 37.410 160.690 38.175 160.830 ;
        RECT 37.410 160.630 37.730 160.690 ;
        RECT 37.885 160.645 38.175 160.690 ;
        RECT 38.345 160.830 38.635 160.875 ;
        RECT 38.790 160.830 39.110 160.890 ;
        RECT 38.345 160.690 39.110 160.830 ;
        RECT 38.345 160.645 38.635 160.690 ;
        RECT 38.790 160.630 39.110 160.690 ;
        RECT 40.185 160.830 40.475 160.875 ;
        RECT 41.090 160.830 41.410 160.890 ;
        RECT 40.185 160.690 41.410 160.830 ;
        RECT 40.185 160.645 40.475 160.690 ;
        RECT 41.090 160.630 41.410 160.690 ;
        RECT 44.770 160.630 45.090 160.890 ;
        RECT 49.830 160.630 50.150 160.890 ;
        RECT 50.750 160.830 51.070 160.890 ;
        RECT 52.145 160.830 52.435 160.875 ;
        RECT 50.750 160.690 52.435 160.830 ;
        RECT 50.750 160.630 51.070 160.690 ;
        RECT 52.145 160.645 52.435 160.690 ;
        RECT 58.570 160.830 58.890 160.890 ;
        RECT 64.105 160.830 64.395 160.875 ;
        RECT 58.570 160.690 64.395 160.830 ;
        RECT 58.570 160.630 58.890 160.690 ;
        RECT 64.105 160.645 64.395 160.690 ;
        RECT 66.865 160.645 67.155 160.875 ;
        RECT 68.245 160.645 68.535 160.875 ;
        RECT 69.165 160.830 69.455 160.875 ;
        RECT 70.085 160.830 70.375 160.875 ;
        RECT 69.165 160.690 70.375 160.830 ;
        RECT 69.165 160.645 69.455 160.690 ;
        RECT 70.085 160.645 70.375 160.690 ;
        RECT 71.450 160.830 71.770 160.890 ;
        RECT 75.130 160.830 75.450 160.890 ;
        RECT 71.450 160.690 75.450 160.830 ;
        RECT 16.250 160.490 16.570 160.550 ;
        RECT 23.165 160.490 23.455 160.535 ;
        RECT 16.250 160.350 23.455 160.490 ;
        RECT 16.250 160.290 16.570 160.350 ;
        RECT 23.165 160.305 23.455 160.350 ;
        RECT 24.045 160.490 24.335 160.535 ;
        RECT 25.235 160.490 25.525 160.535 ;
        RECT 27.755 160.490 28.045 160.535 ;
        RECT 24.045 160.350 28.045 160.490 ;
        RECT 24.045 160.305 24.335 160.350 ;
        RECT 25.235 160.305 25.525 160.350 ;
        RECT 27.755 160.305 28.045 160.350 ;
        RECT 51.225 160.305 51.515 160.535 ;
        RECT 57.675 160.490 57.965 160.535 ;
        RECT 60.195 160.490 60.485 160.535 ;
        RECT 61.385 160.490 61.675 160.535 ;
        RECT 57.675 160.350 61.675 160.490 ;
        RECT 57.675 160.305 57.965 160.350 ;
        RECT 60.195 160.305 60.485 160.350 ;
        RECT 61.385 160.305 61.675 160.350 ;
        RECT 62.265 160.490 62.555 160.535 ;
        RECT 64.550 160.490 64.870 160.550 ;
        RECT 62.265 160.350 64.870 160.490 ;
        RECT 62.265 160.305 62.555 160.350 ;
        RECT 23.650 160.150 23.940 160.195 ;
        RECT 25.750 160.150 26.040 160.195 ;
        RECT 27.320 160.150 27.610 160.195 ;
        RECT 23.650 160.010 27.610 160.150 ;
        RECT 23.650 159.965 23.940 160.010 ;
        RECT 25.750 159.965 26.040 160.010 ;
        RECT 27.320 159.965 27.610 160.010 ;
        RECT 41.105 160.150 41.395 160.195 ;
        RECT 51.300 160.150 51.440 160.305 ;
        RECT 64.550 160.290 64.870 160.350 ;
        RECT 41.105 160.010 51.440 160.150 ;
        RECT 52.590 160.150 52.910 160.210 ;
        RECT 55.365 160.150 55.655 160.195 ;
        RECT 56.270 160.150 56.590 160.210 ;
        RECT 52.590 160.010 56.590 160.150 ;
        RECT 41.105 159.965 41.395 160.010 ;
        RECT 52.590 159.950 52.910 160.010 ;
        RECT 55.365 159.965 55.655 160.010 ;
        RECT 56.270 159.950 56.590 160.010 ;
        RECT 58.110 160.150 58.400 160.195 ;
        RECT 59.680 160.150 59.970 160.195 ;
        RECT 61.780 160.150 62.070 160.195 ;
        RECT 58.110 160.010 62.070 160.150 ;
        RECT 66.940 160.150 67.080 160.645 ;
        RECT 68.320 160.490 68.460 160.645 ;
        RECT 71.450 160.630 71.770 160.690 ;
        RECT 75.130 160.630 75.450 160.690 ;
        RECT 75.605 160.830 75.895 160.875 ;
        RECT 75.605 160.690 76.740 160.830 ;
        RECT 75.605 160.645 75.895 160.690 ;
        RECT 76.600 160.550 76.740 160.690 ;
        RECT 76.970 160.630 77.290 160.890 ;
        RECT 82.045 160.850 82.335 160.875 ;
        RECT 81.660 160.830 82.335 160.850 ;
        RECT 77.520 160.710 82.335 160.830 ;
        RECT 77.520 160.690 81.800 160.710 ;
        RECT 70.530 160.490 70.850 160.550 ;
        RECT 68.320 160.350 70.850 160.490 ;
        RECT 70.530 160.290 70.850 160.350 ;
        RECT 73.305 160.490 73.595 160.535 ;
        RECT 74.210 160.490 74.530 160.550 ;
        RECT 73.305 160.350 74.530 160.490 ;
        RECT 73.305 160.305 73.595 160.350 ;
        RECT 74.210 160.290 74.530 160.350 ;
        RECT 74.685 160.490 74.975 160.535 ;
        RECT 74.685 160.350 75.360 160.490 ;
        RECT 74.685 160.305 74.975 160.350 ;
        RECT 73.765 160.150 74.055 160.195 ;
        RECT 66.940 160.010 74.055 160.150 ;
        RECT 58.110 159.965 58.400 160.010 ;
        RECT 59.680 159.965 59.970 160.010 ;
        RECT 61.780 159.965 62.070 160.010 ;
        RECT 73.765 159.965 74.055 160.010 ;
        RECT 30.065 159.810 30.355 159.855 ;
        RECT 31.430 159.810 31.750 159.870 ;
        RECT 30.065 159.670 31.750 159.810 ;
        RECT 30.065 159.625 30.355 159.670 ;
        RECT 31.430 159.610 31.750 159.670 ;
        RECT 39.710 159.610 40.030 159.870 ;
        RECT 52.130 159.610 52.450 159.870 ;
        RECT 65.930 159.610 66.250 159.870 ;
        RECT 71.910 159.810 72.230 159.870 ;
        RECT 75.220 159.810 75.360 160.350 ;
        RECT 76.050 160.290 76.370 160.550 ;
        RECT 76.510 160.490 76.830 160.550 ;
        RECT 77.520 160.490 77.660 160.690 ;
        RECT 82.045 160.645 82.335 160.710 ;
        RECT 76.510 160.350 77.660 160.490 ;
        RECT 76.510 160.290 76.830 160.350 ;
        RECT 81.110 160.290 81.430 160.550 ;
        RECT 81.570 160.290 81.890 160.550 ;
        RECT 82.120 160.490 82.260 160.645 ;
        RECT 82.490 160.630 82.810 160.890 ;
        RECT 83.410 160.630 83.730 160.890 ;
        RECT 83.870 160.830 84.190 160.890 ;
        RECT 88.945 160.830 89.235 160.875 ;
        RECT 83.870 160.690 89.235 160.830 ;
        RECT 90.860 160.830 91.000 161.370 ;
        RECT 101.810 161.310 102.130 161.370 ;
        RECT 103.665 161.325 103.955 161.370 ;
        RECT 106.410 161.510 106.730 161.570 ;
        RECT 111.930 161.510 112.250 161.570 ;
        RECT 113.325 161.510 113.615 161.555 ;
        RECT 106.410 161.370 107.100 161.510 ;
        RECT 106.410 161.310 106.730 161.370 ;
        RECT 106.960 161.170 107.100 161.370 ;
        RECT 111.930 161.370 113.615 161.510 ;
        RECT 111.930 161.310 112.250 161.370 ;
        RECT 113.325 161.325 113.615 161.370 ;
        RECT 107.650 161.170 107.940 161.215 ;
        RECT 96.840 161.030 106.640 161.170 ;
        RECT 106.960 161.030 107.940 161.170 ;
        RECT 96.840 160.890 96.980 161.030 ;
        RECT 91.705 160.830 91.995 160.875 ;
        RECT 90.860 160.690 91.995 160.830 ;
        RECT 83.870 160.630 84.190 160.690 ;
        RECT 88.945 160.645 89.235 160.690 ;
        RECT 91.705 160.645 91.995 160.690 ;
        RECT 92.150 160.830 92.470 160.890 ;
        RECT 96.750 160.830 97.070 160.890 ;
        RECT 106.500 160.875 106.640 161.030 ;
        RECT 107.650 160.985 107.940 161.030 ;
        RECT 98.045 160.830 98.335 160.875 ;
        RECT 92.150 160.690 97.070 160.830 ;
        RECT 92.150 160.630 92.470 160.690 ;
        RECT 96.750 160.630 97.070 160.690 ;
        RECT 97.300 160.690 98.335 160.830 ;
        RECT 86.630 160.490 86.950 160.550 ;
        RECT 82.120 160.350 86.950 160.490 ;
        RECT 86.630 160.290 86.950 160.350 ;
        RECT 90.770 160.290 91.090 160.550 ;
        RECT 93.530 160.490 93.850 160.550 ;
        RECT 97.300 160.490 97.440 160.690 ;
        RECT 98.045 160.645 98.335 160.690 ;
        RECT 106.425 160.645 106.715 160.875 ;
        RECT 93.530 160.350 97.440 160.490 ;
        RECT 97.645 160.490 97.935 160.535 ;
        RECT 98.835 160.490 99.125 160.535 ;
        RECT 101.355 160.490 101.645 160.535 ;
        RECT 97.645 160.350 101.645 160.490 ;
        RECT 93.530 160.290 93.850 160.350 ;
        RECT 97.645 160.305 97.935 160.350 ;
        RECT 98.835 160.305 99.125 160.350 ;
        RECT 101.355 160.305 101.645 160.350 ;
        RECT 107.305 160.490 107.595 160.535 ;
        RECT 108.495 160.490 108.785 160.535 ;
        RECT 111.015 160.490 111.305 160.535 ;
        RECT 107.305 160.350 111.305 160.490 ;
        RECT 107.305 160.305 107.595 160.350 ;
        RECT 108.495 160.305 108.785 160.350 ;
        RECT 111.015 160.305 111.305 160.350 ;
        RECT 79.745 160.150 80.035 160.195 ;
        RECT 80.650 160.150 80.970 160.210 ;
        RECT 77.520 160.010 79.500 160.150 ;
        RECT 77.520 159.810 77.660 160.010 ;
        RECT 71.910 159.670 77.660 159.810 ;
        RECT 78.350 159.810 78.670 159.870 ;
        RECT 78.825 159.810 79.115 159.855 ;
        RECT 78.350 159.670 79.115 159.810 ;
        RECT 79.360 159.810 79.500 160.010 ;
        RECT 79.745 160.010 80.970 160.150 ;
        RECT 79.745 159.965 80.035 160.010 ;
        RECT 80.650 159.950 80.970 160.010 ;
        RECT 84.345 160.150 84.635 160.195 ;
        RECT 90.860 160.150 91.000 160.290 ;
        RECT 84.345 160.010 91.000 160.150 ;
        RECT 97.250 160.150 97.540 160.195 ;
        RECT 99.350 160.150 99.640 160.195 ;
        RECT 100.920 160.150 101.210 160.195 ;
        RECT 97.250 160.010 101.210 160.150 ;
        RECT 84.345 159.965 84.635 160.010 ;
        RECT 97.250 159.965 97.540 160.010 ;
        RECT 99.350 159.965 99.640 160.010 ;
        RECT 100.920 159.965 101.210 160.010 ;
        RECT 106.910 160.150 107.200 160.195 ;
        RECT 109.010 160.150 109.300 160.195 ;
        RECT 110.580 160.150 110.870 160.195 ;
        RECT 106.910 160.010 110.870 160.150 ;
        RECT 106.910 159.965 107.200 160.010 ;
        RECT 109.010 159.965 109.300 160.010 ;
        RECT 110.580 159.965 110.870 160.010 ;
        RECT 81.110 159.810 81.430 159.870 ;
        RECT 79.360 159.670 81.430 159.810 ;
        RECT 71.910 159.610 72.230 159.670 ;
        RECT 78.350 159.610 78.670 159.670 ;
        RECT 78.825 159.625 79.115 159.670 ;
        RECT 81.110 159.610 81.430 159.670 ;
        RECT 81.570 159.810 81.890 159.870 ;
        RECT 93.070 159.810 93.390 159.870 ;
        RECT 81.570 159.670 93.390 159.810 ;
        RECT 81.570 159.610 81.890 159.670 ;
        RECT 93.070 159.610 93.390 159.670 ;
        RECT 11.120 158.990 150.500 159.470 ;
        RECT 26.830 158.590 27.150 158.850 ;
        RECT 53.050 158.590 53.370 158.850 ;
        RECT 57.650 158.590 57.970 158.850 ;
        RECT 58.570 158.590 58.890 158.850 ;
        RECT 70.530 158.790 70.850 158.850 ;
        RECT 71.005 158.790 71.295 158.835 ;
        RECT 70.530 158.650 71.295 158.790 ;
        RECT 70.530 158.590 70.850 158.650 ;
        RECT 71.005 158.605 71.295 158.650 ;
        RECT 72.830 158.790 73.150 158.850 ;
        RECT 74.225 158.790 74.515 158.835 ;
        RECT 72.830 158.650 74.515 158.790 ;
        RECT 72.830 158.590 73.150 158.650 ;
        RECT 74.225 158.605 74.515 158.650 ;
        RECT 75.145 158.790 75.435 158.835 ;
        RECT 75.590 158.790 75.910 158.850 ;
        RECT 75.145 158.650 75.910 158.790 ;
        RECT 75.145 158.605 75.435 158.650 ;
        RECT 74.300 158.450 74.440 158.605 ;
        RECT 75.590 158.590 75.910 158.650 ;
        RECT 78.350 158.790 78.670 158.850 ;
        RECT 84.790 158.790 85.110 158.850 ;
        RECT 78.350 158.650 85.110 158.790 ;
        RECT 78.350 158.590 78.670 158.650 ;
        RECT 84.790 158.590 85.110 158.650 ;
        RECT 88.945 158.605 89.235 158.835 ;
        RECT 89.020 158.450 89.160 158.605 ;
        RECT 93.530 158.590 93.850 158.850 ;
        RECT 105.030 158.450 105.350 158.510 ;
        RECT 124.810 158.450 125.130 158.510 ;
        RECT 74.300 158.310 78.120 158.450 ;
        RECT 89.020 158.310 92.380 158.450 ;
        RECT 72.845 158.110 73.135 158.155 ;
        RECT 75.130 158.110 75.450 158.170 ;
        RECT 72.845 157.970 75.450 158.110 ;
        RECT 72.845 157.925 73.135 157.970 ;
        RECT 75.130 157.910 75.450 157.970 ;
        RECT 24.990 157.570 25.310 157.830 ;
        RECT 25.450 157.570 25.770 157.830 ;
        RECT 26.385 157.770 26.675 157.815 ;
        RECT 27.765 157.770 28.055 157.815 ;
        RECT 26.385 157.630 28.055 157.770 ;
        RECT 26.385 157.585 26.675 157.630 ;
        RECT 27.765 157.585 28.055 157.630 ;
        RECT 71.910 157.570 72.230 157.830 ;
        RECT 77.980 157.770 78.120 158.310 ;
        RECT 78.825 157.925 79.115 158.155 ;
        RECT 80.205 157.925 80.495 158.155 ;
        RECT 84.805 158.110 85.095 158.155 ;
        RECT 91.245 158.110 91.535 158.155 ;
        RECT 84.805 157.970 86.400 158.110 ;
        RECT 84.805 157.925 85.095 157.970 ;
        RECT 78.365 157.770 78.655 157.815 ;
        RECT 77.980 157.630 78.655 157.770 ;
        RECT 78.365 157.585 78.655 157.630 ;
        RECT 42.010 157.430 42.330 157.490 ;
        RECT 50.305 157.430 50.595 157.475 ;
        RECT 42.010 157.290 50.595 157.430 ;
        RECT 42.010 157.230 42.330 157.290 ;
        RECT 50.305 157.245 50.595 157.290 ;
        RECT 56.745 157.430 57.035 157.475 ;
        RECT 60.410 157.430 60.730 157.490 ;
        RECT 56.745 157.290 60.730 157.430 ;
        RECT 56.745 157.245 57.035 157.290 ;
        RECT 60.410 157.230 60.730 157.290 ;
        RECT 73.305 157.430 73.595 157.475 ;
        RECT 73.305 157.290 78.580 157.430 ;
        RECT 73.305 157.245 73.595 157.290 ;
        RECT 78.440 157.150 78.580 157.290 ;
        RECT 41.090 157.090 41.410 157.150 ;
        RECT 51.210 157.090 51.530 157.150 ;
        RECT 41.090 156.950 51.530 157.090 ;
        RECT 41.090 156.890 41.410 156.950 ;
        RECT 51.210 156.890 51.530 156.950 ;
        RECT 51.670 156.890 51.990 157.150 ;
        RECT 52.145 157.090 52.435 157.135 ;
        RECT 53.050 157.090 53.370 157.150 ;
        RECT 52.145 156.950 53.370 157.090 ;
        RECT 52.145 156.905 52.435 156.950 ;
        RECT 53.050 156.890 53.370 156.950 ;
        RECT 57.190 157.090 57.510 157.150 ;
        RECT 57.745 157.090 58.035 157.135 ;
        RECT 57.190 156.950 58.035 157.090 ;
        RECT 57.190 156.890 57.510 156.950 ;
        RECT 57.745 156.905 58.035 156.950 ;
        RECT 70.990 157.090 71.310 157.150 ;
        RECT 74.210 157.135 74.530 157.150 ;
        RECT 74.210 157.090 74.645 157.135 ;
        RECT 76.510 157.090 76.830 157.150 ;
        RECT 70.990 156.950 76.830 157.090 ;
        RECT 70.990 156.890 71.310 156.950 ;
        RECT 74.210 156.905 74.645 156.950 ;
        RECT 74.210 156.890 74.530 156.905 ;
        RECT 76.510 156.890 76.830 156.950 ;
        RECT 78.350 156.890 78.670 157.150 ;
        RECT 78.900 157.090 79.040 157.925 ;
        RECT 80.280 157.430 80.420 157.925 ;
        RECT 84.330 157.570 84.650 157.830 ;
        RECT 85.265 157.585 85.555 157.815 ;
        RECT 85.340 157.430 85.480 157.585 ;
        RECT 85.710 157.570 86.030 157.830 ;
        RECT 86.260 157.815 86.400 157.970 ;
        RECT 87.180 157.970 91.535 158.110 ;
        RECT 87.180 157.815 87.320 157.970 ;
        RECT 91.245 157.925 91.535 157.970 ;
        RECT 91.690 157.910 92.010 158.170 ;
        RECT 88.010 157.815 88.330 157.830 ;
        RECT 86.190 157.585 86.480 157.815 ;
        RECT 87.105 157.585 87.395 157.815 ;
        RECT 88.010 157.770 88.340 157.815 ;
        RECT 88.010 157.630 88.525 157.770 ;
        RECT 88.010 157.585 88.340 157.630 ;
        RECT 88.010 157.570 88.330 157.585 ;
        RECT 80.280 157.290 85.480 157.430 ;
        RECT 83.410 157.090 83.730 157.150 ;
        RECT 78.900 156.950 83.730 157.090 ;
        RECT 85.340 157.090 85.480 157.290 ;
        RECT 87.550 157.230 87.870 157.490 ;
        RECT 89.390 157.230 89.710 157.490 ;
        RECT 90.310 157.430 90.630 157.490 ;
        RECT 89.940 157.290 90.630 157.430 ;
        RECT 91.780 157.430 91.920 157.910 ;
        RECT 92.240 157.770 92.380 158.310 ;
        RECT 95.920 158.310 125.130 158.450 ;
        RECT 92.610 158.110 92.930 158.170 ;
        RECT 95.920 158.110 96.060 158.310 ;
        RECT 105.030 158.250 105.350 158.310 ;
        RECT 124.810 158.250 125.130 158.310 ;
        RECT 97.225 158.110 97.515 158.155 ;
        RECT 99.050 158.110 99.370 158.170 ;
        RECT 92.610 157.970 96.060 158.110 ;
        RECT 92.610 157.910 92.930 157.970 ;
        RECT 94.925 157.770 95.215 157.815 ;
        RECT 92.240 157.630 95.215 157.770 ;
        RECT 94.925 157.585 95.215 157.630 ;
        RECT 95.370 157.570 95.690 157.830 ;
        RECT 95.920 157.815 96.060 157.970 ;
        RECT 96.840 157.970 97.515 158.110 ;
        RECT 96.840 157.815 96.980 157.970 ;
        RECT 97.225 157.925 97.515 157.970 ;
        RECT 97.760 157.970 99.370 158.110 ;
        RECT 95.845 157.585 96.135 157.815 ;
        RECT 96.765 157.585 97.055 157.815 ;
        RECT 97.760 157.430 97.900 157.970 ;
        RECT 99.050 157.910 99.370 157.970 ;
        RECT 99.525 158.110 99.815 158.155 ;
        RECT 101.810 158.110 102.130 158.170 ;
        RECT 99.525 157.970 102.130 158.110 ;
        RECT 99.525 157.925 99.815 157.970 ;
        RECT 101.810 157.910 102.130 157.970 ;
        RECT 103.190 157.910 103.510 158.170 ;
        RECT 98.130 157.570 98.450 157.830 ;
        RECT 98.605 157.585 98.895 157.815 ;
        RECT 101.350 157.770 101.670 157.830 ;
        RECT 103.665 157.770 103.955 157.815 ;
        RECT 101.350 157.630 103.955 157.770 ;
        RECT 91.780 157.290 97.900 157.430 ;
        RECT 89.940 157.090 90.080 157.290 ;
        RECT 90.310 157.230 90.630 157.290 ;
        RECT 85.340 156.950 90.080 157.090 ;
        RECT 95.830 157.090 96.150 157.150 ;
        RECT 98.680 157.090 98.820 157.585 ;
        RECT 101.350 157.570 101.670 157.630 ;
        RECT 103.665 157.585 103.955 157.630 ;
        RECT 110.090 157.570 110.410 157.830 ;
        RECT 95.830 156.950 98.820 157.090 ;
        RECT 101.350 157.090 101.670 157.150 ;
        RECT 101.825 157.090 102.115 157.135 ;
        RECT 101.350 156.950 102.115 157.090 ;
        RECT 83.410 156.890 83.730 156.950 ;
        RECT 95.830 156.890 96.150 156.950 ;
        RECT 101.350 156.890 101.670 156.950 ;
        RECT 101.825 156.905 102.115 156.950 ;
        RECT 109.170 157.090 109.490 157.150 ;
        RECT 110.565 157.090 110.855 157.135 ;
        RECT 109.170 156.950 110.855 157.090 ;
        RECT 109.170 156.890 109.490 156.950 ;
        RECT 110.565 156.905 110.855 156.950 ;
        RECT 11.120 156.270 151.295 156.750 ;
        RECT 25.450 156.070 25.770 156.130 ;
        RECT 29.145 156.070 29.435 156.115 ;
        RECT 25.450 155.930 29.435 156.070 ;
        RECT 25.450 155.870 25.770 155.930 ;
        RECT 29.145 155.885 29.435 155.930 ;
        RECT 32.350 156.070 32.670 156.130 ;
        RECT 42.470 156.070 42.790 156.130 ;
        RECT 48.005 156.070 48.295 156.115 ;
        RECT 49.830 156.070 50.150 156.130 ;
        RECT 32.350 155.930 34.880 156.070 ;
        RECT 32.350 155.870 32.670 155.930 ;
        RECT 30.525 155.730 30.815 155.775 ;
        RECT 31.430 155.730 31.750 155.790 ;
        RECT 30.525 155.590 34.420 155.730 ;
        RECT 30.525 155.545 30.815 155.590 ;
        RECT 31.430 155.530 31.750 155.590 ;
        RECT 34.280 155.450 34.420 155.590 ;
        RECT 19.010 155.190 19.330 155.450 ;
        RECT 30.065 155.205 30.355 155.435 ;
        RECT 30.140 155.050 30.280 155.205 ;
        RECT 30.970 155.190 31.290 155.450 ;
        RECT 31.890 155.190 32.210 155.450 ;
        RECT 34.190 155.190 34.510 155.450 ;
        RECT 34.740 155.435 34.880 155.930 ;
        RECT 40.260 155.930 47.300 156.070 ;
        RECT 39.710 155.530 40.030 155.790 ;
        RECT 40.260 155.775 40.400 155.930 ;
        RECT 42.470 155.870 42.790 155.930 ;
        RECT 40.185 155.545 40.475 155.775 ;
        RECT 44.770 155.730 45.090 155.790 ;
        RECT 41.180 155.590 46.380 155.730 ;
        RECT 40.745 155.500 41.035 155.545 ;
        RECT 41.180 155.500 41.320 155.590 ;
        RECT 44.770 155.530 45.090 155.590 ;
        RECT 34.665 155.205 34.955 155.435 ;
        RECT 38.805 155.390 39.095 155.435 ;
        RECT 39.250 155.390 39.570 155.450 ;
        RECT 36.120 155.250 39.570 155.390 ;
        RECT 40.745 155.360 41.320 155.500 ;
        RECT 40.745 155.315 41.035 155.360 ;
        RECT 30.140 154.910 32.120 155.050 ;
        RECT 31.980 154.430 32.120 154.910 ;
        RECT 34.740 154.710 34.880 155.205 ;
        RECT 35.110 154.850 35.430 155.110 ;
        RECT 36.120 154.710 36.260 155.250 ;
        RECT 38.805 155.205 39.095 155.250 ;
        RECT 39.250 155.190 39.570 155.250 ;
        RECT 41.565 155.205 41.855 155.435 ;
        RECT 38.330 155.050 38.650 155.110 ;
        RECT 36.580 154.910 38.650 155.050 ;
        RECT 36.580 154.755 36.720 154.910 ;
        RECT 38.330 154.850 38.650 154.910 ;
        RECT 41.090 155.050 41.410 155.110 ;
        RECT 41.640 155.050 41.780 155.205 ;
        RECT 42.010 155.190 42.330 155.450 ;
        RECT 42.930 155.190 43.250 155.450 ;
        RECT 43.865 155.390 44.155 155.435 ;
        RECT 44.325 155.390 44.615 155.435 ;
        RECT 43.865 155.250 44.615 155.390 ;
        RECT 43.865 155.205 44.155 155.250 ;
        RECT 44.325 155.205 44.615 155.250 ;
        RECT 45.230 155.190 45.550 155.450 ;
        RECT 46.240 155.095 46.380 155.590 ;
        RECT 47.160 155.435 47.300 155.930 ;
        RECT 48.005 155.930 50.150 156.070 ;
        RECT 48.005 155.885 48.295 155.930 ;
        RECT 49.830 155.870 50.150 155.930 ;
        RECT 50.380 155.930 53.740 156.070 ;
        RECT 48.450 155.730 48.770 155.790 ;
        RECT 50.380 155.730 50.520 155.930 ;
        RECT 48.450 155.590 50.520 155.730 ;
        RECT 48.450 155.530 48.770 155.590 ;
        RECT 53.080 155.435 53.340 155.480 ;
        RECT 53.600 155.435 53.740 155.930 ;
        RECT 57.190 155.870 57.510 156.130 ;
        RECT 59.950 155.870 60.270 156.130 ;
        RECT 65.930 155.870 66.250 156.130 ;
        RECT 70.990 155.870 71.310 156.130 ;
        RECT 73.750 156.070 74.070 156.130 ;
        RECT 85.265 156.070 85.555 156.115 ;
        RECT 85.710 156.070 86.030 156.130 ;
        RECT 73.750 155.930 84.100 156.070 ;
        RECT 73.750 155.870 74.070 155.930 ;
        RECT 56.730 155.530 57.050 155.790 ;
        RECT 47.085 155.205 47.375 155.435 ;
        RECT 50.305 155.390 50.595 155.435 ;
        RECT 53.065 155.390 53.355 155.435 ;
        RECT 50.305 155.250 53.355 155.390 ;
        RECT 50.305 155.205 50.595 155.250 ;
        RECT 53.065 155.205 53.355 155.250 ;
        RECT 53.525 155.205 53.815 155.435 ;
        RECT 53.080 155.160 53.340 155.205 ;
        RECT 56.270 155.190 56.590 155.450 ;
        RECT 56.820 155.390 56.960 155.530 ;
        RECT 57.205 155.390 57.495 155.435 ;
        RECT 56.820 155.250 57.495 155.390 ;
        RECT 57.205 155.205 57.495 155.250 ;
        RECT 59.045 155.390 59.335 155.435 ;
        RECT 60.040 155.390 60.180 155.870 ;
        RECT 65.440 155.730 65.730 155.775 ;
        RECT 66.020 155.730 66.160 155.870 ;
        RECT 73.840 155.730 73.980 155.870 ;
        RECT 65.440 155.590 66.160 155.730 ;
        RECT 72.460 155.590 73.980 155.730 ;
        RECT 65.440 155.545 65.730 155.590 ;
        RECT 59.045 155.250 60.180 155.390 ;
        RECT 64.105 155.390 64.395 155.435 ;
        RECT 64.550 155.390 64.870 155.450 ;
        RECT 72.460 155.435 72.600 155.590 ;
        RECT 82.950 155.530 83.270 155.790 ;
        RECT 83.410 155.530 83.730 155.790 ;
        RECT 64.105 155.250 64.870 155.390 ;
        RECT 59.045 155.205 59.335 155.250 ;
        RECT 64.105 155.205 64.395 155.250 ;
        RECT 64.550 155.190 64.870 155.250 ;
        RECT 72.385 155.205 72.675 155.435 ;
        RECT 83.040 155.390 83.180 155.530 ;
        RECT 73.840 155.250 83.180 155.390 ;
        RECT 83.960 155.380 84.100 155.930 ;
        RECT 85.265 155.930 86.030 156.070 ;
        RECT 85.265 155.885 85.555 155.930 ;
        RECT 85.710 155.870 86.030 155.930 ;
        RECT 95.830 155.870 96.150 156.130 ;
        RECT 96.305 156.070 96.595 156.115 ;
        RECT 98.130 156.070 98.450 156.130 ;
        RECT 96.305 155.930 98.450 156.070 ;
        RECT 96.305 155.885 96.595 155.930 ;
        RECT 98.130 155.870 98.450 155.930 ;
        RECT 101.810 156.070 102.130 156.130 ;
        RECT 101.810 155.930 102.500 156.070 ;
        RECT 101.810 155.870 102.130 155.930 ;
        RECT 84.330 155.775 84.650 155.790 ;
        RECT 84.330 155.730 84.795 155.775 ;
        RECT 86.170 155.730 86.490 155.790 ;
        RECT 89.390 155.730 89.710 155.790 ;
        RECT 84.330 155.590 89.710 155.730 ;
        RECT 84.330 155.545 84.795 155.590 ;
        RECT 84.330 155.530 84.650 155.545 ;
        RECT 86.170 155.530 86.490 155.590 ;
        RECT 89.390 155.530 89.710 155.590 ;
        RECT 91.230 155.730 91.550 155.790 ;
        RECT 102.360 155.775 102.500 155.930 ;
        RECT 97.225 155.730 97.515 155.775 ;
        RECT 91.230 155.590 97.515 155.730 ;
        RECT 91.230 155.530 91.550 155.590 ;
        RECT 97.225 155.545 97.515 155.590 ;
        RECT 101.285 155.730 101.575 155.775 ;
        RECT 101.285 155.590 102.040 155.730 ;
        RECT 101.285 155.545 101.575 155.590 ;
        RECT 101.900 155.450 102.040 155.590 ;
        RECT 102.285 155.545 102.575 155.775 ;
        RECT 87.105 155.390 87.395 155.435 ;
        RECT 87.550 155.390 87.870 155.450 ;
        RECT 84.420 155.380 87.870 155.390 ;
        RECT 83.960 155.250 87.870 155.380 ;
        RECT 73.840 155.095 73.980 155.250 ;
        RECT 83.960 155.240 84.560 155.250 ;
        RECT 87.105 155.205 87.395 155.250 ;
        RECT 87.550 155.190 87.870 155.250 ;
        RECT 88.010 155.190 88.330 155.450 ;
        RECT 90.310 155.390 90.630 155.450 ;
        RECT 92.625 155.390 92.915 155.435 ;
        RECT 90.310 155.250 92.915 155.390 ;
        RECT 90.310 155.190 90.630 155.250 ;
        RECT 92.625 155.205 92.915 155.250 ;
        RECT 95.050 155.390 95.340 155.435 ;
        RECT 99.065 155.390 99.355 155.435 ;
        RECT 101.810 155.390 102.130 155.450 ;
        RECT 95.050 155.250 98.820 155.390 ;
        RECT 95.050 155.205 95.340 155.250 ;
        RECT 45.705 155.050 45.995 155.095 ;
        RECT 41.090 154.910 41.780 155.050 ;
        RECT 42.100 154.910 45.995 155.050 ;
        RECT 41.090 154.850 41.410 154.910 ;
        RECT 34.740 154.570 36.260 154.710 ;
        RECT 36.505 154.525 36.795 154.755 ;
        RECT 38.790 154.510 39.110 154.770 ;
        RECT 40.170 154.710 40.490 154.770 ;
        RECT 42.100 154.710 42.240 154.910 ;
        RECT 45.705 154.865 45.995 154.910 ;
        RECT 46.165 155.050 46.455 155.095 ;
        RECT 48.465 155.050 48.755 155.095 ;
        RECT 46.165 154.910 48.755 155.050 ;
        RECT 46.165 154.865 46.455 154.910 ;
        RECT 48.465 154.865 48.755 154.910 ;
        RECT 64.985 155.050 65.275 155.095 ;
        RECT 66.175 155.050 66.465 155.095 ;
        RECT 68.695 155.050 68.985 155.095 ;
        RECT 64.985 154.910 68.985 155.050 ;
        RECT 64.985 154.865 65.275 154.910 ;
        RECT 66.175 154.865 66.465 154.910 ;
        RECT 68.695 154.865 68.985 154.910 ;
        RECT 73.765 154.865 74.055 155.095 ;
        RECT 75.590 154.850 75.910 155.110 ;
        RECT 84.790 155.050 85.110 155.110 ;
        RECT 88.100 155.050 88.240 155.190 ;
        RECT 84.790 154.910 88.240 155.050 ;
        RECT 84.790 154.850 85.110 154.910 ;
        RECT 94.005 154.865 94.295 155.095 ;
        RECT 40.170 154.570 42.240 154.710 ;
        RECT 43.850 154.710 44.170 154.770 ;
        RECT 51.670 154.710 51.990 154.770 ;
        RECT 43.850 154.570 51.990 154.710 ;
        RECT 40.170 154.510 40.490 154.570 ;
        RECT 43.850 154.510 44.170 154.570 ;
        RECT 51.670 154.510 51.990 154.570 ;
        RECT 64.590 154.710 64.880 154.755 ;
        RECT 66.690 154.710 66.980 154.755 ;
        RECT 68.260 154.710 68.550 154.755 ;
        RECT 64.590 154.570 68.550 154.710 ;
        RECT 64.590 154.525 64.880 154.570 ;
        RECT 66.690 154.525 66.980 154.570 ;
        RECT 68.260 154.525 68.550 154.570 ;
        RECT 72.845 154.710 73.135 154.755 ;
        RECT 75.680 154.710 75.820 154.850 ;
        RECT 91.230 154.710 91.550 154.770 ;
        RECT 72.845 154.570 75.820 154.710 ;
        RECT 84.420 154.570 91.550 154.710 ;
        RECT 94.080 154.710 94.220 154.865 ;
        RECT 94.450 154.850 94.770 155.110 ;
        RECT 95.830 155.050 96.150 155.110 ;
        RECT 98.680 155.050 98.820 155.250 ;
        RECT 99.065 155.250 102.130 155.390 ;
        RECT 99.065 155.205 99.355 155.250 ;
        RECT 101.810 155.190 102.130 155.250 ;
        RECT 107.790 155.390 108.110 155.450 ;
        RECT 108.265 155.390 108.555 155.435 ;
        RECT 107.790 155.250 108.555 155.390 ;
        RECT 107.790 155.190 108.110 155.250 ;
        RECT 108.265 155.205 108.555 155.250 ;
        RECT 109.170 155.190 109.490 155.450 ;
        RECT 105.490 155.050 105.810 155.110 ;
        RECT 109.260 155.050 109.400 155.190 ;
        RECT 95.830 154.910 98.260 155.050 ;
        RECT 98.680 154.910 101.580 155.050 ;
        RECT 95.830 154.850 96.150 154.910 ;
        RECT 94.910 154.710 95.230 154.770 ;
        RECT 94.080 154.570 95.230 154.710 ;
        RECT 72.845 154.525 73.135 154.570 ;
        RECT 17.170 154.370 17.490 154.430 ;
        RECT 18.105 154.370 18.395 154.415 ;
        RECT 17.170 154.230 18.395 154.370 ;
        RECT 17.170 154.170 17.490 154.230 ;
        RECT 18.105 154.185 18.395 154.230 ;
        RECT 31.890 154.170 32.210 154.430 ;
        RECT 53.065 154.370 53.355 154.415 ;
        RECT 53.985 154.370 54.275 154.415 ;
        RECT 53.065 154.230 54.275 154.370 ;
        RECT 53.065 154.185 53.355 154.230 ;
        RECT 53.985 154.185 54.275 154.230 ;
        RECT 59.965 154.370 60.255 154.415 ;
        RECT 61.790 154.370 62.110 154.430 ;
        RECT 59.965 154.230 62.110 154.370 ;
        RECT 59.965 154.185 60.255 154.230 ;
        RECT 61.790 154.170 62.110 154.230 ;
        RECT 73.290 154.170 73.610 154.430 ;
        RECT 73.750 154.370 74.070 154.430 ;
        RECT 75.130 154.370 75.450 154.430 ;
        RECT 84.420 154.415 84.560 154.570 ;
        RECT 91.230 154.510 91.550 154.570 ;
        RECT 94.910 154.510 95.230 154.570 ;
        RECT 73.750 154.230 75.450 154.370 ;
        RECT 73.750 154.170 74.070 154.230 ;
        RECT 75.130 154.170 75.450 154.230 ;
        RECT 84.345 154.185 84.635 154.415 ;
        RECT 88.010 154.170 88.330 154.430 ;
        RECT 96.290 154.370 96.610 154.430 ;
        RECT 97.225 154.370 97.515 154.415 ;
        RECT 96.290 154.230 97.515 154.370 ;
        RECT 98.120 154.370 98.260 154.910 ;
        RECT 101.440 154.430 101.580 154.910 ;
        RECT 105.490 154.910 109.400 155.050 ;
        RECT 105.490 154.850 105.810 154.910 ;
        RECT 100.445 154.370 100.735 154.415 ;
        RECT 98.120 154.230 100.735 154.370 ;
        RECT 96.290 154.170 96.610 154.230 ;
        RECT 97.225 154.185 97.515 154.230 ;
        RECT 100.445 154.185 100.735 154.230 ;
        RECT 101.350 154.170 101.670 154.430 ;
        RECT 108.710 154.170 109.030 154.430 ;
        RECT 11.120 153.550 150.500 154.030 ;
        RECT 26.845 153.350 27.135 153.395 ;
        RECT 30.970 153.350 31.290 153.410 ;
        RECT 26.845 153.210 31.290 153.350 ;
        RECT 26.845 153.165 27.135 153.210 ;
        RECT 30.970 153.150 31.290 153.210 ;
        RECT 42.010 153.150 42.330 153.410 ;
        RECT 42.470 153.150 42.790 153.410 ;
        RECT 42.930 153.150 43.250 153.410 ;
        RECT 44.785 153.350 45.075 153.395 ;
        RECT 45.230 153.350 45.550 153.410 ;
        RECT 44.785 153.210 45.550 153.350 ;
        RECT 44.785 153.165 45.075 153.210 ;
        RECT 45.230 153.150 45.550 153.210 ;
        RECT 55.365 153.350 55.655 153.395 ;
        RECT 56.270 153.350 56.590 153.410 ;
        RECT 55.365 153.210 56.590 153.350 ;
        RECT 55.365 153.165 55.655 153.210 ;
        RECT 56.270 153.150 56.590 153.210 ;
        RECT 84.790 153.150 85.110 153.410 ;
        RECT 92.165 153.165 92.455 153.395 ;
        RECT 95.370 153.350 95.690 153.410 ;
        RECT 95.845 153.350 96.135 153.395 ;
        RECT 95.370 153.210 96.135 153.350 ;
        RECT 16.290 153.010 16.580 153.055 ;
        RECT 18.390 153.010 18.680 153.055 ;
        RECT 19.960 153.010 20.250 153.055 ;
        RECT 16.290 152.870 20.250 153.010 ;
        RECT 16.290 152.825 16.580 152.870 ;
        RECT 18.390 152.825 18.680 152.870 ;
        RECT 19.960 152.825 20.250 152.870 ;
        RECT 22.705 153.010 22.995 153.055 ;
        RECT 30.510 153.010 30.830 153.070 ;
        RECT 22.705 152.870 30.830 153.010 ;
        RECT 22.705 152.825 22.995 152.870 ;
        RECT 30.510 152.810 30.830 152.870 ;
        RECT 16.685 152.670 16.975 152.715 ;
        RECT 17.875 152.670 18.165 152.715 ;
        RECT 20.395 152.670 20.685 152.715 ;
        RECT 16.685 152.530 20.685 152.670 ;
        RECT 16.685 152.485 16.975 152.530 ;
        RECT 17.875 152.485 18.165 152.530 ;
        RECT 20.395 152.485 20.685 152.530 ;
        RECT 24.530 152.670 24.850 152.730 ;
        RECT 25.005 152.670 25.295 152.715 ;
        RECT 24.530 152.530 25.295 152.670 ;
        RECT 30.600 152.670 30.740 152.810 ;
        RECT 30.600 152.530 31.200 152.670 ;
        RECT 24.530 152.470 24.850 152.530 ;
        RECT 25.005 152.485 25.295 152.530 ;
        RECT 15.805 152.330 16.095 152.375 ;
        RECT 16.250 152.330 16.570 152.390 ;
        RECT 17.170 152.375 17.490 152.390 ;
        RECT 17.140 152.330 17.490 152.375 ;
        RECT 15.805 152.190 16.570 152.330 ;
        RECT 16.975 152.190 17.490 152.330 ;
        RECT 15.805 152.145 16.095 152.190 ;
        RECT 16.250 152.130 16.570 152.190 ;
        RECT 17.140 152.145 17.490 152.190 ;
        RECT 25.465 152.330 25.755 152.375 ;
        RECT 27.290 152.330 27.610 152.390 ;
        RECT 31.060 152.375 31.200 152.530 ;
        RECT 25.465 152.190 27.610 152.330 ;
        RECT 25.465 152.145 25.755 152.190 ;
        RECT 17.170 152.130 17.490 152.145 ;
        RECT 27.290 152.130 27.610 152.190 ;
        RECT 30.525 152.145 30.815 152.375 ;
        RECT 30.985 152.145 31.275 152.375 ;
        RECT 29.590 151.450 29.910 151.710 ;
        RECT 30.600 151.650 30.740 152.145 ;
        RECT 32.350 152.130 32.670 152.390 ;
        RECT 35.110 152.130 35.430 152.390 ;
        RECT 40.170 152.330 40.490 152.390 ;
        RECT 41.565 152.330 41.855 152.375 ;
        RECT 42.100 152.330 42.240 153.150 ;
        RECT 40.170 152.190 42.240 152.330 ;
        RECT 43.020 152.330 43.160 153.150 ;
        RECT 51.670 153.010 51.990 153.070 ;
        RECT 60.410 153.010 60.700 153.055 ;
        RECT 61.980 153.010 62.270 153.055 ;
        RECT 64.080 153.010 64.370 153.055 ;
        RECT 51.670 152.870 54.660 153.010 ;
        RECT 51.670 152.810 51.990 152.870 ;
        RECT 51.300 152.530 54.200 152.670 ;
        RECT 51.300 152.390 51.440 152.530 ;
        RECT 44.325 152.330 44.615 152.375 ;
        RECT 45.245 152.330 45.535 152.375 ;
        RECT 43.020 152.190 44.615 152.330 ;
        RECT 40.170 152.130 40.490 152.190 ;
        RECT 41.565 152.145 41.855 152.190 ;
        RECT 44.325 152.145 44.615 152.190 ;
        RECT 44.860 152.190 45.535 152.330 ;
        RECT 31.430 151.790 31.750 152.050 ;
        RECT 35.200 151.990 35.340 152.130 ;
        RECT 36.950 151.990 37.270 152.050 ;
        RECT 38.790 151.990 39.110 152.050 ;
        RECT 41.090 151.990 41.410 152.050 ;
        RECT 42.025 151.990 42.315 152.035 ;
        RECT 35.200 151.850 42.315 151.990 ;
        RECT 36.950 151.790 37.270 151.850 ;
        RECT 38.790 151.790 39.110 151.850 ;
        RECT 41.090 151.790 41.410 151.850 ;
        RECT 42.025 151.805 42.315 151.850 ;
        RECT 42.945 151.990 43.235 152.035 ;
        RECT 43.850 151.990 44.170 152.050 ;
        RECT 42.945 151.850 44.170 151.990 ;
        RECT 42.945 151.805 43.235 151.850 ;
        RECT 43.850 151.790 44.170 151.850 ;
        RECT 44.860 151.710 45.000 152.190 ;
        RECT 45.245 152.145 45.535 152.190 ;
        RECT 51.210 152.130 51.530 152.390 ;
        RECT 52.605 152.145 52.895 152.375 ;
        RECT 52.130 151.990 52.450 152.050 ;
        RECT 52.680 151.990 52.820 152.145 ;
        RECT 53.050 152.130 53.370 152.390 ;
        RECT 54.060 152.375 54.200 152.530 ;
        RECT 54.520 152.375 54.660 152.870 ;
        RECT 60.410 152.870 64.370 153.010 ;
        RECT 60.410 152.825 60.700 152.870 ;
        RECT 61.980 152.825 62.270 152.870 ;
        RECT 64.080 152.825 64.370 152.870 ;
        RECT 80.205 153.010 80.495 153.055 ;
        RECT 80.205 152.870 86.860 153.010 ;
        RECT 80.205 152.825 80.495 152.870 ;
        RECT 59.975 152.670 60.265 152.715 ;
        RECT 62.495 152.670 62.785 152.715 ;
        RECT 63.685 152.670 63.975 152.715 ;
        RECT 59.975 152.530 63.975 152.670 ;
        RECT 59.975 152.485 60.265 152.530 ;
        RECT 62.495 152.485 62.785 152.530 ;
        RECT 63.685 152.485 63.975 152.530 ;
        RECT 67.325 152.670 67.615 152.715 ;
        RECT 67.770 152.670 68.090 152.730 ;
        RECT 67.325 152.530 68.090 152.670 ;
        RECT 67.325 152.485 67.615 152.530 ;
        RECT 67.770 152.470 68.090 152.530 ;
        RECT 78.825 152.670 79.115 152.715 ;
        RECT 82.490 152.670 82.810 152.730 ;
        RECT 78.825 152.530 84.560 152.670 ;
        RECT 78.825 152.485 79.115 152.530 ;
        RECT 82.490 152.470 82.810 152.530 ;
        RECT 53.985 152.145 54.275 152.375 ;
        RECT 54.445 152.145 54.735 152.375 ;
        RECT 61.790 152.330 62.110 152.390 ;
        RECT 63.230 152.330 63.520 152.375 ;
        RECT 61.790 152.190 63.520 152.330 ;
        RECT 61.790 152.130 62.110 152.190 ;
        RECT 63.230 152.145 63.520 152.190 ;
        RECT 64.550 152.130 64.870 152.390 ;
        RECT 66.390 152.130 66.710 152.390 ;
        RECT 72.845 152.145 73.135 152.375 ;
        RECT 73.290 152.330 73.610 152.390 ;
        RECT 73.765 152.330 74.055 152.375 ;
        RECT 73.290 152.190 74.055 152.330 ;
        RECT 52.130 151.850 52.820 151.990 ;
        RECT 72.920 151.990 73.060 152.145 ;
        RECT 73.290 152.130 73.610 152.190 ;
        RECT 73.765 152.145 74.055 152.190 ;
        RECT 74.210 152.130 74.530 152.390 ;
        RECT 74.670 152.330 74.990 152.390 ;
        RECT 76.985 152.330 77.275 152.375 ;
        RECT 74.670 152.190 77.275 152.330 ;
        RECT 74.670 152.130 74.990 152.190 ;
        RECT 76.985 152.145 77.275 152.190 ;
        RECT 78.350 152.130 78.670 152.390 ;
        RECT 84.420 152.375 84.560 152.530 ;
        RECT 83.885 152.330 84.175 152.375 ;
        RECT 83.500 152.190 84.175 152.330 ;
        RECT 76.050 151.990 76.370 152.050 ;
        RECT 72.920 151.850 76.370 151.990 ;
        RECT 52.130 151.790 52.450 151.850 ;
        RECT 73.840 151.710 73.980 151.850 ;
        RECT 76.050 151.790 76.370 151.850 ;
        RECT 83.500 151.710 83.640 152.190 ;
        RECT 83.885 152.145 84.175 152.190 ;
        RECT 84.345 152.145 84.635 152.375 ;
        RECT 85.725 152.330 86.015 152.375 ;
        RECT 86.170 152.330 86.490 152.390 ;
        RECT 85.340 152.190 86.490 152.330 ;
        RECT 86.720 152.330 86.860 152.870 ;
        RECT 87.090 152.810 87.410 153.070 ;
        RECT 92.240 153.010 92.380 153.165 ;
        RECT 95.370 153.150 95.690 153.210 ;
        RECT 95.845 153.165 96.135 153.210 ;
        RECT 96.380 153.210 96.995 153.350 ;
        RECT 96.380 153.010 96.520 153.210 ;
        RECT 92.240 152.870 96.520 153.010 ;
        RECT 96.855 152.670 96.995 153.210 ;
        RECT 98.130 153.150 98.450 153.410 ;
        RECT 102.270 153.350 102.590 153.410 ;
        RECT 108.265 153.350 108.555 153.395 ;
        RECT 102.270 153.210 118.140 153.350 ;
        RECT 102.270 153.150 102.590 153.210 ;
        RECT 108.265 153.165 108.555 153.210 ;
        RECT 111.010 152.810 111.330 153.070 ;
        RECT 113.770 153.010 114.060 153.055 ;
        RECT 115.340 153.010 115.630 153.055 ;
        RECT 117.440 153.010 117.730 153.055 ;
        RECT 113.770 152.870 117.730 153.010 ;
        RECT 113.770 152.825 114.060 152.870 ;
        RECT 115.340 152.825 115.630 152.870 ;
        RECT 117.440 152.825 117.730 152.870 ;
        RECT 118.000 152.715 118.140 153.210 ;
        RECT 113.335 152.670 113.625 152.715 ;
        RECT 115.855 152.670 116.145 152.715 ;
        RECT 117.045 152.670 117.335 152.715 ;
        RECT 96.855 152.530 97.440 152.670 ;
        RECT 87.105 152.330 87.395 152.375 ;
        RECT 91.230 152.330 91.550 152.390 ;
        RECT 86.720 152.190 91.550 152.330 ;
        RECT 85.340 152.035 85.480 152.190 ;
        RECT 85.725 152.145 86.015 152.190 ;
        RECT 86.170 152.130 86.490 152.190 ;
        RECT 87.105 152.145 87.395 152.190 ;
        RECT 91.230 152.130 91.550 152.190 ;
        RECT 93.530 152.130 93.850 152.390 ;
        RECT 93.990 152.130 94.310 152.390 ;
        RECT 94.465 152.145 94.755 152.375 ;
        RECT 95.265 152.330 95.555 152.375 ;
        RECT 95.125 152.300 95.555 152.330 ;
        RECT 95.830 152.300 96.150 152.390 ;
        RECT 95.125 152.160 96.150 152.300 ;
        RECT 95.265 152.145 95.555 152.160 ;
        RECT 85.265 151.805 85.555 152.035 ;
        RECT 31.890 151.650 32.210 151.710 ;
        RECT 30.600 151.510 32.210 151.650 ;
        RECT 31.890 151.450 32.210 151.510 ;
        RECT 44.770 151.450 45.090 151.710 ;
        RECT 57.650 151.450 57.970 151.710 ;
        RECT 65.470 151.450 65.790 151.710 ;
        RECT 71.925 151.650 72.215 151.695 ;
        RECT 72.370 151.650 72.690 151.710 ;
        RECT 71.925 151.510 72.690 151.650 ;
        RECT 71.925 151.465 72.215 151.510 ;
        RECT 72.370 151.450 72.690 151.510 ;
        RECT 73.750 151.450 74.070 151.710 ;
        RECT 76.510 151.450 76.830 151.710 ;
        RECT 83.410 151.650 83.730 151.710 ;
        RECT 86.185 151.650 86.475 151.695 ;
        RECT 83.410 151.510 86.475 151.650 ;
        RECT 94.540 151.650 94.680 152.145 ;
        RECT 95.830 152.130 96.150 152.160 ;
        RECT 96.675 152.330 96.965 152.375 ;
        RECT 96.675 152.145 96.980 152.330 ;
        RECT 96.290 151.650 96.610 151.710 ;
        RECT 94.540 151.510 96.610 151.650 ;
        RECT 96.840 151.650 96.980 152.145 ;
        RECT 97.300 151.990 97.440 152.530 ;
        RECT 113.335 152.530 117.335 152.670 ;
        RECT 113.335 152.485 113.625 152.530 ;
        RECT 115.855 152.485 116.145 152.530 ;
        RECT 117.045 152.485 117.335 152.530 ;
        RECT 117.925 152.670 118.215 152.715 ;
        RECT 118.830 152.670 119.150 152.730 ;
        RECT 122.970 152.670 123.290 152.730 ;
        RECT 117.925 152.530 123.290 152.670 ;
        RECT 117.925 152.485 118.215 152.530 ;
        RECT 118.830 152.470 119.150 152.530 ;
        RECT 122.970 152.470 123.290 152.530 ;
        RECT 97.670 152.130 97.990 152.390 ;
        RECT 100.890 152.330 101.210 152.390 ;
        RECT 101.825 152.330 102.115 152.375 ;
        RECT 100.890 152.190 102.115 152.330 ;
        RECT 100.890 152.130 101.210 152.190 ;
        RECT 101.825 152.145 102.115 152.190 ;
        RECT 99.065 151.990 99.355 152.035 ;
        RECT 97.300 151.850 99.355 151.990 ;
        RECT 99.065 151.805 99.355 151.850 ;
        RECT 109.170 151.990 109.490 152.050 ;
        RECT 116.590 151.990 116.880 152.035 ;
        RECT 109.170 151.850 116.880 151.990 ;
        RECT 109.170 151.790 109.490 151.850 ;
        RECT 116.590 151.805 116.880 151.850 ;
        RECT 97.210 151.650 97.530 151.710 ;
        RECT 96.840 151.510 97.530 151.650 ;
        RECT 83.410 151.450 83.730 151.510 ;
        RECT 86.185 151.465 86.475 151.510 ;
        RECT 96.290 151.450 96.610 151.510 ;
        RECT 97.210 151.450 97.530 151.510 ;
        RECT 11.120 150.830 151.295 151.310 ;
        RECT 19.010 150.430 19.330 150.690 ;
        RECT 29.590 150.630 29.910 150.690 ;
        RECT 22.090 150.490 29.910 150.630 ;
        RECT 19.945 149.950 20.235 149.995 ;
        RECT 22.090 149.950 22.230 150.490 ;
        RECT 29.590 150.430 29.910 150.490 ;
        RECT 40.630 150.630 40.950 150.690 ;
        RECT 41.565 150.630 41.855 150.675 ;
        RECT 40.630 150.490 41.855 150.630 ;
        RECT 40.630 150.430 40.950 150.490 ;
        RECT 41.565 150.445 41.855 150.490 ;
        RECT 74.210 150.630 74.530 150.690 ;
        RECT 74.685 150.630 74.975 150.675 ;
        RECT 74.210 150.490 74.975 150.630 ;
        RECT 74.210 150.430 74.530 150.490 ;
        RECT 74.685 150.445 74.975 150.490 ;
        RECT 76.510 150.430 76.830 150.690 ;
        RECT 94.910 150.430 95.230 150.690 ;
        RECT 96.305 150.630 96.595 150.675 ;
        RECT 98.130 150.630 98.450 150.690 ;
        RECT 96.305 150.490 98.450 150.630 ;
        RECT 96.305 150.445 96.595 150.490 ;
        RECT 98.130 150.430 98.450 150.490 ;
        RECT 108.710 150.430 109.030 150.690 ;
        RECT 109.170 150.430 109.490 150.690 ;
        RECT 111.010 150.430 111.330 150.690 ;
        RECT 39.265 150.290 39.555 150.335 ;
        RECT 39.265 150.150 41.320 150.290 ;
        RECT 39.265 150.105 39.555 150.150 ;
        RECT 19.945 149.810 22.230 149.950 ;
        RECT 30.970 149.950 31.290 150.010 ;
        RECT 33.745 149.950 34.035 149.995 ;
        RECT 35.570 149.950 35.890 150.010 ;
        RECT 38.790 149.995 39.110 150.010 ;
        RECT 38.755 149.950 39.110 149.995 ;
        RECT 30.970 149.810 35.890 149.950 ;
        RECT 38.595 149.810 39.110 149.950 ;
        RECT 19.945 149.765 20.235 149.810 ;
        RECT 30.970 149.750 31.290 149.810 ;
        RECT 33.745 149.765 34.035 149.810 ;
        RECT 35.570 149.750 35.890 149.810 ;
        RECT 38.755 149.765 39.110 149.810 ;
        RECT 39.725 149.950 40.015 149.995 ;
        RECT 40.170 149.950 40.490 150.010 ;
        RECT 41.180 149.995 41.320 150.150 ;
        RECT 39.725 149.810 40.490 149.950 ;
        RECT 39.725 149.765 40.015 149.810 ;
        RECT 38.790 149.750 39.110 149.765 ;
        RECT 20.390 149.610 20.710 149.670 ;
        RECT 20.865 149.610 21.155 149.655 ;
        RECT 34.190 149.610 34.510 149.670 ;
        RECT 39.800 149.610 39.940 149.765 ;
        RECT 40.170 149.750 40.490 149.810 ;
        RECT 41.105 149.765 41.395 149.995 ;
        RECT 42.025 149.950 42.315 149.995 ;
        RECT 45.690 149.950 46.010 150.010 ;
        RECT 53.525 149.950 53.815 149.995 ;
        RECT 42.025 149.810 53.815 149.950 ;
        RECT 42.025 149.765 42.315 149.810 ;
        RECT 45.690 149.750 46.010 149.810 ;
        RECT 53.525 149.765 53.815 149.810 ;
        RECT 75.590 149.750 75.910 150.010 ;
        RECT 76.065 149.950 76.355 149.995 ;
        RECT 76.600 149.950 76.740 150.430 ;
        RECT 95.000 150.290 95.140 150.430 ;
        RECT 108.800 150.290 108.940 150.430 ;
        RECT 95.000 150.150 95.600 150.290 ;
        RECT 76.065 149.810 76.740 149.950 ;
        RECT 76.065 149.765 76.355 149.810 ;
        RECT 93.085 149.765 93.375 149.995 ;
        RECT 93.530 149.950 93.850 150.010 ;
        RECT 93.530 149.810 94.045 149.950 ;
        RECT 20.390 149.470 22.230 149.610 ;
        RECT 20.390 149.410 20.710 149.470 ;
        RECT 20.865 149.425 21.155 149.470 ;
        RECT 22.090 148.930 22.230 149.470 ;
        RECT 34.190 149.470 39.940 149.610 ;
        RECT 34.190 149.410 34.510 149.470 ;
        RECT 51.210 149.410 51.530 149.670 ;
        RECT 51.670 149.610 51.990 149.670 ;
        RECT 53.065 149.610 53.355 149.655 ;
        RECT 51.670 149.470 53.355 149.610 ;
        RECT 51.670 149.410 51.990 149.470 ;
        RECT 53.065 149.425 53.355 149.470 ;
        RECT 74.685 149.610 74.975 149.655 ;
        RECT 79.270 149.610 79.590 149.670 ;
        RECT 74.685 149.470 79.590 149.610 ;
        RECT 74.685 149.425 74.975 149.470 ;
        RECT 79.270 149.410 79.590 149.470 ;
        RECT 27.290 149.270 27.610 149.330 ;
        RECT 31.905 149.270 32.195 149.315 ;
        RECT 27.290 149.130 32.195 149.270 ;
        RECT 27.290 149.070 27.610 149.130 ;
        RECT 31.905 149.085 32.195 149.130 ;
        RECT 56.730 149.270 57.050 149.330 ;
        RECT 61.790 149.270 62.110 149.330 ;
        RECT 56.730 149.130 62.110 149.270 ;
        RECT 93.160 149.270 93.300 149.765 ;
        RECT 93.530 149.750 93.850 149.810 ;
        RECT 94.450 149.750 94.770 150.010 ;
        RECT 95.460 149.995 95.600 150.150 ;
        RECT 106.960 150.150 108.940 150.290 ;
        RECT 111.100 150.290 111.240 150.430 ;
        RECT 113.310 150.290 113.630 150.350 ;
        RECT 120.670 150.290 120.990 150.350 ;
        RECT 111.100 150.150 113.080 150.290 ;
        RECT 94.925 149.765 95.215 149.995 ;
        RECT 95.410 149.765 95.700 149.995 ;
        RECT 98.145 149.950 98.435 149.995 ;
        RECT 95.920 149.810 103.420 149.950 ;
        RECT 95.000 149.610 95.140 149.765 ;
        RECT 95.920 149.610 96.060 149.810 ;
        RECT 98.145 149.765 98.435 149.810 ;
        RECT 95.000 149.470 96.060 149.610 ;
        RECT 96.765 149.610 97.055 149.655 ;
        RECT 99.050 149.610 99.370 149.670 ;
        RECT 96.765 149.470 99.370 149.610 ;
        RECT 96.765 149.425 97.055 149.470 ;
        RECT 99.050 149.410 99.370 149.470 ;
        RECT 101.810 149.410 102.130 149.670 ;
        RECT 103.280 149.655 103.420 149.810 ;
        RECT 103.650 149.750 103.970 150.010 ;
        RECT 105.030 149.950 105.350 150.010 ;
        RECT 106.960 149.995 107.100 150.150 ;
        RECT 105.965 149.950 106.255 149.995 ;
        RECT 105.030 149.810 106.255 149.950 ;
        RECT 105.030 149.750 105.350 149.810 ;
        RECT 105.965 149.765 106.255 149.810 ;
        RECT 106.885 149.765 107.175 149.995 ;
        RECT 107.345 149.765 107.635 149.995 ;
        RECT 103.205 149.610 103.495 149.655 ;
        RECT 103.205 149.470 103.880 149.610 ;
        RECT 103.205 149.425 103.495 149.470 ;
        RECT 97.225 149.270 97.515 149.315 ;
        RECT 93.160 149.130 97.515 149.270 ;
        RECT 56.730 149.070 57.050 149.130 ;
        RECT 61.790 149.070 62.110 149.130 ;
        RECT 97.225 149.085 97.515 149.130 ;
        RECT 103.740 148.990 103.880 149.470 ;
        RECT 107.420 149.270 107.560 149.765 ;
        RECT 107.790 149.750 108.110 150.010 ;
        RECT 108.250 149.950 108.570 150.010 ;
        RECT 109.645 149.950 109.935 149.995 ;
        RECT 108.250 149.810 109.935 149.950 ;
        RECT 108.250 149.750 108.570 149.810 ;
        RECT 109.645 149.765 109.935 149.810 ;
        RECT 111.470 149.750 111.790 150.010 ;
        RECT 112.940 149.995 113.080 150.150 ;
        RECT 113.310 150.150 120.990 150.290 ;
        RECT 113.310 150.090 113.630 150.150 ;
        RECT 120.670 150.090 120.990 150.150 ;
        RECT 112.865 149.765 113.155 149.995 ;
        RECT 114.690 149.750 115.010 150.010 ;
        RECT 122.110 149.950 122.400 149.995 ;
        RECT 115.700 149.810 122.400 149.950 ;
        RECT 107.880 149.610 108.020 149.750 ;
        RECT 110.565 149.610 110.855 149.655 ;
        RECT 113.325 149.610 113.615 149.655 ;
        RECT 107.880 149.470 113.615 149.610 ;
        RECT 110.565 149.425 110.855 149.470 ;
        RECT 113.325 149.425 113.615 149.470 ;
        RECT 115.700 149.315 115.840 149.810 ;
        RECT 122.110 149.765 122.400 149.810 ;
        RECT 122.970 149.950 123.290 150.010 ;
        RECT 123.445 149.950 123.735 149.995 ;
        RECT 122.970 149.810 123.735 149.950 ;
        RECT 122.970 149.750 123.290 149.810 ;
        RECT 123.445 149.765 123.735 149.810 ;
        RECT 118.855 149.610 119.145 149.655 ;
        RECT 121.375 149.610 121.665 149.655 ;
        RECT 122.565 149.610 122.855 149.655 ;
        RECT 118.855 149.470 122.855 149.610 ;
        RECT 118.855 149.425 119.145 149.470 ;
        RECT 121.375 149.425 121.665 149.470 ;
        RECT 122.565 149.425 122.855 149.470 ;
        RECT 107.420 149.130 109.860 149.270 ;
        RECT 109.720 148.990 109.860 149.130 ;
        RECT 115.625 149.085 115.915 149.315 ;
        RECT 119.290 149.270 119.580 149.315 ;
        RECT 120.860 149.270 121.150 149.315 ;
        RECT 122.960 149.270 123.250 149.315 ;
        RECT 119.290 149.130 123.250 149.270 ;
        RECT 119.290 149.085 119.580 149.130 ;
        RECT 120.860 149.085 121.150 149.130 ;
        RECT 122.960 149.085 123.250 149.130 ;
        RECT 24.990 148.930 25.310 148.990 ;
        RECT 37.410 148.930 37.730 148.990 ;
        RECT 22.090 148.790 37.730 148.930 ;
        RECT 24.990 148.730 25.310 148.790 ;
        RECT 37.410 148.730 37.730 148.790 ;
        RECT 54.445 148.930 54.735 148.975 ;
        RECT 68.230 148.930 68.550 148.990 ;
        RECT 54.445 148.790 68.550 148.930 ;
        RECT 54.445 148.745 54.735 148.790 ;
        RECT 68.230 148.730 68.550 148.790 ;
        RECT 94.910 148.930 95.230 148.990 ;
        RECT 97.685 148.930 97.975 148.975 ;
        RECT 94.910 148.790 97.975 148.930 ;
        RECT 94.910 148.730 95.230 148.790 ;
        RECT 97.685 148.745 97.975 148.790 ;
        RECT 103.650 148.730 103.970 148.990 ;
        RECT 109.630 148.730 109.950 148.990 ;
        RECT 110.090 148.730 110.410 148.990 ;
        RECT 116.530 148.730 116.850 148.990 ;
        RECT 11.120 148.110 150.500 148.590 ;
        RECT 30.510 147.910 30.830 147.970 ;
        RECT 18.640 147.770 30.830 147.910 ;
        RECT 18.640 147.275 18.780 147.770 ;
        RECT 23.240 147.615 23.380 147.770 ;
        RECT 30.510 147.710 30.830 147.770 ;
        RECT 45.690 147.710 46.010 147.970 ;
        RECT 51.210 147.910 51.530 147.970 ;
        RECT 51.685 147.910 51.975 147.955 ;
        RECT 52.605 147.910 52.895 147.955 ;
        RECT 51.210 147.770 52.895 147.910 ;
        RECT 51.210 147.710 51.530 147.770 ;
        RECT 51.685 147.725 51.975 147.770 ;
        RECT 52.605 147.725 52.895 147.770 ;
        RECT 60.500 147.770 66.115 147.910 ;
        RECT 20.405 147.385 20.695 147.615 ;
        RECT 23.165 147.385 23.455 147.615 ;
        RECT 23.625 147.570 23.915 147.615 ;
        RECT 24.070 147.570 24.390 147.630 ;
        RECT 23.625 147.430 25.680 147.570 ;
        RECT 23.625 147.385 23.915 147.430 ;
        RECT 18.565 147.045 18.855 147.275 ;
        RECT 20.480 146.890 20.620 147.385 ;
        RECT 24.070 147.370 24.390 147.430 ;
        RECT 20.865 147.230 21.155 147.275 ;
        RECT 20.865 147.090 24.760 147.230 ;
        RECT 20.865 147.045 21.155 147.090 ;
        RECT 21.325 146.890 21.615 146.935 ;
        RECT 23.610 146.890 23.930 146.950 ;
        RECT 24.620 146.935 24.760 147.090 ;
        RECT 25.540 146.935 25.680 147.430 ;
        RECT 26.385 147.230 26.675 147.275 ;
        RECT 29.145 147.230 29.435 147.275 ;
        RECT 26.385 147.090 29.435 147.230 ;
        RECT 30.600 147.230 30.740 147.710 ;
        RECT 38.370 147.570 38.660 147.615 ;
        RECT 40.470 147.570 40.760 147.615 ;
        RECT 42.040 147.570 42.330 147.615 ;
        RECT 38.370 147.430 42.330 147.570 ;
        RECT 38.370 147.385 38.660 147.430 ;
        RECT 40.470 147.385 40.760 147.430 ;
        RECT 42.040 147.385 42.330 147.430 ;
        RECT 44.785 147.385 45.075 147.615 ;
        RECT 54.445 147.570 54.735 147.615 ;
        RECT 60.500 147.570 60.640 147.770 ;
        RECT 54.445 147.430 60.640 147.570 ;
        RECT 54.445 147.385 54.735 147.430 ;
        RECT 38.765 147.230 39.055 147.275 ;
        RECT 39.955 147.230 40.245 147.275 ;
        RECT 42.475 147.230 42.765 147.275 ;
        RECT 30.600 147.090 32.580 147.230 ;
        RECT 26.385 147.045 26.675 147.090 ;
        RECT 29.145 147.045 29.435 147.090 ;
        RECT 20.480 146.750 23.930 146.890 ;
        RECT 21.325 146.705 21.615 146.750 ;
        RECT 23.610 146.690 23.930 146.750 ;
        RECT 24.545 146.705 24.835 146.935 ;
        RECT 25.465 146.705 25.755 146.935 ;
        RECT 26.830 146.690 27.150 146.950 ;
        RECT 27.305 146.705 27.595 146.935 ;
        RECT 25.005 146.550 25.295 146.595 ;
        RECT 27.380 146.550 27.520 146.705 ;
        RECT 27.750 146.690 28.070 146.950 ;
        RECT 30.065 146.890 30.355 146.935 ;
        RECT 30.970 146.890 31.290 146.950 ;
        RECT 32.440 146.935 32.580 147.090 ;
        RECT 38.765 147.090 42.765 147.230 ;
        RECT 38.765 147.045 39.055 147.090 ;
        RECT 39.955 147.045 40.245 147.090 ;
        RECT 42.475 147.045 42.765 147.090 ;
        RECT 30.065 146.750 31.290 146.890 ;
        RECT 30.065 146.705 30.355 146.750 ;
        RECT 30.970 146.690 31.290 146.750 ;
        RECT 31.445 146.705 31.735 146.935 ;
        RECT 32.365 146.705 32.655 146.935 ;
        RECT 25.005 146.410 27.520 146.550 ;
        RECT 31.520 146.550 31.660 146.705 ;
        RECT 34.190 146.690 34.510 146.950 ;
        RECT 37.870 146.690 38.190 146.950 ;
        RECT 44.860 146.890 45.000 147.385 ;
        RECT 53.050 147.230 53.370 147.290 ;
        RECT 50.840 147.090 56.500 147.230 ;
        RECT 50.840 146.935 50.980 147.090 ;
        RECT 53.050 147.030 53.370 147.090 ;
        RECT 56.360 146.950 56.500 147.090 ;
        RECT 57.190 147.030 57.510 147.290 ;
        RECT 58.585 147.230 58.875 147.275 ;
        RECT 58.585 147.090 59.260 147.230 ;
        RECT 58.585 147.045 58.875 147.090 ;
        RECT 47.545 146.890 47.835 146.935 ;
        RECT 48.005 146.890 48.295 146.935 ;
        RECT 44.860 146.750 48.295 146.890 ;
        RECT 47.545 146.705 47.835 146.750 ;
        RECT 48.005 146.705 48.295 146.750 ;
        RECT 50.765 146.705 51.055 146.935 ;
        RECT 51.685 146.705 51.975 146.935 ;
        RECT 52.145 146.890 52.435 146.935 ;
        RECT 52.145 146.750 53.280 146.890 ;
        RECT 52.145 146.705 52.435 146.750 ;
        RECT 34.280 146.550 34.420 146.690 ;
        RECT 31.520 146.410 34.420 146.550 ;
        RECT 39.220 146.550 39.510 146.595 ;
        RECT 39.710 146.550 40.030 146.610 ;
        RECT 39.220 146.410 40.030 146.550 ;
        RECT 25.005 146.365 25.295 146.410 ;
        RECT 25.540 146.270 25.680 146.410 ;
        RECT 39.220 146.365 39.510 146.410 ;
        RECT 39.710 146.350 40.030 146.410 ;
        RECT 40.170 146.550 40.490 146.610 ;
        RECT 46.625 146.550 46.915 146.595 ;
        RECT 40.170 146.410 46.915 146.550 ;
        RECT 51.760 146.550 51.900 146.705 ;
        RECT 51.760 146.410 52.360 146.550 ;
        RECT 40.170 146.350 40.490 146.410 ;
        RECT 46.625 146.365 46.915 146.410 ;
        RECT 52.220 146.270 52.360 146.410 ;
        RECT 53.140 146.270 53.280 146.750 ;
        RECT 53.525 146.705 53.815 146.935 ;
        RECT 53.600 146.550 53.740 146.705 ;
        RECT 56.270 146.690 56.590 146.950 ;
        RECT 56.745 146.890 57.035 146.935 ;
        RECT 58.110 146.890 58.430 146.950 ;
        RECT 56.745 146.750 58.430 146.890 ;
        RECT 56.745 146.705 57.035 146.750 ;
        RECT 58.110 146.690 58.430 146.750 ;
        RECT 59.120 146.550 59.260 147.090 ;
        RECT 59.505 146.890 59.795 146.935 ;
        RECT 60.500 146.890 60.640 147.430 ;
        RECT 60.885 147.385 61.175 147.615 ;
        RECT 61.790 147.570 62.110 147.630 ;
        RECT 61.790 147.430 62.940 147.570 ;
        RECT 60.960 147.230 61.100 147.385 ;
        RECT 61.790 147.370 62.110 147.430 ;
        RECT 62.265 147.230 62.555 147.275 ;
        RECT 60.960 147.090 62.555 147.230 ;
        RECT 62.800 147.230 62.940 147.430 ;
        RECT 64.565 147.230 64.855 147.275 ;
        RECT 65.010 147.230 65.330 147.290 ;
        RECT 62.800 147.090 65.330 147.230 ;
        RECT 65.975 147.230 66.115 147.770 ;
        RECT 68.690 147.710 69.010 147.970 ;
        RECT 104.145 147.910 104.435 147.955 ;
        RECT 105.065 147.910 105.355 147.955 ;
        RECT 104.145 147.770 105.355 147.910 ;
        RECT 104.145 147.725 104.435 147.770 ;
        RECT 105.065 147.725 105.355 147.770 ;
        RECT 108.250 147.710 108.570 147.970 ;
        RECT 114.690 147.910 115.010 147.970 ;
        RECT 116.545 147.910 116.835 147.955 ;
        RECT 114.690 147.770 116.835 147.910 ;
        RECT 114.690 147.710 115.010 147.770 ;
        RECT 116.545 147.725 116.835 147.770 ;
        RECT 77.890 147.570 78.210 147.630 ;
        RECT 88.485 147.570 88.775 147.615 ;
        RECT 94.450 147.570 94.770 147.630 ;
        RECT 102.270 147.570 102.590 147.630 ;
        RECT 109.630 147.570 109.950 147.630 ;
        RECT 77.890 147.430 88.240 147.570 ;
        RECT 77.890 147.370 78.210 147.430 ;
        RECT 66.405 147.230 66.695 147.275 ;
        RECT 65.975 147.090 66.695 147.230 ;
        RECT 62.265 147.045 62.555 147.090 ;
        RECT 64.565 147.045 64.855 147.090 ;
        RECT 65.010 147.030 65.330 147.090 ;
        RECT 66.405 147.045 66.695 147.090 ;
        RECT 67.310 147.030 67.630 147.290 ;
        RECT 79.745 147.230 80.035 147.275 ;
        RECT 86.185 147.230 86.475 147.275 ;
        RECT 71.080 147.090 80.035 147.230 ;
        RECT 59.505 146.750 60.640 146.890 ;
        RECT 59.505 146.705 59.795 146.750 ;
        RECT 62.725 146.705 63.015 146.935 ;
        RECT 64.105 146.705 64.395 146.935 ;
        RECT 65.950 146.890 66.240 146.935 ;
        RECT 65.950 146.750 66.620 146.890 ;
        RECT 65.950 146.705 66.240 146.750 ;
        RECT 60.885 146.550 61.175 146.595 ;
        RECT 53.600 146.410 56.960 146.550 ;
        RECT 59.120 146.410 62.020 146.550 ;
        RECT 56.820 146.270 56.960 146.410 ;
        RECT 60.885 146.365 61.175 146.410 ;
        RECT 61.880 146.270 62.020 146.410 ;
        RECT 25.450 146.010 25.770 146.270 ;
        RECT 28.685 146.210 28.975 146.255 ;
        RECT 38.790 146.210 39.110 146.270 ;
        RECT 28.685 146.070 39.110 146.210 ;
        RECT 28.685 146.025 28.975 146.070 ;
        RECT 38.790 146.010 39.110 146.070 ;
        RECT 47.070 146.210 47.390 146.270 ;
        RECT 48.925 146.210 49.215 146.255 ;
        RECT 47.070 146.070 49.215 146.210 ;
        RECT 47.070 146.010 47.390 146.070 ;
        RECT 48.925 146.025 49.215 146.070 ;
        RECT 52.130 146.010 52.450 146.270 ;
        RECT 53.050 146.010 53.370 146.270 ;
        RECT 56.730 146.010 57.050 146.270 ;
        RECT 59.950 146.010 60.270 146.270 ;
        RECT 61.330 146.010 61.650 146.270 ;
        RECT 61.790 146.010 62.110 146.270 ;
        RECT 62.800 146.210 62.940 146.705 ;
        RECT 64.180 146.550 64.320 146.705 ;
        RECT 64.180 146.410 66.160 146.550 ;
        RECT 66.020 146.270 66.160 146.410 ;
        RECT 65.025 146.210 65.315 146.255 ;
        RECT 62.800 146.070 65.315 146.210 ;
        RECT 65.025 146.025 65.315 146.070 ;
        RECT 65.930 146.010 66.250 146.270 ;
        RECT 66.480 146.210 66.620 146.750 ;
        RECT 66.850 146.690 67.170 146.950 ;
        RECT 68.230 146.890 68.550 146.950 ;
        RECT 69.585 146.890 69.875 146.985 ;
        RECT 68.230 146.755 69.875 146.890 ;
        RECT 68.230 146.750 69.840 146.755 ;
        RECT 68.230 146.690 68.550 146.750 ;
        RECT 70.070 146.690 70.390 146.950 ;
        RECT 71.080 146.935 71.220 147.090 ;
        RECT 79.745 147.045 80.035 147.090 ;
        RECT 81.200 147.090 86.475 147.230 ;
        RECT 71.005 146.705 71.295 146.935 ;
        RECT 71.465 146.890 71.755 146.935 ;
        RECT 78.810 146.890 79.130 146.950 ;
        RECT 81.200 146.935 81.340 147.090 ;
        RECT 86.185 147.045 86.475 147.090 ;
        RECT 81.125 146.890 81.415 146.935 ;
        RECT 71.465 146.750 78.580 146.890 ;
        RECT 71.465 146.705 71.755 146.750 ;
        RECT 77.430 146.350 77.750 146.610 ;
        RECT 78.440 146.270 78.580 146.750 ;
        RECT 78.810 146.750 81.415 146.890 ;
        RECT 78.810 146.690 79.130 146.750 ;
        RECT 81.125 146.705 81.415 146.750 ;
        RECT 81.585 146.705 81.875 146.935 ;
        RECT 82.045 146.890 82.335 146.935 ;
        RECT 82.490 146.890 82.810 146.950 ;
        RECT 82.045 146.750 82.810 146.890 ;
        RECT 82.045 146.705 82.335 146.750 ;
        RECT 81.660 146.550 81.800 146.705 ;
        RECT 82.490 146.690 82.810 146.750 ;
        RECT 82.965 146.890 83.255 146.935 ;
        RECT 83.410 146.890 83.730 146.950 ;
        RECT 82.965 146.750 83.730 146.890 ;
        RECT 82.965 146.705 83.255 146.750 ;
        RECT 83.410 146.690 83.730 146.750 ;
        RECT 86.630 146.690 86.950 146.950 ;
        RECT 88.100 146.890 88.240 147.430 ;
        RECT 88.485 147.430 94.770 147.570 ;
        RECT 88.485 147.385 88.775 147.430 ;
        RECT 94.450 147.370 94.770 147.430 ;
        RECT 99.600 147.430 103.420 147.570 ;
        RECT 99.600 146.935 99.740 147.430 ;
        RECT 102.270 147.370 102.590 147.430 ;
        RECT 99.970 147.230 100.290 147.290 ;
        RECT 102.745 147.230 103.035 147.275 ;
        RECT 99.970 147.090 103.035 147.230 ;
        RECT 99.970 147.030 100.290 147.090 ;
        RECT 102.745 147.045 103.035 147.090 ;
        RECT 99.525 146.890 99.815 146.935 ;
        RECT 88.100 146.750 99.815 146.890 ;
        RECT 99.525 146.705 99.815 146.750 ;
        RECT 88.930 146.550 89.250 146.610 ;
        RECT 93.530 146.550 93.850 146.610 ;
        RECT 81.660 146.410 93.850 146.550 ;
        RECT 102.820 146.550 102.960 147.045 ;
        RECT 103.280 146.935 103.420 147.430 ;
        RECT 109.630 147.430 115.380 147.570 ;
        RECT 109.630 147.370 109.950 147.430 ;
        RECT 107.345 147.230 107.635 147.275 ;
        RECT 111.025 147.230 111.315 147.275 ;
        RECT 111.470 147.230 111.790 147.290 ;
        RECT 107.345 147.090 111.790 147.230 ;
        RECT 107.345 147.045 107.635 147.090 ;
        RECT 111.025 147.045 111.315 147.090 ;
        RECT 111.470 147.030 111.790 147.090 ;
        RECT 112.020 147.090 114.920 147.230 ;
        RECT 103.205 146.890 103.495 146.935 ;
        RECT 107.805 146.890 108.095 146.935 ;
        RECT 103.205 146.750 108.095 146.890 ;
        RECT 103.205 146.705 103.495 146.750 ;
        RECT 107.805 146.705 108.095 146.750 ;
        RECT 108.725 146.705 109.015 146.935 ;
        RECT 108.800 146.550 108.940 146.705 ;
        RECT 110.550 146.690 110.870 146.950 ;
        RECT 112.020 146.890 112.160 147.090 ;
        RECT 111.100 146.750 112.160 146.890 ;
        RECT 111.100 146.550 111.240 146.750 ;
        RECT 113.310 146.690 113.630 146.950 ;
        RECT 114.245 146.890 114.535 146.935 ;
        RECT 113.860 146.750 114.535 146.890 ;
        RECT 102.820 146.410 111.240 146.550 ;
        RECT 111.470 146.550 111.790 146.610 ;
        RECT 113.400 146.550 113.540 146.690 ;
        RECT 111.470 146.410 113.540 146.550 ;
        RECT 88.930 146.350 89.250 146.410 ;
        RECT 93.530 146.350 93.850 146.410 ;
        RECT 111.470 146.350 111.790 146.410 ;
        RECT 66.850 146.210 67.170 146.270 ;
        RECT 66.480 146.070 67.170 146.210 ;
        RECT 66.850 146.010 67.170 146.070 ;
        RECT 77.890 146.010 78.210 146.270 ;
        RECT 78.350 146.010 78.670 146.270 ;
        RECT 79.270 146.210 79.590 146.270 ;
        RECT 99.970 146.210 100.290 146.270 ;
        RECT 79.270 146.070 100.290 146.210 ;
        RECT 79.270 146.010 79.590 146.070 ;
        RECT 99.970 146.010 100.290 146.070 ;
        RECT 112.405 146.210 112.695 146.255 ;
        RECT 113.860 146.210 114.000 146.750 ;
        RECT 114.245 146.705 114.535 146.750 ;
        RECT 114.780 146.595 114.920 147.090 ;
        RECT 115.240 146.935 115.380 147.430 ;
        RECT 116.085 147.385 116.375 147.615 ;
        RECT 115.165 146.705 115.455 146.935 ;
        RECT 116.160 146.890 116.300 147.385 ;
        RECT 117.465 146.890 117.755 146.935 ;
        RECT 116.160 146.750 117.755 146.890 ;
        RECT 117.465 146.705 117.755 146.750 ;
        RECT 117.910 146.890 118.230 146.950 ;
        RECT 119.290 146.890 119.610 146.950 ;
        RECT 117.910 146.750 119.610 146.890 ;
        RECT 117.910 146.690 118.230 146.750 ;
        RECT 119.290 146.690 119.610 146.750 ;
        RECT 114.705 146.550 114.995 146.595 ;
        RECT 116.530 146.550 116.850 146.610 ;
        RECT 114.705 146.410 116.850 146.550 ;
        RECT 114.705 146.365 114.995 146.410 ;
        RECT 116.530 146.350 116.850 146.410 ;
        RECT 112.405 146.070 114.000 146.210 ;
        RECT 112.405 146.025 112.695 146.070 ;
        RECT 11.120 145.390 151.295 145.870 ;
        RECT 24.070 144.990 24.390 145.250 ;
        RECT 25.450 144.990 25.770 145.250 ;
        RECT 39.710 144.990 40.030 145.250 ;
        RECT 57.650 144.990 57.970 145.250 ;
        RECT 61.330 144.990 61.650 145.250 ;
        RECT 65.010 145.190 65.330 145.250 ;
        RECT 70.070 145.190 70.390 145.250 ;
        RECT 70.545 145.190 70.835 145.235 ;
        RECT 65.010 145.050 70.835 145.190 ;
        RECT 65.010 144.990 65.330 145.050 ;
        RECT 70.070 144.990 70.390 145.050 ;
        RECT 70.545 145.005 70.835 145.050 ;
        RECT 77.430 145.190 77.750 145.250 ;
        RECT 77.905 145.190 78.195 145.235 ;
        RECT 77.430 145.050 78.195 145.190 ;
        RECT 77.430 144.990 77.750 145.050 ;
        RECT 77.905 145.005 78.195 145.050 ;
        RECT 78.350 145.190 78.670 145.250 ;
        RECT 79.745 145.190 80.035 145.235 ;
        RECT 78.350 145.050 80.035 145.190 ;
        RECT 78.350 144.990 78.670 145.050 ;
        RECT 79.745 145.005 80.035 145.050 ;
        RECT 86.170 144.990 86.490 145.250 ;
        RECT 88.930 144.990 89.250 145.250 ;
        RECT 94.910 144.990 95.230 145.250 ;
        RECT 24.160 144.555 24.300 144.990 ;
        RECT 25.540 144.555 25.680 144.990 ;
        RECT 35.570 144.850 35.890 144.910 ;
        RECT 57.740 144.850 57.880 144.990 ;
        RECT 35.570 144.710 57.880 144.850 ;
        RECT 35.570 144.650 35.890 144.710 ;
        RECT 24.085 144.325 24.375 144.555 ;
        RECT 25.005 144.325 25.295 144.555 ;
        RECT 25.465 144.325 25.755 144.555 ;
        RECT 24.530 144.170 24.850 144.230 ;
        RECT 24.160 144.030 24.850 144.170 ;
        RECT 24.160 143.875 24.300 144.030 ;
        RECT 24.530 143.970 24.850 144.030 ;
        RECT 24.085 143.645 24.375 143.875 ;
        RECT 25.080 143.830 25.220 144.325 ;
        RECT 25.540 144.170 25.680 144.325 ;
        RECT 27.290 144.310 27.610 144.570 ;
        RECT 38.330 144.310 38.650 144.570 ;
        RECT 39.265 144.510 39.555 144.555 ;
        RECT 40.645 144.510 40.935 144.555 ;
        RECT 39.265 144.370 40.935 144.510 ;
        RECT 39.265 144.325 39.555 144.370 ;
        RECT 40.645 144.325 40.935 144.370 ;
        RECT 47.070 144.510 47.390 144.570 ;
        RECT 50.765 144.510 51.055 144.555 ;
        RECT 47.070 144.370 51.055 144.510 ;
        RECT 47.070 144.310 47.390 144.370 ;
        RECT 50.765 144.325 51.055 144.370 ;
        RECT 51.670 144.310 51.990 144.570 ;
        RECT 61.420 144.555 61.560 144.990 ;
        RECT 61.790 144.850 62.110 144.910 ;
        RECT 66.850 144.850 67.170 144.910 ;
        RECT 72.370 144.895 72.690 144.910 ;
        RECT 61.790 144.710 67.170 144.850 ;
        RECT 61.790 144.650 62.110 144.710 ;
        RECT 66.850 144.650 67.170 144.710 ;
        RECT 72.340 144.850 72.690 144.895 ;
        RECT 83.885 144.850 84.175 144.895 ;
        RECT 86.945 144.850 87.235 144.895 ;
        RECT 72.340 144.710 72.840 144.850 ;
        RECT 78.900 144.710 87.235 144.850 ;
        RECT 72.340 144.665 72.690 144.710 ;
        RECT 72.370 144.650 72.690 144.665 ;
        RECT 78.900 144.570 79.040 144.710 ;
        RECT 83.885 144.665 84.175 144.710 ;
        RECT 86.945 144.665 87.235 144.710 ;
        RECT 88.025 144.850 88.315 144.895 ;
        RECT 102.745 144.850 103.035 144.895 ;
        RECT 103.190 144.850 103.510 144.910 ;
        RECT 88.025 144.710 93.760 144.850 ;
        RECT 88.025 144.665 88.315 144.710 ;
        RECT 65.010 144.555 65.330 144.570 ;
        RECT 61.360 144.325 61.650 144.555 ;
        RECT 64.980 144.325 65.330 144.555 ;
        RECT 65.010 144.310 65.330 144.325 ;
        RECT 78.810 144.310 79.130 144.570 ;
        RECT 79.745 144.510 80.035 144.555 ;
        RECT 82.030 144.510 82.350 144.570 ;
        RECT 90.860 144.555 91.000 144.710 ;
        RECT 79.745 144.370 82.350 144.510 ;
        RECT 79.745 144.325 80.035 144.370 ;
        RECT 82.030 144.310 82.350 144.370 ;
        RECT 82.965 144.325 83.255 144.555 ;
        RECT 89.865 144.510 90.155 144.555 ;
        RECT 89.865 144.370 90.265 144.510 ;
        RECT 89.865 144.325 90.155 144.370 ;
        RECT 90.785 144.325 91.075 144.555 ;
        RECT 26.845 144.170 27.135 144.215 ;
        RECT 25.540 144.030 27.135 144.170 ;
        RECT 26.845 143.985 27.135 144.030 ;
        RECT 27.380 143.830 27.520 144.310 ;
        RECT 29.145 144.170 29.435 144.215 ;
        RECT 31.430 144.170 31.750 144.230 ;
        RECT 29.145 144.030 31.750 144.170 ;
        RECT 29.145 143.985 29.435 144.030 ;
        RECT 31.430 143.970 31.750 144.030 ;
        RECT 37.410 143.970 37.730 144.230 ;
        RECT 48.910 144.170 49.230 144.230 ;
        RECT 51.760 144.170 51.900 144.310 ;
        RECT 48.910 144.030 51.900 144.170 ;
        RECT 53.050 144.170 53.370 144.230 ;
        RECT 58.110 144.170 58.430 144.230 ;
        RECT 53.050 144.030 58.430 144.170 ;
        RECT 48.910 143.970 49.230 144.030 ;
        RECT 53.050 143.970 53.370 144.030 ;
        RECT 58.110 143.970 58.430 144.030 ;
        RECT 60.425 144.170 60.715 144.215 ;
        RECT 60.425 144.030 61.100 144.170 ;
        RECT 60.425 143.985 60.715 144.030 ;
        RECT 25.080 143.690 27.520 143.830 ;
        RECT 37.500 143.490 37.640 143.970 ;
        RECT 51.685 143.830 51.975 143.875 ;
        RECT 56.730 143.830 57.050 143.890 ;
        RECT 59.030 143.830 59.350 143.890 ;
        RECT 51.685 143.690 59.350 143.830 ;
        RECT 51.685 143.645 51.975 143.690 ;
        RECT 56.730 143.630 57.050 143.690 ;
        RECT 59.030 143.630 59.350 143.690 ;
        RECT 60.960 143.550 61.100 144.030 ;
        RECT 63.645 143.985 63.935 144.215 ;
        RECT 64.525 144.170 64.815 144.215 ;
        RECT 65.715 144.170 66.005 144.215 ;
        RECT 68.235 144.170 68.525 144.215 ;
        RECT 71.005 144.170 71.295 144.215 ;
        RECT 64.525 144.030 68.525 144.170 ;
        RECT 64.525 143.985 64.815 144.030 ;
        RECT 65.715 143.985 66.005 144.030 ;
        RECT 68.235 143.985 68.525 144.030 ;
        RECT 70.390 144.030 71.295 144.170 ;
        RECT 60.870 143.490 61.190 143.550 ;
        RECT 37.500 143.350 61.190 143.490 ;
        RECT 60.870 143.290 61.190 143.350 ;
        RECT 61.790 143.490 62.110 143.550 ;
        RECT 62.265 143.490 62.555 143.535 ;
        RECT 61.790 143.350 62.555 143.490 ;
        RECT 63.720 143.490 63.860 143.985 ;
        RECT 64.130 143.830 64.420 143.875 ;
        RECT 66.230 143.830 66.520 143.875 ;
        RECT 67.800 143.830 68.090 143.875 ;
        RECT 64.130 143.690 68.090 143.830 ;
        RECT 64.130 143.645 64.420 143.690 ;
        RECT 66.230 143.645 66.520 143.690 ;
        RECT 67.800 143.645 68.090 143.690 ;
        RECT 64.550 143.490 64.870 143.550 ;
        RECT 70.390 143.490 70.530 144.030 ;
        RECT 71.005 143.985 71.295 144.030 ;
        RECT 71.885 144.170 72.175 144.215 ;
        RECT 73.075 144.170 73.365 144.215 ;
        RECT 75.595 144.170 75.885 144.215 ;
        RECT 71.885 144.030 75.885 144.170 ;
        RECT 71.885 143.985 72.175 144.030 ;
        RECT 73.075 143.985 73.365 144.030 ;
        RECT 75.595 143.985 75.885 144.030 ;
        RECT 78.350 143.970 78.670 144.230 ;
        RECT 83.040 144.170 83.180 144.325 ;
        RECT 89.940 144.170 90.080 144.325 ;
        RECT 93.070 144.310 93.390 144.570 ;
        RECT 93.620 144.510 93.760 144.710 ;
        RECT 102.745 144.710 103.510 144.850 ;
        RECT 102.745 144.665 103.035 144.710 ;
        RECT 103.190 144.650 103.510 144.710 ;
        RECT 103.650 144.510 103.970 144.570 ;
        RECT 93.620 144.370 103.970 144.510 ;
        RECT 103.650 144.310 103.970 144.370 ;
        RECT 115.625 144.510 115.915 144.555 ;
        RECT 116.530 144.510 116.850 144.570 ;
        RECT 115.625 144.370 116.850 144.510 ;
        RECT 115.625 144.325 115.915 144.370 ;
        RECT 116.530 144.310 116.850 144.370 ;
        RECT 92.625 144.170 92.915 144.215 ;
        RECT 83.040 144.030 92.915 144.170 ;
        RECT 71.490 143.830 71.780 143.875 ;
        RECT 73.590 143.830 73.880 143.875 ;
        RECT 75.160 143.830 75.450 143.875 ;
        RECT 71.490 143.690 75.450 143.830 ;
        RECT 71.490 143.645 71.780 143.690 ;
        RECT 73.590 143.645 73.880 143.690 ;
        RECT 75.160 143.645 75.450 143.690 ;
        RECT 63.720 143.350 70.530 143.490 ;
        RECT 78.440 143.490 78.580 143.970 ;
        RECT 79.285 143.830 79.575 143.875 ;
        RECT 82.950 143.830 83.270 143.890 ;
        RECT 79.285 143.690 83.270 143.830 ;
        RECT 79.285 143.645 79.575 143.690 ;
        RECT 82.950 143.630 83.270 143.690 ;
        RECT 87.640 143.550 87.780 144.030 ;
        RECT 92.625 143.985 92.915 144.030 ;
        RECT 102.270 143.830 102.590 143.890 ;
        RECT 104.125 143.830 104.415 143.875 ;
        RECT 102.270 143.690 104.415 143.830 ;
        RECT 102.270 143.630 102.590 143.690 ;
        RECT 104.125 143.645 104.415 143.690 ;
        RECT 83.410 143.490 83.730 143.550 ;
        RECT 78.440 143.350 83.730 143.490 ;
        RECT 61.790 143.290 62.110 143.350 ;
        RECT 62.265 143.305 62.555 143.350 ;
        RECT 64.550 143.290 64.870 143.350 ;
        RECT 83.410 143.290 83.730 143.350 ;
        RECT 87.105 143.490 87.395 143.535 ;
        RECT 87.550 143.490 87.870 143.550 ;
        RECT 87.105 143.350 87.870 143.490 ;
        RECT 87.105 143.305 87.395 143.350 ;
        RECT 87.550 143.290 87.870 143.350 ;
        RECT 105.030 143.290 105.350 143.550 ;
        RECT 116.545 143.490 116.835 143.535 ;
        RECT 119.750 143.490 120.070 143.550 ;
        RECT 116.545 143.350 120.070 143.490 ;
        RECT 116.545 143.305 116.835 143.350 ;
        RECT 119.750 143.290 120.070 143.350 ;
        RECT 11.120 142.670 150.500 143.150 ;
        RECT 38.330 142.270 38.650 142.530 ;
        RECT 47.070 142.470 47.390 142.530 ;
        RECT 42.560 142.330 47.390 142.470 ;
        RECT 42.560 141.835 42.700 142.330 ;
        RECT 45.780 142.175 45.920 142.330 ;
        RECT 47.070 142.270 47.390 142.330 ;
        RECT 53.050 142.270 53.370 142.530 ;
        RECT 65.010 142.470 65.330 142.530 ;
        RECT 65.485 142.470 65.775 142.515 ;
        RECT 65.010 142.330 65.775 142.470 ;
        RECT 65.010 142.270 65.330 142.330 ;
        RECT 65.485 142.285 65.775 142.330 ;
        RECT 105.030 142.270 105.350 142.530 ;
        RECT 43.865 142.130 44.155 142.175 ;
        RECT 43.865 141.990 45.460 142.130 ;
        RECT 43.865 141.945 44.155 141.990 ;
        RECT 42.485 141.790 42.775 141.835 ;
        RECT 37.040 141.650 42.775 141.790 ;
        RECT 45.320 141.790 45.460 141.990 ;
        RECT 45.705 141.945 45.995 142.175 ;
        RECT 53.140 142.130 53.280 142.270 ;
        RECT 46.240 141.990 53.280 142.130 ;
        RECT 60.870 142.130 61.190 142.190 ;
        RECT 60.870 141.990 70.530 142.130 ;
        RECT 46.240 141.790 46.380 141.990 ;
        RECT 45.320 141.650 46.380 141.790 ;
        RECT 37.040 141.510 37.180 141.650 ;
        RECT 42.485 141.605 42.775 141.650 ;
        RECT 18.550 141.250 18.870 141.510 ;
        RECT 28.225 141.265 28.515 141.495 ;
        RECT 28.670 141.450 28.990 141.510 ;
        RECT 29.145 141.450 29.435 141.495 ;
        RECT 30.970 141.450 31.290 141.510 ;
        RECT 28.670 141.310 31.290 141.450 ;
        RECT 24.530 141.110 24.850 141.170 ;
        RECT 28.300 141.110 28.440 141.265 ;
        RECT 28.670 141.250 28.990 141.310 ;
        RECT 29.145 141.265 29.435 141.310 ;
        RECT 30.970 141.250 31.290 141.310 ;
        RECT 32.350 141.450 32.670 141.510 ;
        RECT 35.585 141.450 35.875 141.495 ;
        RECT 32.350 141.310 35.875 141.450 ;
        RECT 32.350 141.250 32.670 141.310 ;
        RECT 35.585 141.265 35.875 141.310 ;
        RECT 36.950 141.250 37.270 141.510 ;
        RECT 47.620 141.495 47.760 141.990 ;
        RECT 60.870 141.930 61.190 141.990 ;
        RECT 65.470 141.790 65.790 141.850 ;
        RECT 48.080 141.650 65.790 141.790 ;
        RECT 70.390 141.790 70.530 141.990 ;
        RECT 94.450 141.790 94.770 141.850 ;
        RECT 70.390 141.650 94.770 141.790 ;
        RECT 37.425 141.450 37.715 141.495 ;
        RECT 37.425 141.310 47.300 141.450 ;
        RECT 37.425 141.265 37.715 141.310 ;
        RECT 33.730 141.110 34.050 141.170 ;
        RECT 24.530 140.970 34.050 141.110 ;
        RECT 24.530 140.910 24.850 140.970 ;
        RECT 33.730 140.910 34.050 140.970 ;
        RECT 36.490 140.910 36.810 141.170 ;
        RECT 17.170 140.770 17.490 140.830 ;
        RECT 17.645 140.770 17.935 140.815 ;
        RECT 17.170 140.630 17.935 140.770 ;
        RECT 17.170 140.570 17.490 140.630 ;
        RECT 17.645 140.585 17.935 140.630 ;
        RECT 29.130 140.570 29.450 140.830 ;
        RECT 30.970 140.770 31.290 140.830 ;
        RECT 31.890 140.770 32.210 140.830 ;
        RECT 37.500 140.770 37.640 141.265 ;
        RECT 44.310 141.110 44.630 141.170 ;
        RECT 47.160 141.110 47.300 141.310 ;
        RECT 47.545 141.265 47.835 141.495 ;
        RECT 48.080 141.110 48.220 141.650 ;
        RECT 65.470 141.590 65.790 141.650 ;
        RECT 94.450 141.590 94.770 141.650 ;
        RECT 103.190 141.790 103.510 141.850 ;
        RECT 104.125 141.790 104.415 141.835 ;
        RECT 103.190 141.650 104.415 141.790 ;
        RECT 103.190 141.590 103.510 141.650 ;
        RECT 104.125 141.605 104.415 141.650 ;
        RECT 52.605 141.450 52.895 141.495 ;
        RECT 57.650 141.450 57.970 141.510 ;
        RECT 52.605 141.310 57.970 141.450 ;
        RECT 52.605 141.265 52.895 141.310 ;
        RECT 57.650 141.250 57.970 141.310 ;
        RECT 61.790 141.450 62.110 141.510 ;
        RECT 66.405 141.450 66.695 141.495 ;
        RECT 61.790 141.310 66.695 141.450 ;
        RECT 61.790 141.250 62.110 141.310 ;
        RECT 66.405 141.265 66.695 141.310 ;
        RECT 76.510 141.250 76.830 141.510 ;
        RECT 77.430 141.250 77.750 141.510 ;
        RECT 99.970 141.450 100.290 141.510 ;
        RECT 102.745 141.450 103.035 141.495 ;
        RECT 99.970 141.310 103.035 141.450 ;
        RECT 99.970 141.250 100.290 141.310 ;
        RECT 102.745 141.265 103.035 141.310 ;
        RECT 103.650 141.250 103.970 141.510 ;
        RECT 44.310 140.970 45.460 141.110 ;
        RECT 47.160 140.970 48.220 141.110 ;
        RECT 104.200 141.110 104.340 141.605 ;
        RECT 105.120 141.495 105.260 142.270 ;
        RECT 114.245 142.130 114.535 142.175 ;
        RECT 112.480 141.990 114.535 142.130 ;
        RECT 107.345 141.790 107.635 141.835 ;
        RECT 105.580 141.650 107.635 141.790 ;
        RECT 105.580 141.510 105.720 141.650 ;
        RECT 107.345 141.605 107.635 141.650 ;
        RECT 109.645 141.790 109.935 141.835 ;
        RECT 109.645 141.650 112.160 141.790 ;
        RECT 109.645 141.605 109.935 141.650 ;
        RECT 105.045 141.265 105.335 141.495 ;
        RECT 105.490 141.250 105.810 141.510 ;
        RECT 105.950 141.250 106.270 141.510 ;
        RECT 107.790 141.450 108.110 141.510 ;
        RECT 110.090 141.450 110.410 141.510 ;
        RECT 107.790 141.310 110.410 141.450 ;
        RECT 107.790 141.250 108.110 141.310 ;
        RECT 110.090 141.250 110.410 141.310 ;
        RECT 111.025 141.450 111.315 141.495 ;
        RECT 111.470 141.450 111.790 141.510 ;
        RECT 112.020 141.495 112.160 141.650 ;
        RECT 112.480 141.495 112.620 141.990 ;
        RECT 114.245 141.945 114.535 141.990 ;
        RECT 116.990 142.130 117.280 142.175 ;
        RECT 118.560 142.130 118.850 142.175 ;
        RECT 120.660 142.130 120.950 142.175 ;
        RECT 116.990 141.990 120.950 142.130 ;
        RECT 116.990 141.945 117.280 141.990 ;
        RECT 118.560 141.945 118.850 141.990 ;
        RECT 120.660 141.945 120.950 141.990 ;
        RECT 116.555 141.790 116.845 141.835 ;
        RECT 119.075 141.790 119.365 141.835 ;
        RECT 120.265 141.790 120.555 141.835 ;
        RECT 116.555 141.650 120.555 141.790 ;
        RECT 116.555 141.605 116.845 141.650 ;
        RECT 119.075 141.605 119.365 141.650 ;
        RECT 120.265 141.605 120.555 141.650 ;
        RECT 111.025 141.310 111.790 141.450 ;
        RECT 111.025 141.265 111.315 141.310 ;
        RECT 111.470 141.250 111.790 141.310 ;
        RECT 111.945 141.265 112.235 141.495 ;
        RECT 112.405 141.265 112.695 141.495 ;
        RECT 112.865 141.265 113.155 141.495 ;
        RECT 121.145 141.450 121.435 141.495 ;
        RECT 118.920 141.310 121.435 141.450 ;
        RECT 112.480 141.110 112.620 141.265 ;
        RECT 104.200 140.970 112.620 141.110 ;
        RECT 44.310 140.910 44.630 140.970 ;
        RECT 30.970 140.630 37.640 140.770 ;
        RECT 30.970 140.570 31.290 140.630 ;
        RECT 31.890 140.570 32.210 140.630 ;
        RECT 44.770 140.570 45.090 140.830 ;
        RECT 45.320 140.815 45.460 140.970 ;
        RECT 45.245 140.585 45.535 140.815 ;
        RECT 47.070 140.770 47.390 140.830 ;
        RECT 75.590 140.770 75.910 140.830 ;
        RECT 47.070 140.630 75.910 140.770 ;
        RECT 47.070 140.570 47.390 140.630 ;
        RECT 75.590 140.570 75.910 140.630 ;
        RECT 76.970 140.570 77.290 140.830 ;
        RECT 101.825 140.770 102.115 140.815 ;
        RECT 102.730 140.770 103.050 140.830 ;
        RECT 101.825 140.630 103.050 140.770 ;
        RECT 101.825 140.585 102.115 140.630 ;
        RECT 102.730 140.570 103.050 140.630 ;
        RECT 105.490 140.570 105.810 140.830 ;
        RECT 108.250 140.770 108.570 140.830 ;
        RECT 109.630 140.770 109.950 140.830 ;
        RECT 112.940 140.770 113.080 141.265 ;
        RECT 118.370 141.110 118.690 141.170 ;
        RECT 118.920 141.110 119.060 141.310 ;
        RECT 121.145 141.265 121.435 141.310 ;
        RECT 118.370 140.970 119.060 141.110 ;
        RECT 119.750 141.155 120.070 141.170 ;
        RECT 118.370 140.910 118.690 140.970 ;
        RECT 119.750 140.925 120.100 141.155 ;
        RECT 119.750 140.910 120.070 140.925 ;
        RECT 108.250 140.630 113.080 140.770 ;
        RECT 108.250 140.570 108.570 140.630 ;
        RECT 109.630 140.570 109.950 140.630 ;
        RECT 113.770 140.570 114.090 140.830 ;
        RECT 11.120 139.950 151.295 140.430 ;
        RECT 37.870 139.750 38.190 139.810 ;
        RECT 38.805 139.750 39.095 139.795 ;
        RECT 47.070 139.750 47.390 139.810 ;
        RECT 22.090 139.610 39.095 139.750 ;
        RECT 16.250 139.410 16.570 139.470 ;
        RECT 22.090 139.410 22.230 139.610 ;
        RECT 37.870 139.550 38.190 139.610 ;
        RECT 38.805 139.565 39.095 139.610 ;
        RECT 45.780 139.610 47.390 139.750 ;
        RECT 16.250 139.270 22.230 139.410 ;
        RECT 23.610 139.410 23.930 139.470 ;
        RECT 28.670 139.410 28.990 139.470 ;
        RECT 23.610 139.270 28.990 139.410 ;
        RECT 16.250 139.210 16.570 139.270 ;
        RECT 23.610 139.210 23.930 139.270 ;
        RECT 15.805 139.070 16.095 139.115 ;
        RECT 16.340 139.070 16.480 139.210 ;
        RECT 17.170 139.115 17.490 139.130 ;
        RECT 24.160 139.115 24.300 139.270 ;
        RECT 28.670 139.210 28.990 139.270 ;
        RECT 29.130 139.410 29.450 139.470 ;
        RECT 29.605 139.410 29.895 139.455 ;
        RECT 29.130 139.270 29.895 139.410 ;
        RECT 29.130 139.210 29.450 139.270 ;
        RECT 29.605 139.225 29.895 139.270 ;
        RECT 31.445 139.410 31.735 139.455 ;
        RECT 33.730 139.410 34.050 139.470 ;
        RECT 31.445 139.270 34.050 139.410 ;
        RECT 31.445 139.225 31.735 139.270 ;
        RECT 33.730 139.210 34.050 139.270 ;
        RECT 17.140 139.070 17.490 139.115 ;
        RECT 15.805 138.930 16.480 139.070 ;
        RECT 16.975 138.930 17.490 139.070 ;
        RECT 15.805 138.885 16.095 138.930 ;
        RECT 17.140 138.885 17.490 138.930 ;
        RECT 24.085 138.885 24.375 139.115 ;
        RECT 27.765 139.070 28.055 139.115 ;
        RECT 26.000 138.930 28.055 139.070 ;
        RECT 17.170 138.870 17.490 138.885 ;
        RECT 16.685 138.730 16.975 138.775 ;
        RECT 17.875 138.730 18.165 138.775 ;
        RECT 20.395 138.730 20.685 138.775 ;
        RECT 16.685 138.590 20.685 138.730 ;
        RECT 16.685 138.545 16.975 138.590 ;
        RECT 17.875 138.545 18.165 138.590 ;
        RECT 20.395 138.545 20.685 138.590 ;
        RECT 24.530 138.530 24.850 138.790 ;
        RECT 16.290 138.390 16.580 138.435 ;
        RECT 18.390 138.390 18.680 138.435 ;
        RECT 19.960 138.390 20.250 138.435 ;
        RECT 16.290 138.250 20.250 138.390 ;
        RECT 16.290 138.205 16.580 138.250 ;
        RECT 18.390 138.205 18.680 138.250 ;
        RECT 19.960 138.205 20.250 138.250 ;
        RECT 22.705 138.390 22.995 138.435 ;
        RECT 24.620 138.390 24.760 138.530 ;
        RECT 26.000 138.450 26.140 138.930 ;
        RECT 27.765 138.885 28.055 138.930 ;
        RECT 30.970 138.870 31.290 139.130 ;
        RECT 31.890 138.870 32.210 139.130 ;
        RECT 32.810 139.070 33.130 139.130 ;
        RECT 45.780 139.070 45.920 139.610 ;
        RECT 47.070 139.550 47.390 139.610 ;
        RECT 58.585 139.750 58.875 139.795 ;
        RECT 59.950 139.750 60.270 139.810 ;
        RECT 58.585 139.610 60.270 139.750 ;
        RECT 58.585 139.565 58.875 139.610 ;
        RECT 59.950 139.550 60.270 139.610 ;
        RECT 60.410 139.750 60.730 139.810 ;
        RECT 61.345 139.750 61.635 139.795 ;
        RECT 60.410 139.610 61.635 139.750 ;
        RECT 60.410 139.550 60.730 139.610 ;
        RECT 61.345 139.565 61.635 139.610 ;
        RECT 75.605 139.565 75.895 139.795 ;
        RECT 79.270 139.750 79.590 139.810 ;
        RECT 87.105 139.750 87.395 139.795 ;
        RECT 89.850 139.750 90.170 139.810 ;
        RECT 105.030 139.750 105.350 139.810 ;
        RECT 79.270 139.610 82.720 139.750 ;
        RECT 46.165 139.410 46.455 139.455 ;
        RECT 47.545 139.410 47.835 139.455 ;
        RECT 49.370 139.410 49.690 139.470 ;
        RECT 46.165 139.270 49.690 139.410 ;
        RECT 46.165 139.225 46.455 139.270 ;
        RECT 47.545 139.225 47.835 139.270 ;
        RECT 49.370 139.210 49.690 139.270 ;
        RECT 56.285 139.410 56.575 139.455 ;
        RECT 64.550 139.410 64.870 139.470 ;
        RECT 56.285 139.270 64.870 139.410 ;
        RECT 56.285 139.225 56.575 139.270 ;
        RECT 64.550 139.210 64.870 139.270 ;
        RECT 65.470 139.210 65.790 139.470 ;
        RECT 75.680 139.410 75.820 139.565 ;
        RECT 79.270 139.550 79.590 139.610 ;
        RECT 76.510 139.410 76.830 139.470 ;
        RECT 76.985 139.410 77.275 139.455 ;
        RECT 75.680 139.270 77.275 139.410 ;
        RECT 76.510 139.210 76.830 139.270 ;
        RECT 76.985 139.225 77.275 139.270 ;
        RECT 77.430 139.410 77.750 139.470 ;
        RECT 77.905 139.410 78.195 139.455 ;
        RECT 78.825 139.410 79.115 139.455 ;
        RECT 77.430 139.270 79.115 139.410 ;
        RECT 77.430 139.210 77.750 139.270 ;
        RECT 77.905 139.225 78.195 139.270 ;
        RECT 78.825 139.225 79.115 139.270 ;
        RECT 81.355 139.410 81.645 139.455 ;
        RECT 82.030 139.410 82.350 139.470 ;
        RECT 81.355 139.270 82.350 139.410 ;
        RECT 81.355 139.225 81.645 139.270 ;
        RECT 82.030 139.210 82.350 139.270 ;
        RECT 32.810 138.930 45.920 139.070 ;
        RECT 32.810 138.870 33.130 138.930 ;
        RECT 57.650 138.870 57.970 139.130 ;
        RECT 59.030 138.870 59.350 139.130 ;
        RECT 59.505 138.885 59.795 139.115 ;
        RECT 73.765 139.070 74.055 139.115 ;
        RECT 79.270 139.070 79.590 139.130 ;
        RECT 79.745 139.070 80.035 139.115 ;
        RECT 73.765 138.930 79.040 139.070 ;
        RECT 73.765 138.885 74.055 138.930 ;
        RECT 28.685 138.730 28.975 138.775 ;
        RECT 31.430 138.730 31.750 138.790 ;
        RECT 28.685 138.590 31.750 138.730 ;
        RECT 28.685 138.545 28.975 138.590 ;
        RECT 31.430 138.530 31.750 138.590 ;
        RECT 53.510 138.730 53.830 138.790 ;
        RECT 55.350 138.730 55.670 138.790 ;
        RECT 59.580 138.730 59.720 138.885 ;
        RECT 53.510 138.590 59.720 138.730 ;
        RECT 53.510 138.530 53.830 138.590 ;
        RECT 55.350 138.530 55.670 138.590 ;
        RECT 59.950 138.530 60.270 138.790 ;
        RECT 73.305 138.730 73.595 138.775 ;
        RECT 78.350 138.730 78.670 138.790 ;
        RECT 73.305 138.590 78.670 138.730 ;
        RECT 73.305 138.545 73.595 138.590 ;
        RECT 22.705 138.250 24.760 138.390 ;
        RECT 22.705 138.205 22.995 138.250 ;
        RECT 25.910 138.190 26.230 138.450 ;
        RECT 27.290 138.390 27.610 138.450 ;
        RECT 27.765 138.390 28.055 138.435 ;
        RECT 27.290 138.250 28.055 138.390 ;
        RECT 27.290 138.190 27.610 138.250 ;
        RECT 27.765 138.205 28.055 138.250 ;
        RECT 73.380 138.110 73.520 138.545 ;
        RECT 78.350 138.530 78.670 138.590 ;
        RECT 77.890 138.390 78.210 138.450 ;
        RECT 78.900 138.390 79.040 138.930 ;
        RECT 79.270 138.930 80.035 139.070 ;
        RECT 79.270 138.870 79.590 138.930 ;
        RECT 79.745 138.885 80.035 138.930 ;
        RECT 80.190 138.870 80.510 139.130 ;
        RECT 80.665 138.885 80.955 139.115 ;
        RECT 82.580 139.070 82.720 139.610 ;
        RECT 87.105 139.610 90.170 139.750 ;
        RECT 87.105 139.565 87.395 139.610 ;
        RECT 89.850 139.550 90.170 139.610 ;
        RECT 101.440 139.610 105.350 139.750 ;
        RECT 86.170 139.410 86.490 139.470 ;
        RECT 96.750 139.410 97.070 139.470 ;
        RECT 97.270 139.410 97.560 139.455 ;
        RECT 84.420 139.270 85.940 139.410 ;
        RECT 84.420 139.130 84.560 139.270 ;
        RECT 84.330 139.070 84.650 139.130 ;
        RECT 82.580 138.930 84.650 139.070 ;
        RECT 77.890 138.250 79.040 138.390 ;
        RECT 77.890 138.190 78.210 138.250 ;
        RECT 25.450 138.050 25.770 138.110 ;
        RECT 30.065 138.050 30.355 138.095 ;
        RECT 25.450 137.910 30.355 138.050 ;
        RECT 25.450 137.850 25.770 137.910 ;
        RECT 30.065 137.865 30.355 137.910 ;
        RECT 56.730 137.850 57.050 138.110 ;
        RECT 60.410 137.850 60.730 138.110 ;
        RECT 66.850 138.050 67.170 138.110 ;
        RECT 72.830 138.050 73.150 138.110 ;
        RECT 66.850 137.910 73.150 138.050 ;
        RECT 66.850 137.850 67.170 137.910 ;
        RECT 72.830 137.850 73.150 137.910 ;
        RECT 73.290 137.850 73.610 138.110 ;
        RECT 76.050 137.850 76.370 138.110 ;
        RECT 80.740 138.050 80.880 138.885 ;
        RECT 82.045 138.730 82.335 138.775 ;
        RECT 82.580 138.730 82.720 138.930 ;
        RECT 84.330 138.870 84.650 138.930 ;
        RECT 85.265 138.885 85.555 139.115 ;
        RECT 85.800 139.070 85.940 139.270 ;
        RECT 86.170 139.270 89.160 139.410 ;
        RECT 86.170 139.210 86.490 139.270 ;
        RECT 86.645 139.070 86.935 139.115 ;
        RECT 85.800 138.930 86.935 139.070 ;
        RECT 86.645 138.885 86.935 138.930 ;
        RECT 82.045 138.590 82.720 138.730 ;
        RECT 85.340 138.730 85.480 138.885 ;
        RECT 87.550 138.870 87.870 139.130 ;
        RECT 89.020 139.115 89.160 139.270 ;
        RECT 89.480 139.270 96.520 139.410 ;
        RECT 89.480 139.130 89.620 139.270 ;
        RECT 88.945 138.885 89.235 139.115 ;
        RECT 89.390 138.870 89.710 139.130 ;
        RECT 89.850 138.870 90.170 139.130 ;
        RECT 96.380 139.070 96.520 139.270 ;
        RECT 96.750 139.270 97.560 139.410 ;
        RECT 96.750 139.210 97.070 139.270 ;
        RECT 97.270 139.225 97.560 139.270 ;
        RECT 101.440 139.070 101.580 139.610 ;
        RECT 105.030 139.550 105.350 139.610 ;
        RECT 105.950 139.550 106.270 139.810 ;
        RECT 107.345 139.750 107.635 139.795 ;
        RECT 107.790 139.750 108.110 139.810 ;
        RECT 107.345 139.610 108.110 139.750 ;
        RECT 107.345 139.565 107.635 139.610 ;
        RECT 107.790 139.550 108.110 139.610 ;
        RECT 113.770 139.550 114.090 139.810 ;
        RECT 116.530 139.550 116.850 139.810 ;
        RECT 102.270 139.410 102.590 139.470 ;
        RECT 103.665 139.410 103.955 139.455 ;
        RECT 102.270 139.270 103.955 139.410 ;
        RECT 106.040 139.410 106.180 139.550 ;
        RECT 106.425 139.410 106.715 139.455 ;
        RECT 106.040 139.270 106.715 139.410 ;
        RECT 107.880 139.410 108.020 139.550 ;
        RECT 107.880 139.270 108.480 139.410 ;
        RECT 102.270 139.210 102.590 139.270 ;
        RECT 103.665 139.225 103.955 139.270 ;
        RECT 106.425 139.225 106.715 139.270 ;
        RECT 96.380 138.930 101.580 139.070 ;
        RECT 101.825 139.070 102.115 139.115 ;
        RECT 105.490 139.070 105.810 139.130 ;
        RECT 107.805 139.070 108.095 139.115 ;
        RECT 101.825 138.930 108.095 139.070 ;
        RECT 101.825 138.885 102.115 138.930 ;
        RECT 105.490 138.870 105.810 138.930 ;
        RECT 107.805 138.885 108.095 138.930 ;
        RECT 87.640 138.730 87.780 138.870 ;
        RECT 94.015 138.730 94.305 138.775 ;
        RECT 96.535 138.730 96.825 138.775 ;
        RECT 97.725 138.730 98.015 138.775 ;
        RECT 85.340 138.590 91.920 138.730 ;
        RECT 82.045 138.545 82.335 138.590 ;
        RECT 81.110 138.390 81.430 138.450 ;
        RECT 81.110 138.250 89.160 138.390 ;
        RECT 81.110 138.190 81.430 138.250 ;
        RECT 89.020 138.110 89.160 138.250 ;
        RECT 82.490 138.050 82.810 138.110 ;
        RECT 80.740 137.910 82.810 138.050 ;
        RECT 82.490 137.850 82.810 137.910 ;
        RECT 83.410 138.050 83.730 138.110 ;
        RECT 86.170 138.050 86.490 138.110 ;
        RECT 83.410 137.910 86.490 138.050 ;
        RECT 83.410 137.850 83.730 137.910 ;
        RECT 86.170 137.850 86.490 137.910 ;
        RECT 88.930 137.850 89.250 138.110 ;
        RECT 91.780 138.095 91.920 138.590 ;
        RECT 94.015 138.590 98.015 138.730 ;
        RECT 94.015 138.545 94.305 138.590 ;
        RECT 96.535 138.545 96.825 138.590 ;
        RECT 97.725 138.545 98.015 138.590 ;
        RECT 98.590 138.530 98.910 138.790 ;
        RECT 101.350 138.530 101.670 138.790 ;
        RECT 102.285 138.545 102.575 138.775 ;
        RECT 92.150 138.390 92.470 138.450 ;
        RECT 94.450 138.390 94.740 138.435 ;
        RECT 96.020 138.390 96.310 138.435 ;
        RECT 98.120 138.390 98.410 138.435 ;
        RECT 92.150 138.250 94.220 138.390 ;
        RECT 92.150 138.190 92.470 138.250 ;
        RECT 91.705 138.050 91.995 138.095 ;
        RECT 93.530 138.050 93.850 138.110 ;
        RECT 91.705 137.910 93.850 138.050 ;
        RECT 94.080 138.050 94.220 138.250 ;
        RECT 94.450 138.250 98.410 138.390 ;
        RECT 94.450 138.205 94.740 138.250 ;
        RECT 96.020 138.205 96.310 138.250 ;
        RECT 98.120 138.205 98.410 138.250 ;
        RECT 100.445 138.050 100.735 138.095 ;
        RECT 94.080 137.910 100.735 138.050 ;
        RECT 102.360 138.050 102.500 138.545 ;
        RECT 102.730 138.530 103.050 138.790 ;
        RECT 103.190 138.390 103.510 138.450 ;
        RECT 105.045 138.390 105.335 138.435 ;
        RECT 108.340 138.390 108.480 139.270 ;
        RECT 113.860 139.070 114.000 139.550 ;
        RECT 115.625 139.070 115.915 139.115 ;
        RECT 113.860 138.930 115.915 139.070 ;
        RECT 115.625 138.885 115.915 138.930 ;
        RECT 110.090 138.730 110.410 138.790 ;
        RECT 114.705 138.730 114.995 138.775 ;
        RECT 117.910 138.730 118.230 138.790 ;
        RECT 110.090 138.590 118.230 138.730 ;
        RECT 110.090 138.530 110.410 138.590 ;
        RECT 114.705 138.545 114.995 138.590 ;
        RECT 117.910 138.530 118.230 138.590 ;
        RECT 103.190 138.250 105.335 138.390 ;
        RECT 103.190 138.190 103.510 138.250 ;
        RECT 105.045 138.205 105.335 138.250 ;
        RECT 105.580 138.250 108.480 138.390 ;
        RECT 105.580 138.050 105.720 138.250 ;
        RECT 102.360 137.910 105.720 138.050 ;
        RECT 91.705 137.865 91.995 137.910 ;
        RECT 93.530 137.850 93.850 137.910 ;
        RECT 100.445 137.865 100.735 137.910 ;
        RECT 106.410 137.850 106.730 138.110 ;
        RECT 11.120 137.230 150.500 137.710 ;
        RECT 18.550 136.830 18.870 137.090 ;
        RECT 25.450 137.030 25.770 137.090 ;
        RECT 22.090 136.890 25.770 137.030 ;
        RECT 22.090 136.350 22.230 136.890 ;
        RECT 25.450 136.830 25.770 136.890 ;
        RECT 25.910 136.830 26.230 137.090 ;
        RECT 31.890 137.030 32.210 137.090 ;
        RECT 29.220 136.890 32.210 137.030 ;
        RECT 19.560 136.210 22.230 136.350 ;
        RECT 26.000 136.350 26.140 136.830 ;
        RECT 29.220 136.735 29.360 136.890 ;
        RECT 31.890 136.830 32.210 136.890 ;
        RECT 36.490 137.030 36.810 137.090 ;
        RECT 37.425 137.030 37.715 137.075 ;
        RECT 36.490 136.890 37.715 137.030 ;
        RECT 36.490 136.830 36.810 136.890 ;
        RECT 37.425 136.845 37.715 136.890 ;
        RECT 46.625 137.030 46.915 137.075 ;
        RECT 47.070 137.030 47.390 137.090 ;
        RECT 46.625 136.890 47.390 137.030 ;
        RECT 46.625 136.845 46.915 136.890 ;
        RECT 47.070 136.830 47.390 136.890 ;
        RECT 47.545 137.030 47.835 137.075 ;
        RECT 47.545 136.890 53.280 137.030 ;
        RECT 47.545 136.845 47.835 136.890 ;
        RECT 29.145 136.505 29.435 136.735 ;
        RECT 48.005 136.690 48.295 136.735 ;
        RECT 41.640 136.550 48.295 136.690 ;
        RECT 53.140 136.690 53.280 136.890 ;
        RECT 53.510 136.830 53.830 137.090 ;
        RECT 57.190 137.030 57.510 137.090 ;
        RECT 59.965 137.030 60.255 137.075 ;
        RECT 60.870 137.030 61.190 137.090 ;
        RECT 57.190 136.890 61.190 137.030 ;
        RECT 57.190 136.830 57.510 136.890 ;
        RECT 59.965 136.845 60.255 136.890 ;
        RECT 60.870 136.830 61.190 136.890 ;
        RECT 62.265 136.845 62.555 137.075 ;
        RECT 67.770 137.030 68.090 137.090 ;
        RECT 71.465 137.030 71.755 137.075 ;
        RECT 73.290 137.030 73.610 137.090 ;
        RECT 67.770 136.890 69.840 137.030 ;
        RECT 60.410 136.690 60.730 136.750 ;
        RECT 62.340 136.690 62.480 136.845 ;
        RECT 67.770 136.830 68.090 136.890 ;
        RECT 53.140 136.550 62.480 136.690 ;
        RECT 65.050 136.690 65.340 136.735 ;
        RECT 67.150 136.690 67.440 136.735 ;
        RECT 68.720 136.690 69.010 136.735 ;
        RECT 65.050 136.550 69.010 136.690 ;
        RECT 26.845 136.350 27.135 136.395 ;
        RECT 26.000 136.210 27.135 136.350 ;
        RECT 19.560 136.055 19.700 136.210 ;
        RECT 26.845 136.165 27.135 136.210 ;
        RECT 39.725 136.350 40.015 136.395 ;
        RECT 41.640 136.350 41.780 136.550 ;
        RECT 48.005 136.505 48.295 136.550 ;
        RECT 60.410 136.490 60.730 136.550 ;
        RECT 65.050 136.505 65.340 136.550 ;
        RECT 67.150 136.505 67.440 136.550 ;
        RECT 68.720 136.505 69.010 136.550 ;
        RECT 39.725 136.210 41.780 136.350 ;
        RECT 39.725 136.165 40.015 136.210 ;
        RECT 19.485 135.825 19.775 136.055 ;
        RECT 20.390 135.810 20.710 136.070 ;
        RECT 27.290 135.810 27.610 136.070 ;
        RECT 38.790 136.010 39.110 136.070 ;
        RECT 41.640 136.055 41.780 136.210 ;
        RECT 44.310 136.350 44.630 136.410 ;
        RECT 45.705 136.350 45.995 136.395 ;
        RECT 44.310 136.210 48.220 136.350 ;
        RECT 44.310 136.150 44.630 136.210 ;
        RECT 45.705 136.165 45.995 136.210 ;
        RECT 39.265 136.010 39.555 136.055 ;
        RECT 38.790 135.870 39.555 136.010 ;
        RECT 38.790 135.810 39.110 135.870 ;
        RECT 39.265 135.825 39.555 135.870 ;
        RECT 41.565 135.825 41.855 136.055 ;
        RECT 42.945 136.010 43.235 136.055 ;
        RECT 44.400 136.010 44.540 136.150 ;
        RECT 42.945 135.870 44.540 136.010 ;
        RECT 42.945 135.825 43.235 135.870 ;
        RECT 39.340 135.670 39.480 135.825 ;
        RECT 44.770 135.810 45.090 136.070 ;
        RECT 48.080 136.055 48.220 136.210 ;
        RECT 52.130 136.150 52.450 136.410 ;
        RECT 58.585 136.165 58.875 136.395 ;
        RECT 59.030 136.350 59.350 136.410 ;
        RECT 62.250 136.350 62.570 136.410 ;
        RECT 59.030 136.210 62.570 136.350 ;
        RECT 46.625 135.825 46.915 136.055 ;
        RECT 48.005 135.825 48.295 136.055 ;
        RECT 48.925 135.825 49.215 136.055 ;
        RECT 51.670 136.010 51.990 136.070 ;
        RECT 53.050 136.010 53.370 136.070 ;
        RECT 51.670 135.870 53.370 136.010 ;
        RECT 42.025 135.670 42.315 135.715 ;
        RECT 44.325 135.670 44.615 135.715 ;
        RECT 39.340 135.530 44.615 135.670 ;
        RECT 44.860 135.670 45.000 135.810 ;
        RECT 46.700 135.670 46.840 135.825 ;
        RECT 49.000 135.670 49.140 135.825 ;
        RECT 51.670 135.810 51.990 135.870 ;
        RECT 53.050 135.810 53.370 135.870 ;
        RECT 57.190 135.810 57.510 136.070 ;
        RECT 58.125 136.010 58.415 136.055 ;
        RECT 58.660 136.010 58.800 136.165 ;
        RECT 59.030 136.150 59.350 136.210 ;
        RECT 62.250 136.150 62.570 136.210 ;
        RECT 64.550 136.150 64.870 136.410 ;
        RECT 65.445 136.350 65.735 136.395 ;
        RECT 66.635 136.350 66.925 136.395 ;
        RECT 69.155 136.350 69.445 136.395 ;
        RECT 65.445 136.210 69.445 136.350 ;
        RECT 65.445 136.165 65.735 136.210 ;
        RECT 66.635 136.165 66.925 136.210 ;
        RECT 69.155 136.165 69.445 136.210 ;
        RECT 58.125 135.870 58.800 136.010 ;
        RECT 59.490 136.010 59.810 136.070 ;
        RECT 60.885 136.010 61.175 136.055 ;
        RECT 59.490 135.870 61.175 136.010 ;
        RECT 58.125 135.825 58.415 135.870 ;
        RECT 59.490 135.810 59.810 135.870 ;
        RECT 60.885 135.825 61.175 135.870 ;
        RECT 44.860 135.530 49.140 135.670 ;
        RECT 42.025 135.485 42.315 135.530 ;
        RECT 44.325 135.485 44.615 135.530 ;
        RECT 43.850 135.130 44.170 135.390 ;
        RECT 53.140 135.330 53.280 135.810 ;
        RECT 57.650 135.670 57.970 135.730 ;
        RECT 59.950 135.670 60.270 135.730 ;
        RECT 63.185 135.670 63.475 135.715 ;
        RECT 57.650 135.530 63.475 135.670 ;
        RECT 57.650 135.470 57.970 135.530 ;
        RECT 59.950 135.470 60.270 135.530 ;
        RECT 63.185 135.485 63.475 135.530 ;
        RECT 65.900 135.670 66.190 135.715 ;
        RECT 67.770 135.670 68.090 135.730 ;
        RECT 65.900 135.530 68.090 135.670 ;
        RECT 69.700 135.670 69.840 136.890 ;
        RECT 71.465 136.890 73.610 137.030 ;
        RECT 71.465 136.845 71.755 136.890 ;
        RECT 73.290 136.830 73.610 136.890 ;
        RECT 76.050 137.030 76.370 137.090 ;
        RECT 76.985 137.030 77.275 137.075 ;
        RECT 83.425 137.030 83.715 137.075 ;
        RECT 96.750 137.030 97.070 137.090 ;
        RECT 97.685 137.030 97.975 137.075 ;
        RECT 76.050 136.890 77.275 137.030 ;
        RECT 76.050 136.830 76.370 136.890 ;
        RECT 76.985 136.845 77.275 136.890 ;
        RECT 83.040 136.890 83.715 137.030 ;
        RECT 82.030 136.690 82.350 136.750 ;
        RECT 83.040 136.690 83.180 136.890 ;
        RECT 83.425 136.845 83.715 136.890 ;
        RECT 94.080 136.890 95.600 137.030 ;
        RECT 94.080 136.690 94.220 136.890 ;
        RECT 82.030 136.550 83.180 136.690 ;
        RECT 83.500 136.550 94.220 136.690 ;
        RECT 82.030 136.490 82.350 136.550 ;
        RECT 72.830 136.350 73.150 136.410 ;
        RECT 83.500 136.350 83.640 136.550 ;
        RECT 72.830 136.210 83.640 136.350 ;
        RECT 72.830 136.150 73.150 136.210 ;
        RECT 84.330 136.150 84.650 136.410 ;
        RECT 88.930 136.150 89.250 136.410 ;
        RECT 90.325 136.350 90.615 136.395 ;
        RECT 90.325 136.210 93.300 136.350 ;
        RECT 90.325 136.165 90.615 136.210 ;
        RECT 80.190 136.010 80.510 136.070 ;
        RECT 82.045 136.010 82.335 136.055 ;
        RECT 75.680 135.870 78.120 136.010 ;
        RECT 75.680 135.730 75.820 135.870 ;
        RECT 74.225 135.670 74.515 135.715 ;
        RECT 69.700 135.530 74.515 135.670 ;
        RECT 65.900 135.485 66.190 135.530 ;
        RECT 67.770 135.470 68.090 135.530 ;
        RECT 74.225 135.485 74.515 135.530 ;
        RECT 75.590 135.470 75.910 135.730 ;
        RECT 76.970 135.715 77.290 135.730 ;
        RECT 77.980 135.715 78.120 135.870 ;
        RECT 80.190 135.870 82.335 136.010 ;
        RECT 80.190 135.810 80.510 135.870 ;
        RECT 82.045 135.825 82.335 135.870 ;
        RECT 83.410 135.810 83.730 136.070 ;
        RECT 83.885 136.010 84.175 136.055 ;
        RECT 84.420 136.010 84.560 136.150 ;
        RECT 83.885 135.870 84.560 136.010 ;
        RECT 83.885 135.825 84.175 135.870 ;
        RECT 84.790 135.810 85.110 136.070 ;
        RECT 88.485 135.825 88.775 136.055 ;
        RECT 89.850 136.010 90.170 136.070 ;
        RECT 93.160 136.055 93.300 136.210 ;
        RECT 92.165 136.010 92.455 136.055 ;
        RECT 89.850 135.870 92.455 136.010 ;
        RECT 76.905 135.485 77.290 135.715 ;
        RECT 77.905 135.485 78.195 135.715 ;
        RECT 76.970 135.470 77.290 135.485 ;
        RECT 78.350 135.470 78.670 135.730 ;
        RECT 82.490 135.670 82.810 135.730 ;
        RECT 88.560 135.670 88.700 135.825 ;
        RECT 89.850 135.810 90.170 135.870 ;
        RECT 92.165 135.825 92.455 135.870 ;
        RECT 93.085 135.825 93.375 136.055 ;
        RECT 82.490 135.530 88.700 135.670 ;
        RECT 92.240 135.670 92.380 135.825 ;
        RECT 93.530 135.810 93.850 136.070 ;
        RECT 94.080 136.055 94.220 136.550 ;
        RECT 94.925 136.505 95.215 136.735 ;
        RECT 95.460 136.690 95.600 136.890 ;
        RECT 96.750 136.890 97.975 137.030 ;
        RECT 96.750 136.830 97.070 136.890 ;
        RECT 97.685 136.845 97.975 136.890 ;
        RECT 96.290 136.690 96.610 136.750 ;
        RECT 108.250 136.690 108.570 136.750 ;
        RECT 95.460 136.550 108.570 136.690 ;
        RECT 94.450 136.150 94.770 136.410 ;
        RECT 95.000 136.350 95.140 136.505 ;
        RECT 96.290 136.490 96.610 136.550 ;
        RECT 108.250 136.490 108.570 136.550 ;
        RECT 95.000 136.210 96.520 136.350 ;
        RECT 94.005 135.825 94.295 136.055 ;
        RECT 94.540 136.010 94.680 136.150 ;
        RECT 96.380 136.055 96.520 136.210 ;
        RECT 95.385 136.010 95.675 136.055 ;
        RECT 94.540 135.870 95.675 136.010 ;
        RECT 95.385 135.825 95.675 135.870 ;
        RECT 96.305 135.825 96.595 136.055 ;
        RECT 97.225 136.010 97.515 136.055 ;
        RECT 98.605 136.010 98.895 136.055 ;
        RECT 97.225 135.870 98.895 136.010 ;
        RECT 97.225 135.825 97.515 135.870 ;
        RECT 98.605 135.825 98.895 135.870 ;
        RECT 106.870 135.670 107.190 135.730 ;
        RECT 111.470 135.670 111.790 135.730 ;
        RECT 92.240 135.530 111.790 135.670 ;
        RECT 82.490 135.470 82.810 135.530 ;
        RECT 59.490 135.330 59.810 135.390 ;
        RECT 53.140 135.190 59.810 135.330 ;
        RECT 59.490 135.130 59.810 135.190 ;
        RECT 61.330 135.130 61.650 135.390 ;
        RECT 62.250 135.375 62.570 135.390 ;
        RECT 62.185 135.145 62.570 135.375 ;
        RECT 62.250 135.130 62.570 135.145 ;
        RECT 72.370 135.130 72.690 135.390 ;
        RECT 73.225 135.330 73.515 135.375 ;
        RECT 73.750 135.330 74.070 135.390 ;
        RECT 73.225 135.190 74.070 135.330 ;
        RECT 73.225 135.145 73.515 135.190 ;
        RECT 73.750 135.130 74.070 135.190 ;
        RECT 76.050 135.130 76.370 135.390 ;
        RECT 78.440 135.330 78.580 135.470 ;
        RECT 83.870 135.330 84.190 135.390 ;
        RECT 78.440 135.190 84.190 135.330 ;
        RECT 83.870 135.130 84.190 135.190 ;
        RECT 84.330 135.130 84.650 135.390 ;
        RECT 88.560 135.330 88.700 135.530 ;
        RECT 106.870 135.470 107.190 135.530 ;
        RECT 111.470 135.470 111.790 135.530 ;
        RECT 92.150 135.330 92.470 135.390 ;
        RECT 88.560 135.190 92.470 135.330 ;
        RECT 92.150 135.130 92.470 135.190 ;
        RECT 94.450 135.330 94.770 135.390 ;
        RECT 110.090 135.330 110.410 135.390 ;
        RECT 94.450 135.190 110.410 135.330 ;
        RECT 94.450 135.130 94.770 135.190 ;
        RECT 110.090 135.130 110.410 135.190 ;
        RECT 11.120 134.510 151.295 134.990 ;
        RECT 31.430 134.310 31.750 134.370 ;
        RECT 31.905 134.310 32.195 134.355 ;
        RECT 54.445 134.310 54.735 134.355 ;
        RECT 57.190 134.310 57.510 134.370 ;
        RECT 68.230 134.310 68.550 134.370 ;
        RECT 69.150 134.310 69.470 134.370 ;
        RECT 31.430 134.170 32.195 134.310 ;
        RECT 31.430 134.110 31.750 134.170 ;
        RECT 31.905 134.125 32.195 134.170 ;
        RECT 36.580 134.170 40.400 134.310 ;
        RECT 30.050 133.770 30.370 134.030 ;
        RECT 31.980 133.970 32.120 134.125 ;
        RECT 31.980 133.830 35.800 133.970 ;
        RECT 30.140 133.630 30.280 133.770 ;
        RECT 35.660 133.690 35.800 133.830 ;
        RECT 36.580 133.725 36.720 134.170 ;
        RECT 32.365 133.630 32.655 133.675 ;
        RECT 30.140 133.490 32.655 133.630 ;
        RECT 32.365 133.445 32.655 133.490 ;
        RECT 35.570 133.430 35.890 133.690 ;
        RECT 36.505 133.495 36.795 133.725 ;
        RECT 36.950 133.620 37.270 133.690 ;
        RECT 38.805 133.630 39.095 133.675 ;
        RECT 37.500 133.620 39.095 133.630 ;
        RECT 36.950 133.490 39.095 133.620 ;
        RECT 36.950 133.480 37.640 133.490 ;
        RECT 36.950 133.430 37.270 133.480 ;
        RECT 38.805 133.445 39.095 133.490 ;
        RECT 39.250 133.430 39.570 133.690 ;
        RECT 39.725 133.445 40.015 133.675 ;
        RECT 36.045 132.950 36.335 132.995 ;
        RECT 39.800 132.950 39.940 133.445 ;
        RECT 36.045 132.810 39.940 132.950 ;
        RECT 40.260 132.950 40.400 134.170 ;
        RECT 40.720 134.170 54.200 134.310 ;
        RECT 40.720 133.675 40.860 134.170 ;
        RECT 43.850 133.970 44.170 134.030 ;
        RECT 42.560 133.830 46.380 133.970 ;
        RECT 42.560 133.675 42.700 133.830 ;
        RECT 43.850 133.770 44.170 133.830 ;
        RECT 46.240 133.675 46.380 133.830 ;
        RECT 46.610 133.770 46.930 134.030 ;
        RECT 51.670 133.970 51.990 134.030 ;
        RECT 47.160 133.830 51.990 133.970 ;
        RECT 54.060 133.970 54.200 134.170 ;
        RECT 54.445 134.170 57.510 134.310 ;
        RECT 54.445 134.125 54.735 134.170 ;
        RECT 57.190 134.110 57.510 134.170 ;
        RECT 65.100 134.170 68.000 134.310 ;
        RECT 65.100 133.970 65.240 134.170 ;
        RECT 67.860 133.970 68.000 134.170 ;
        RECT 68.230 134.170 69.470 134.310 ;
        RECT 68.230 134.110 68.550 134.170 ;
        RECT 69.150 134.110 69.470 134.170 ;
        RECT 73.750 134.310 74.070 134.370 ;
        RECT 104.125 134.310 104.415 134.355 ;
        RECT 73.750 134.170 89.160 134.310 ;
        RECT 73.750 134.110 74.070 134.170 ;
        RECT 89.020 134.030 89.160 134.170 ;
        RECT 104.125 134.170 107.560 134.310 ;
        RECT 104.125 134.125 104.415 134.170 ;
        RECT 75.130 133.970 75.450 134.030 ;
        RECT 54.060 133.830 65.240 133.970 ;
        RECT 65.560 133.830 67.080 133.970 ;
        RECT 40.645 133.445 40.935 133.675 ;
        RECT 41.565 133.445 41.855 133.675 ;
        RECT 42.485 133.445 42.775 133.675 ;
        RECT 44.785 133.445 45.075 133.675 ;
        RECT 46.165 133.445 46.455 133.675 ;
        RECT 41.640 133.290 41.780 133.445 ;
        RECT 42.945 133.290 43.235 133.335 ;
        RECT 41.640 133.150 44.080 133.290 ;
        RECT 42.945 133.105 43.235 133.150 ;
        RECT 43.940 132.950 44.080 133.150 ;
        RECT 44.310 133.090 44.630 133.350 ;
        RECT 44.860 133.290 45.000 133.445 ;
        RECT 47.160 133.290 47.300 133.830 ;
        RECT 51.670 133.770 51.990 133.830 ;
        RECT 47.545 133.445 47.835 133.675 ;
        RECT 52.145 133.630 52.435 133.675 ;
        RECT 60.870 133.630 61.190 133.690 ;
        RECT 65.560 133.675 65.700 133.830 ;
        RECT 52.145 133.490 61.190 133.630 ;
        RECT 52.145 133.445 52.435 133.490 ;
        RECT 44.860 133.150 47.300 133.290 ;
        RECT 46.610 132.950 46.930 133.010 ;
        RECT 40.260 132.810 43.620 132.950 ;
        RECT 43.940 132.810 46.930 132.950 ;
        RECT 36.045 132.765 36.335 132.810 ;
        RECT 37.410 132.410 37.730 132.670 ;
        RECT 42.470 132.410 42.790 132.670 ;
        RECT 43.480 132.610 43.620 132.810 ;
        RECT 46.610 132.750 46.930 132.810 ;
        RECT 47.620 132.950 47.760 133.445 ;
        RECT 60.870 133.430 61.190 133.490 ;
        RECT 65.485 133.445 65.775 133.675 ;
        RECT 66.405 133.445 66.695 133.675 ;
        RECT 57.650 132.950 57.970 133.010 ;
        RECT 47.620 132.810 57.970 132.950 ;
        RECT 66.480 132.950 66.620 133.445 ;
        RECT 66.940 133.290 67.080 133.830 ;
        RECT 67.860 133.830 75.450 133.970 ;
        RECT 67.860 133.630 68.000 133.830 ;
        RECT 75.130 133.770 75.450 133.830 ;
        RECT 88.930 133.770 89.250 134.030 ;
        RECT 107.420 134.015 107.560 134.170 ;
        RECT 105.045 133.970 105.335 134.015 ;
        RECT 102.360 133.830 105.335 133.970 ;
        RECT 68.705 133.630 68.995 133.675 ;
        RECT 67.860 133.490 68.995 133.630 ;
        RECT 68.705 133.445 68.995 133.490 ;
        RECT 70.085 133.630 70.375 133.675 ;
        RECT 72.370 133.630 72.690 133.690 ;
        RECT 70.085 133.490 72.690 133.630 ;
        RECT 70.085 133.445 70.375 133.490 ;
        RECT 72.370 133.430 72.690 133.490 ;
        RECT 101.350 133.630 101.670 133.690 ;
        RECT 102.360 133.675 102.500 133.830 ;
        RECT 105.045 133.785 105.335 133.830 ;
        RECT 107.345 133.785 107.635 134.015 ;
        RECT 102.285 133.630 102.575 133.675 ;
        RECT 101.350 133.490 102.575 133.630 ;
        RECT 101.350 133.430 101.670 133.490 ;
        RECT 102.285 133.445 102.575 133.490 ;
        RECT 104.110 133.430 104.430 133.690 ;
        RECT 104.570 133.430 104.890 133.690 ;
        RECT 106.425 133.630 106.715 133.675 ;
        RECT 106.870 133.630 107.190 133.690 ;
        RECT 106.425 133.490 107.190 133.630 ;
        RECT 106.425 133.445 106.715 133.490 ;
        RECT 106.870 133.430 107.190 133.490 ;
        RECT 107.805 133.445 108.095 133.675 ;
        RECT 67.770 133.290 68.090 133.350 ;
        RECT 66.940 133.150 68.090 133.290 ;
        RECT 67.770 133.090 68.090 133.150 ;
        RECT 69.625 133.290 69.915 133.335 ;
        RECT 76.050 133.290 76.370 133.350 ;
        RECT 69.625 133.150 76.370 133.290 ;
        RECT 69.625 133.105 69.915 133.150 ;
        RECT 76.050 133.090 76.370 133.150 ;
        RECT 102.745 133.105 103.035 133.335 ;
        RECT 104.200 133.290 104.340 133.430 ;
        RECT 107.880 133.290 108.020 133.445 ;
        RECT 108.250 133.430 108.570 133.690 ;
        RECT 110.090 133.430 110.410 133.690 ;
        RECT 110.565 133.445 110.855 133.675 ;
        RECT 111.485 133.630 111.775 133.675 ;
        RECT 111.945 133.630 112.235 133.675 ;
        RECT 111.485 133.490 112.235 133.630 ;
        RECT 111.485 133.445 111.775 133.490 ;
        RECT 111.945 133.445 112.235 133.490 ;
        RECT 110.640 133.290 110.780 133.445 ;
        RECT 104.200 133.150 108.020 133.290 ;
        RECT 109.260 133.150 110.780 133.290 ;
        RECT 73.750 132.950 74.070 133.010 ;
        RECT 66.480 132.810 74.070 132.950 ;
        RECT 47.620 132.610 47.760 132.810 ;
        RECT 57.650 132.750 57.970 132.810 ;
        RECT 73.750 132.750 74.070 132.810 ;
        RECT 74.670 132.950 74.990 133.010 ;
        RECT 102.820 132.950 102.960 133.105 ;
        RECT 106.410 132.950 106.730 133.010 ;
        RECT 109.260 132.995 109.400 133.150 ;
        RECT 74.670 132.810 90.540 132.950 ;
        RECT 102.820 132.810 106.730 132.950 ;
        RECT 74.670 132.750 74.990 132.810 ;
        RECT 90.400 132.670 90.540 132.810 ;
        RECT 106.410 132.750 106.730 132.810 ;
        RECT 109.185 132.765 109.475 132.995 ;
        RECT 43.480 132.470 47.760 132.610 ;
        RECT 48.450 132.410 48.770 132.670 ;
        RECT 53.050 132.410 53.370 132.670 ;
        RECT 56.270 132.610 56.590 132.670 ;
        RECT 65.930 132.610 66.250 132.670 ;
        RECT 56.270 132.470 66.250 132.610 ;
        RECT 56.270 132.410 56.590 132.470 ;
        RECT 65.930 132.410 66.250 132.470 ;
        RECT 67.785 132.610 68.075 132.655 ;
        RECT 69.150 132.610 69.470 132.670 ;
        RECT 67.785 132.470 69.470 132.610 ;
        RECT 67.785 132.425 68.075 132.470 ;
        RECT 69.150 132.410 69.470 132.470 ;
        RECT 76.970 132.610 77.290 132.670 ;
        RECT 82.950 132.610 83.270 132.670 ;
        RECT 76.970 132.470 83.270 132.610 ;
        RECT 76.970 132.410 77.290 132.470 ;
        RECT 82.950 132.410 83.270 132.470 ;
        RECT 90.310 132.410 90.630 132.670 ;
        RECT 112.850 132.410 113.170 132.670 ;
        RECT 11.120 131.790 150.500 132.270 ;
        RECT 27.290 131.390 27.610 131.650 ;
        RECT 37.410 131.390 37.730 131.650 ;
        RECT 42.470 131.390 42.790 131.650 ;
        RECT 48.450 131.590 48.770 131.650 ;
        RECT 43.480 131.450 48.770 131.590 ;
        RECT 30.050 131.250 30.340 131.295 ;
        RECT 31.620 131.250 31.910 131.295 ;
        RECT 33.720 131.250 34.010 131.295 ;
        RECT 30.050 131.110 34.010 131.250 ;
        RECT 30.050 131.065 30.340 131.110 ;
        RECT 31.620 131.065 31.910 131.110 ;
        RECT 33.720 131.065 34.010 131.110 ;
        RECT 29.615 130.910 29.905 130.955 ;
        RECT 32.135 130.910 32.425 130.955 ;
        RECT 33.325 130.910 33.615 130.955 ;
        RECT 37.500 130.910 37.640 131.390 ;
        RECT 29.615 130.770 33.615 130.910 ;
        RECT 29.615 130.725 29.905 130.770 ;
        RECT 32.135 130.725 32.425 130.770 ;
        RECT 33.325 130.725 33.615 130.770 ;
        RECT 33.820 130.770 37.640 130.910 ;
        RECT 32.925 130.570 33.215 130.615 ;
        RECT 33.820 130.570 33.960 130.770 ;
        RECT 32.925 130.430 33.960 130.570 ;
        RECT 34.205 130.570 34.495 130.615 ;
        RECT 37.870 130.570 38.190 130.630 ;
        RECT 41.550 130.570 41.870 130.630 ;
        RECT 34.205 130.430 41.870 130.570 ;
        RECT 42.560 130.570 42.700 131.390 ;
        RECT 43.480 130.615 43.620 131.450 ;
        RECT 48.450 131.390 48.770 131.450 ;
        RECT 52.605 131.590 52.895 131.635 ;
        RECT 54.890 131.590 55.210 131.650 ;
        RECT 52.605 131.450 55.210 131.590 ;
        RECT 52.605 131.405 52.895 131.450 ;
        RECT 54.890 131.390 55.210 131.450 ;
        RECT 56.730 131.390 57.050 131.650 ;
        RECT 60.425 131.590 60.715 131.635 ;
        RECT 61.330 131.590 61.650 131.650 ;
        RECT 60.425 131.450 61.650 131.590 ;
        RECT 60.425 131.405 60.715 131.450 ;
        RECT 61.330 131.390 61.650 131.450 ;
        RECT 65.930 131.590 66.250 131.650 ;
        RECT 82.950 131.590 83.270 131.650 ;
        RECT 99.050 131.590 99.370 131.650 ;
        RECT 65.930 131.450 78.120 131.590 ;
        RECT 65.930 131.390 66.250 131.450 ;
        RECT 44.325 131.250 44.615 131.295 ;
        RECT 56.270 131.250 56.590 131.310 ;
        RECT 44.325 131.110 56.590 131.250 ;
        RECT 44.325 131.065 44.615 131.110 ;
        RECT 56.270 131.050 56.590 131.110 ;
        RECT 55.350 130.910 55.670 130.970 ;
        RECT 52.680 130.770 55.670 130.910 ;
        RECT 42.945 130.570 43.235 130.615 ;
        RECT 42.560 130.430 43.235 130.570 ;
        RECT 32.925 130.385 33.215 130.430 ;
        RECT 34.205 130.385 34.495 130.430 ;
        RECT 37.870 130.370 38.190 130.430 ;
        RECT 41.550 130.370 41.870 130.430 ;
        RECT 42.945 130.385 43.235 130.430 ;
        RECT 43.405 130.385 43.695 130.615 ;
        RECT 44.785 130.570 45.075 130.615 ;
        RECT 48.910 130.570 49.230 130.630 ;
        RECT 52.680 130.615 52.820 130.770 ;
        RECT 55.350 130.710 55.670 130.770 ;
        RECT 55.825 130.910 56.115 130.955 ;
        RECT 56.820 130.910 56.960 131.390 ;
        RECT 57.650 131.250 57.970 131.310 ;
        RECT 73.765 131.250 74.055 131.295 ;
        RECT 57.650 131.110 60.180 131.250 ;
        RECT 57.650 131.050 57.970 131.110 ;
        RECT 60.040 130.955 60.180 131.110 ;
        RECT 73.765 131.110 76.905 131.250 ;
        RECT 73.765 131.065 74.055 131.110 ;
        RECT 59.965 130.910 60.255 130.955 ;
        RECT 75.590 130.910 75.910 130.970 ;
        RECT 55.825 130.770 58.800 130.910 ;
        RECT 55.825 130.725 56.115 130.770 ;
        RECT 44.785 130.430 49.230 130.570 ;
        RECT 44.785 130.385 45.075 130.430 ;
        RECT 44.310 130.230 44.630 130.290 ;
        RECT 44.860 130.230 45.000 130.385 ;
        RECT 48.910 130.370 49.230 130.430 ;
        RECT 52.605 130.385 52.895 130.615 ;
        RECT 53.985 130.570 54.275 130.615 ;
        RECT 55.900 130.570 56.040 130.725 ;
        RECT 53.985 130.430 56.040 130.570 ;
        RECT 53.985 130.385 54.275 130.430 ;
        RECT 56.285 130.385 56.575 130.615 ;
        RECT 56.745 130.570 57.035 130.615 ;
        RECT 57.650 130.570 57.970 130.630 ;
        RECT 58.660 130.615 58.800 130.770 ;
        RECT 59.965 130.770 68.920 130.910 ;
        RECT 59.965 130.725 60.255 130.770 ;
        RECT 56.745 130.430 57.970 130.570 ;
        RECT 56.745 130.385 57.035 130.430 ;
        RECT 43.480 130.090 45.000 130.230 ;
        RECT 53.525 130.230 53.815 130.275 ;
        RECT 56.360 130.230 56.500 130.385 ;
        RECT 57.650 130.370 57.970 130.430 ;
        RECT 58.585 130.385 58.875 130.615 ;
        RECT 57.190 130.230 57.510 130.290 ;
        RECT 68.245 130.230 68.535 130.275 ;
        RECT 53.525 130.090 57.510 130.230 ;
        RECT 43.480 129.950 43.620 130.090 ;
        RECT 44.310 130.030 44.630 130.090 ;
        RECT 53.525 130.045 53.815 130.090 ;
        RECT 57.190 130.030 57.510 130.090 ;
        RECT 59.120 130.090 68.535 130.230 ;
        RECT 68.780 130.230 68.920 130.770 ;
        RECT 70.390 130.770 75.910 130.910 ;
        RECT 69.165 130.570 69.455 130.615 ;
        RECT 70.390 130.570 70.530 130.770 ;
        RECT 75.590 130.710 75.910 130.770 ;
        RECT 69.165 130.430 70.530 130.570 ;
        RECT 69.165 130.385 69.455 130.430 ;
        RECT 74.685 130.385 74.975 130.615 ;
        RECT 73.750 130.230 74.070 130.290 ;
        RECT 68.780 130.090 74.070 130.230 ;
        RECT 74.760 130.230 74.900 130.385 ;
        RECT 75.130 130.370 75.450 130.630 ;
        RECT 76.765 130.615 76.905 131.110 ;
        RECT 77.980 130.910 78.120 131.450 ;
        RECT 82.950 131.450 88.240 131.590 ;
        RECT 82.950 131.390 83.270 131.450 ;
        RECT 78.810 131.050 79.130 131.310 ;
        RECT 79.285 130.910 79.575 130.955 ;
        RECT 77.980 130.770 79.575 130.910 ;
        RECT 79.285 130.725 79.575 130.770 ;
        RECT 76.690 130.385 76.980 130.615 ;
        RECT 80.665 130.570 80.955 130.615 ;
        RECT 82.030 130.570 82.350 130.630 ;
        RECT 78.900 130.430 82.350 130.570 ;
        RECT 83.040 130.570 83.180 131.390 ;
        RECT 83.425 131.250 83.715 131.295 ;
        RECT 84.330 131.250 84.650 131.310 ;
        RECT 83.425 131.110 84.650 131.250 ;
        RECT 88.100 131.250 88.240 131.450 ;
        RECT 99.050 131.450 114.460 131.590 ;
        RECT 99.050 131.390 99.370 131.450 ;
        RECT 100.445 131.250 100.735 131.295 ;
        RECT 104.570 131.250 104.890 131.310 ;
        RECT 88.100 131.110 88.700 131.250 ;
        RECT 83.425 131.065 83.715 131.110 ;
        RECT 84.330 131.050 84.650 131.110 ;
        RECT 84.420 130.910 84.560 131.050 ;
        RECT 84.420 130.770 88.240 130.910 ;
        RECT 84.345 130.570 84.635 130.615 ;
        RECT 83.040 130.430 84.635 130.570 ;
        RECT 78.900 130.230 79.040 130.430 ;
        RECT 80.665 130.385 80.955 130.430 ;
        RECT 82.030 130.370 82.350 130.430 ;
        RECT 84.345 130.385 84.635 130.430 ;
        RECT 85.250 130.570 85.570 130.630 ;
        RECT 88.100 130.615 88.240 130.770 ;
        RECT 88.560 130.615 88.700 131.110 ;
        RECT 100.445 131.110 104.890 131.250 ;
        RECT 100.445 131.065 100.735 131.110 ;
        RECT 104.570 131.050 104.890 131.110 ;
        RECT 107.345 131.065 107.635 131.295 ;
        RECT 110.090 131.250 110.380 131.295 ;
        RECT 111.660 131.250 111.950 131.295 ;
        RECT 113.760 131.250 114.050 131.295 ;
        RECT 110.090 131.110 114.050 131.250 ;
        RECT 110.090 131.065 110.380 131.110 ;
        RECT 111.660 131.065 111.950 131.110 ;
        RECT 113.760 131.065 114.050 131.110 ;
        RECT 99.065 130.910 99.355 130.955 ;
        RECT 104.110 130.910 104.430 130.970 ;
        RECT 107.420 130.910 107.560 131.065 ;
        RECT 114.320 130.955 114.460 131.450 ;
        RECT 118.370 131.390 118.690 131.650 ;
        RECT 99.065 130.770 107.560 130.910 ;
        RECT 109.655 130.910 109.945 130.955 ;
        RECT 112.175 130.910 112.465 130.955 ;
        RECT 113.365 130.910 113.655 130.955 ;
        RECT 109.655 130.770 113.655 130.910 ;
        RECT 99.065 130.725 99.355 130.770 ;
        RECT 104.110 130.710 104.430 130.770 ;
        RECT 109.655 130.725 109.945 130.770 ;
        RECT 112.175 130.725 112.465 130.770 ;
        RECT 113.365 130.725 113.655 130.770 ;
        RECT 114.245 130.910 114.535 130.955 ;
        RECT 118.460 130.910 118.600 131.390 ;
        RECT 114.245 130.770 118.600 130.910 ;
        RECT 114.245 130.725 114.535 130.770 ;
        RECT 86.645 130.570 86.935 130.615 ;
        RECT 85.250 130.430 86.935 130.570 ;
        RECT 85.250 130.370 85.570 130.430 ;
        RECT 86.645 130.385 86.935 130.430 ;
        RECT 88.025 130.385 88.315 130.615 ;
        RECT 88.485 130.385 88.775 130.615 ;
        RECT 98.605 130.570 98.895 130.615 ;
        RECT 102.270 130.570 102.590 130.630 ;
        RECT 98.605 130.430 102.590 130.570 ;
        RECT 98.605 130.385 98.895 130.430 ;
        RECT 102.270 130.370 102.590 130.430 ;
        RECT 112.850 130.615 113.170 130.630 ;
        RECT 112.850 130.570 113.200 130.615 ;
        RECT 112.850 130.430 113.365 130.570 ;
        RECT 112.850 130.385 113.200 130.430 ;
        RECT 112.850 130.370 113.170 130.385 ;
        RECT 74.760 130.090 79.040 130.230 ;
        RECT 79.270 130.230 79.590 130.290 ;
        RECT 79.745 130.230 80.035 130.275 ;
        RECT 79.270 130.090 80.035 130.230 ;
        RECT 59.120 129.950 59.260 130.090 ;
        RECT 68.245 130.045 68.535 130.090 ;
        RECT 42.010 129.690 42.330 129.950 ;
        RECT 43.390 129.690 43.710 129.950 ;
        RECT 54.430 129.690 54.750 129.950 ;
        RECT 59.030 129.690 59.350 129.950 ;
        RECT 60.410 129.890 60.730 129.950 ;
        RECT 61.345 129.890 61.635 129.935 ;
        RECT 60.410 129.750 61.635 129.890 ;
        RECT 60.410 129.690 60.730 129.750 ;
        RECT 61.345 129.705 61.635 129.750 ;
        RECT 66.390 129.890 66.710 129.950 ;
        RECT 67.325 129.890 67.615 129.935 ;
        RECT 66.390 129.750 67.615 129.890 ;
        RECT 68.320 129.890 68.460 130.045 ;
        RECT 73.750 130.030 74.070 130.090 ;
        RECT 79.270 130.030 79.590 130.090 ;
        RECT 79.745 130.045 80.035 130.090 ;
        RECT 84.790 130.230 85.110 130.290 ;
        RECT 87.565 130.230 87.855 130.275 ;
        RECT 84.790 130.090 87.855 130.230 ;
        RECT 84.790 130.030 85.110 130.090 ;
        RECT 87.565 130.045 87.855 130.090 ;
        RECT 74.670 129.890 74.990 129.950 ;
        RECT 68.320 129.750 74.990 129.890 ;
        RECT 66.390 129.690 66.710 129.750 ;
        RECT 67.325 129.705 67.615 129.750 ;
        RECT 74.670 129.690 74.990 129.750 ;
        RECT 76.050 129.690 76.370 129.950 ;
        RECT 76.985 129.890 77.275 129.935 ;
        RECT 81.585 129.890 81.875 129.935 ;
        RECT 76.985 129.750 81.875 129.890 ;
        RECT 76.985 129.705 77.275 129.750 ;
        RECT 81.585 129.705 81.875 129.750 ;
        RECT 85.250 129.690 85.570 129.950 ;
        RECT 86.170 129.690 86.490 129.950 ;
        RECT 89.390 129.690 89.710 129.950 ;
        RECT 11.120 129.070 151.295 129.550 ;
        RECT 39.250 128.870 39.570 128.930 ;
        RECT 51.685 128.870 51.975 128.915 ;
        RECT 53.050 128.870 53.370 128.930 ;
        RECT 54.430 128.870 54.750 128.930 ;
        RECT 59.965 128.870 60.255 128.915 ;
        RECT 61.345 128.870 61.635 128.915 ;
        RECT 39.250 128.730 53.370 128.870 ;
        RECT 39.250 128.670 39.570 128.730 ;
        RECT 51.685 128.685 51.975 128.730 ;
        RECT 53.050 128.670 53.370 128.730 ;
        RECT 53.600 128.730 54.750 128.870 ;
        RECT 53.600 128.530 53.740 128.730 ;
        RECT 54.430 128.670 54.750 128.730 ;
        RECT 56.590 128.730 59.720 128.870 ;
        RECT 53.140 128.390 53.740 128.530 ;
        RECT 53.970 128.530 54.290 128.590 ;
        RECT 56.590 128.530 56.730 128.730 ;
        RECT 53.970 128.390 56.730 128.530 ;
        RECT 42.010 127.990 42.330 128.250 ;
        RECT 42.945 128.005 43.235 128.235 ;
        RECT 43.865 128.190 44.155 128.235 ;
        RECT 44.325 128.190 44.615 128.235 ;
        RECT 43.865 128.050 44.615 128.190 ;
        RECT 43.865 128.005 44.155 128.050 ;
        RECT 44.325 128.005 44.615 128.050 ;
        RECT 48.925 128.005 49.215 128.235 ;
        RECT 49.845 128.190 50.135 128.235 ;
        RECT 51.670 128.190 51.960 128.235 ;
        RECT 52.130 128.190 52.450 128.250 ;
        RECT 49.845 128.050 50.980 128.190 ;
        RECT 49.845 128.005 50.135 128.050 ;
        RECT 43.020 127.850 43.160 128.005 ;
        RECT 49.000 127.850 49.140 128.005 ;
        RECT 43.020 127.710 49.140 127.850 ;
        RECT 45.230 126.970 45.550 127.230 ;
        RECT 49.000 127.170 49.140 127.710 ;
        RECT 49.370 127.650 49.690 127.910 ;
        RECT 50.840 127.555 50.980 128.050 ;
        RECT 51.670 128.050 52.820 128.190 ;
        RECT 51.670 128.005 51.960 128.050 ;
        RECT 52.130 127.990 52.450 128.050 ;
        RECT 50.765 127.325 51.055 127.555 ;
        RECT 52.680 127.510 52.820 128.050 ;
        RECT 53.140 127.850 53.280 128.390 ;
        RECT 53.970 128.330 54.290 128.390 ;
        RECT 59.030 128.330 59.350 128.590 ;
        RECT 59.580 128.530 59.720 128.730 ;
        RECT 59.965 128.730 61.635 128.870 ;
        RECT 59.965 128.685 60.255 128.730 ;
        RECT 61.345 128.685 61.635 128.730 ;
        RECT 66.850 128.670 67.170 128.930 ;
        RECT 73.765 128.685 74.055 128.915 ;
        RECT 75.130 128.870 75.450 128.930 ;
        RECT 75.605 128.870 75.895 128.915 ;
        RECT 79.270 128.870 79.590 128.930 ;
        RECT 82.490 128.870 82.810 128.930 ;
        RECT 75.130 128.730 79.590 128.870 ;
        RECT 66.940 128.530 67.080 128.670 ;
        RECT 59.580 128.390 67.080 128.530 ;
        RECT 73.840 128.530 73.980 128.685 ;
        RECT 75.130 128.670 75.450 128.730 ;
        RECT 75.605 128.685 75.895 128.730 ;
        RECT 79.270 128.670 79.590 128.730 ;
        RECT 81.200 128.730 82.810 128.870 ;
        RECT 78.810 128.530 79.130 128.590 ;
        RECT 73.840 128.390 79.130 128.530 ;
        RECT 59.120 128.190 59.260 128.330 ;
        RECT 56.590 128.050 59.260 128.190 ;
        RECT 53.525 127.850 53.815 127.895 ;
        RECT 53.140 127.710 53.815 127.850 ;
        RECT 53.525 127.665 53.815 127.710 ;
        RECT 53.985 127.850 54.275 127.895 ;
        RECT 54.890 127.850 55.210 127.910 ;
        RECT 53.985 127.710 55.210 127.850 ;
        RECT 53.985 127.665 54.275 127.710 ;
        RECT 54.890 127.650 55.210 127.710 ;
        RECT 54.430 127.510 54.750 127.570 ;
        RECT 52.680 127.370 54.750 127.510 ;
        RECT 54.430 127.310 54.750 127.370 ;
        RECT 56.590 127.170 56.730 128.050 ;
        RECT 60.410 127.990 60.730 128.250 ;
        RECT 60.960 128.235 61.100 128.390 ;
        RECT 60.885 128.005 61.175 128.235 ;
        RECT 61.805 128.190 62.095 128.235 ;
        RECT 63.185 128.190 63.475 128.235 ;
        RECT 66.865 128.190 67.155 128.235 ;
        RECT 61.805 128.050 63.475 128.190 ;
        RECT 61.805 128.005 62.095 128.050 ;
        RECT 63.185 128.005 63.475 128.050 ;
        RECT 64.640 128.050 67.155 128.190 ;
        RECT 64.640 127.910 64.780 128.050 ;
        RECT 66.865 128.005 67.155 128.050 ;
        RECT 67.310 128.190 67.630 128.250 ;
        RECT 68.145 128.190 68.435 128.235 ;
        RECT 67.310 128.050 68.435 128.190 ;
        RECT 67.310 127.990 67.630 128.050 ;
        RECT 68.145 128.005 68.435 128.050 ;
        RECT 64.550 127.650 64.870 127.910 ;
        RECT 77.060 127.895 77.200 128.390 ;
        RECT 78.810 128.330 79.130 128.390 ;
        RECT 81.200 128.235 81.340 128.730 ;
        RECT 82.490 128.670 82.810 128.730 ;
        RECT 84.345 128.870 84.635 128.915 ;
        RECT 84.790 128.870 85.110 128.930 ;
        RECT 84.345 128.730 85.110 128.870 ;
        RECT 84.345 128.685 84.635 128.730 ;
        RECT 84.790 128.670 85.110 128.730 ;
        RECT 86.170 128.670 86.490 128.930 ;
        RECT 89.390 128.670 89.710 128.930 ;
        RECT 81.585 128.530 81.875 128.575 ;
        RECT 85.250 128.530 85.570 128.590 ;
        RECT 81.585 128.390 85.570 128.530 ;
        RECT 81.585 128.345 81.875 128.390 ;
        RECT 85.250 128.330 85.570 128.390 ;
        RECT 77.445 128.005 77.735 128.235 ;
        RECT 81.125 128.005 81.415 128.235 ;
        RECT 82.045 128.005 82.335 128.235 ;
        RECT 65.945 127.665 66.235 127.895 ;
        RECT 67.745 127.850 68.035 127.895 ;
        RECT 68.935 127.850 69.225 127.895 ;
        RECT 71.455 127.850 71.745 127.895 ;
        RECT 67.745 127.710 71.745 127.850 ;
        RECT 67.745 127.665 68.035 127.710 ;
        RECT 68.935 127.665 69.225 127.710 ;
        RECT 71.455 127.665 71.745 127.710 ;
        RECT 76.985 127.665 77.275 127.895 ;
        RECT 77.520 127.850 77.660 128.005 ;
        RECT 82.120 127.850 82.260 128.005 ;
        RECT 82.490 127.990 82.810 128.250 ;
        RECT 83.410 127.990 83.730 128.250 ;
        RECT 86.260 128.235 86.400 128.670 ;
        RECT 89.480 128.530 89.620 128.670 ;
        RECT 88.100 128.390 89.620 128.530 ;
        RECT 88.100 128.235 88.240 128.390 ;
        RECT 90.310 128.330 90.630 128.590 ;
        RECT 86.185 128.005 86.475 128.235 ;
        RECT 88.025 128.005 88.315 128.235 ;
        RECT 88.945 128.005 89.235 128.235 ;
        RECT 89.405 128.005 89.695 128.235 ;
        RECT 96.810 128.190 97.100 128.235 ;
        RECT 93.160 128.050 97.100 128.190 ;
        RECT 83.500 127.850 83.640 127.990 ;
        RECT 89.020 127.850 89.160 128.005 ;
        RECT 77.520 127.710 83.640 127.850 ;
        RECT 85.340 127.710 89.160 127.850 ;
        RECT 89.480 127.850 89.620 128.005 ;
        RECT 92.610 127.850 92.930 127.910 ;
        RECT 89.480 127.710 92.930 127.850 ;
        RECT 60.870 127.510 61.190 127.570 ;
        RECT 65.010 127.510 65.330 127.570 ;
        RECT 66.020 127.510 66.160 127.665 ;
        RECT 60.870 127.370 66.160 127.510 ;
        RECT 67.350 127.510 67.640 127.555 ;
        RECT 69.450 127.510 69.740 127.555 ;
        RECT 71.020 127.510 71.310 127.555 ;
        RECT 67.350 127.370 71.310 127.510 ;
        RECT 60.870 127.310 61.190 127.370 ;
        RECT 65.010 127.310 65.330 127.370 ;
        RECT 67.350 127.325 67.640 127.370 ;
        RECT 69.450 127.325 69.740 127.370 ;
        RECT 71.020 127.325 71.310 127.370 ;
        RECT 82.490 127.510 82.810 127.570 ;
        RECT 85.340 127.555 85.480 127.710 ;
        RECT 92.610 127.650 92.930 127.710 ;
        RECT 82.490 127.370 85.020 127.510 ;
        RECT 82.490 127.310 82.810 127.370 ;
        RECT 49.000 127.030 56.730 127.170 ;
        RECT 59.030 126.970 59.350 127.230 ;
        RECT 84.880 127.170 85.020 127.370 ;
        RECT 85.265 127.325 85.555 127.555 ;
        RECT 90.325 127.510 90.615 127.555 ;
        RECT 93.160 127.510 93.300 128.050 ;
        RECT 96.810 128.005 97.100 128.050 ;
        RECT 98.145 128.190 98.435 128.235 ;
        RECT 99.050 128.190 99.370 128.250 ;
        RECT 98.145 128.050 99.370 128.190 ;
        RECT 98.145 128.005 98.435 128.050 ;
        RECT 99.050 127.990 99.370 128.050 ;
        RECT 93.555 127.850 93.845 127.895 ;
        RECT 96.075 127.850 96.365 127.895 ;
        RECT 97.265 127.850 97.555 127.895 ;
        RECT 93.555 127.710 97.555 127.850 ;
        RECT 93.555 127.665 93.845 127.710 ;
        RECT 96.075 127.665 96.365 127.710 ;
        RECT 97.265 127.665 97.555 127.710 ;
        RECT 85.800 127.370 90.080 127.510 ;
        RECT 85.800 127.170 85.940 127.370 ;
        RECT 84.880 127.030 85.940 127.170 ;
        RECT 87.565 127.170 87.855 127.215 ;
        RECT 88.930 127.170 89.250 127.230 ;
        RECT 87.565 127.030 89.250 127.170 ;
        RECT 89.940 127.170 90.080 127.370 ;
        RECT 90.325 127.370 93.300 127.510 ;
        RECT 93.990 127.510 94.280 127.555 ;
        RECT 95.560 127.510 95.850 127.555 ;
        RECT 97.660 127.510 97.950 127.555 ;
        RECT 93.990 127.370 97.950 127.510 ;
        RECT 90.325 127.325 90.615 127.370 ;
        RECT 93.990 127.325 94.280 127.370 ;
        RECT 95.560 127.325 95.850 127.370 ;
        RECT 97.660 127.325 97.950 127.370 ;
        RECT 91.230 127.170 91.550 127.230 ;
        RECT 89.940 127.030 91.550 127.170 ;
        RECT 87.565 126.985 87.855 127.030 ;
        RECT 88.930 126.970 89.250 127.030 ;
        RECT 91.230 126.970 91.550 127.030 ;
        RECT 11.120 126.350 150.500 126.830 ;
        RECT 39.725 126.150 40.015 126.195 ;
        RECT 43.390 126.150 43.710 126.210 ;
        RECT 39.725 126.010 43.710 126.150 ;
        RECT 39.725 125.965 40.015 126.010 ;
        RECT 43.390 125.950 43.710 126.010 ;
        RECT 64.565 126.150 64.855 126.195 ;
        RECT 65.010 126.150 65.330 126.210 ;
        RECT 64.565 126.010 65.330 126.150 ;
        RECT 64.565 125.965 64.855 126.010 ;
        RECT 65.010 125.950 65.330 126.010 ;
        RECT 66.405 126.150 66.695 126.195 ;
        RECT 67.310 126.150 67.630 126.210 ;
        RECT 66.405 126.010 67.630 126.150 ;
        RECT 66.405 125.965 66.695 126.010 ;
        RECT 67.310 125.950 67.630 126.010 ;
        RECT 92.610 126.150 92.930 126.210 ;
        RECT 95.845 126.150 96.135 126.195 ;
        RECT 92.610 126.010 96.135 126.150 ;
        RECT 92.610 125.950 92.930 126.010 ;
        RECT 95.845 125.965 96.135 126.010 ;
        RECT 42.470 125.810 42.760 125.855 ;
        RECT 44.040 125.810 44.330 125.855 ;
        RECT 46.140 125.810 46.430 125.855 ;
        RECT 42.470 125.670 46.430 125.810 ;
        RECT 42.470 125.625 42.760 125.670 ;
        RECT 44.040 125.625 44.330 125.670 ;
        RECT 46.140 125.625 46.430 125.670 ;
        RECT 58.150 125.810 58.440 125.855 ;
        RECT 60.250 125.810 60.540 125.855 ;
        RECT 61.820 125.810 62.110 125.855 ;
        RECT 58.150 125.670 62.110 125.810 ;
        RECT 58.150 125.625 58.440 125.670 ;
        RECT 60.250 125.625 60.540 125.670 ;
        RECT 61.820 125.625 62.110 125.670 ;
        RECT 42.035 125.470 42.325 125.515 ;
        RECT 44.555 125.470 44.845 125.515 ;
        RECT 45.745 125.470 46.035 125.515 ;
        RECT 42.035 125.330 46.035 125.470 ;
        RECT 42.035 125.285 42.325 125.330 ;
        RECT 44.555 125.285 44.845 125.330 ;
        RECT 45.745 125.285 46.035 125.330 ;
        RECT 58.545 125.470 58.835 125.515 ;
        RECT 59.735 125.470 60.025 125.515 ;
        RECT 62.255 125.470 62.545 125.515 ;
        RECT 58.545 125.330 62.545 125.470 ;
        RECT 58.545 125.285 58.835 125.330 ;
        RECT 59.735 125.285 60.025 125.330 ;
        RECT 62.255 125.285 62.545 125.330 ;
        RECT 66.390 125.270 66.710 125.530 ;
        RECT 91.230 125.470 91.550 125.530 ;
        RECT 91.705 125.470 91.995 125.515 ;
        RECT 91.230 125.330 91.995 125.470 ;
        RECT 91.230 125.270 91.550 125.330 ;
        RECT 91.705 125.285 91.995 125.330 ;
        RECT 41.550 125.130 41.870 125.190 ;
        RECT 46.625 125.130 46.915 125.175 ;
        RECT 57.665 125.130 57.955 125.175 ;
        RECT 64.550 125.130 64.870 125.190 ;
        RECT 41.550 124.990 47.760 125.130 ;
        RECT 41.550 124.930 41.870 124.990 ;
        RECT 46.625 124.945 46.915 124.990 ;
        RECT 45.230 124.835 45.550 124.850 ;
        RECT 45.230 124.790 45.580 124.835 ;
        RECT 45.230 124.650 45.745 124.790 ;
        RECT 45.230 124.605 45.580 124.650 ;
        RECT 45.230 124.590 45.550 124.605 ;
        RECT 47.620 124.510 47.760 124.990 ;
        RECT 57.665 124.990 64.870 125.130 ;
        RECT 57.665 124.945 57.955 124.990 ;
        RECT 64.550 124.930 64.870 124.990 ;
        RECT 65.485 125.130 65.775 125.175 ;
        RECT 66.480 125.130 66.620 125.270 ;
        RECT 65.485 124.990 66.620 125.130 ;
        RECT 94.925 125.130 95.215 125.175 ;
        RECT 95.385 125.130 95.675 125.175 ;
        RECT 94.925 124.990 95.675 125.130 ;
        RECT 65.485 124.945 65.775 124.990 ;
        RECT 94.925 124.945 95.215 124.990 ;
        RECT 95.385 124.945 95.675 124.990 ;
        RECT 96.290 124.930 96.610 125.190 ;
        RECT 59.030 124.835 59.350 124.850 ;
        RECT 59.000 124.790 59.350 124.835 ;
        RECT 58.835 124.650 59.350 124.790 ;
        RECT 59.000 124.605 59.350 124.650 ;
        RECT 59.030 124.590 59.350 124.605 ;
        RECT 47.530 124.250 47.850 124.510 ;
        RECT 11.120 123.630 151.295 124.110 ;
        RECT 54.430 123.230 54.750 123.490 ;
        RECT 48.880 123.090 49.170 123.135 ;
        RECT 49.370 123.090 49.690 123.150 ;
        RECT 48.880 122.950 49.690 123.090 ;
        RECT 48.880 122.905 49.170 122.950 ;
        RECT 49.370 122.890 49.690 122.950 ;
        RECT 47.530 122.550 47.850 122.810 ;
        RECT 48.425 122.410 48.715 122.455 ;
        RECT 49.615 122.410 49.905 122.455 ;
        RECT 52.135 122.410 52.425 122.455 ;
        RECT 48.425 122.270 52.425 122.410 ;
        RECT 48.425 122.225 48.715 122.270 ;
        RECT 49.615 122.225 49.905 122.270 ;
        RECT 52.135 122.225 52.425 122.270 ;
        RECT 48.030 122.070 48.320 122.115 ;
        RECT 50.130 122.070 50.420 122.115 ;
        RECT 51.700 122.070 51.990 122.115 ;
        RECT 48.030 121.930 51.990 122.070 ;
        RECT 48.030 121.885 48.320 121.930 ;
        RECT 50.130 121.885 50.420 121.930 ;
        RECT 51.700 121.885 51.990 121.930 ;
        RECT 11.120 120.910 150.500 121.390 ;
        RECT 11.120 118.190 151.295 118.670 ;
        RECT 11.120 115.470 150.500 115.950 ;
        RECT 11.120 112.750 151.295 113.230 ;
        RECT 11.120 110.030 150.500 110.510 ;
        RECT 11.120 107.310 151.295 107.790 ;
        RECT 11.120 104.590 150.500 105.070 ;
        RECT 11.120 101.870 151.295 102.350 ;
        RECT 11.120 99.150 150.500 99.630 ;
        RECT 11.120 96.430 151.295 96.910 ;
        RECT 11.120 93.710 150.500 94.190 ;
        RECT 11.120 90.990 151.295 91.470 ;
        RECT 11.120 88.270 150.500 88.750 ;
        RECT 11.120 85.550 151.295 86.030 ;
        RECT 11.120 82.830 150.500 83.310 ;
        RECT 11.120 80.110 151.295 80.590 ;
        RECT 11.120 77.390 150.500 77.870 ;
        RECT 11.120 74.670 151.295 75.150 ;
        RECT 54.810 56.250 77.300 59.710 ;
        RECT 54.810 52.430 77.350 56.250 ;
        RECT 54.810 50.390 84.840 52.430 ;
        RECT 95.020 51.750 105.690 60.270 ;
        RECT 117.080 52.030 134.980 58.630 ;
        RECT 94.700 50.580 105.900 51.750 ;
        RECT 54.840 50.350 84.840 50.390 ;
        RECT 54.840 50.340 77.780 50.350 ;
        RECT 54.840 37.380 60.790 50.340 ;
        RECT 61.530 49.540 63.410 50.340 ;
        RECT 61.910 49.290 63.030 49.540 ;
        RECT 64.200 49.490 66.080 50.340 ;
        RECT 64.630 49.300 65.640 49.490 ;
        RECT 64.635 49.290 65.635 49.300 ;
        RECT 63.210 49.240 64.390 49.270 ;
        RECT 61.540 49.030 61.770 49.240 ;
        RECT 61.540 49.020 61.780 49.030 ;
        RECT 61.530 48.370 61.780 49.020 ;
        RECT 63.180 48.370 64.430 49.240 ;
        RECT 65.840 48.370 66.070 49.240 ;
        RECT 61.530 48.190 66.070 48.370 ;
        RECT 61.530 48.110 61.780 48.190 ;
        RECT 61.530 47.230 61.770 48.110 ;
        RECT 63.180 47.280 64.430 48.190 ;
        RECT 65.840 47.280 66.070 48.190 ;
        RECT 66.710 47.690 77.780 50.340 ;
        RECT 78.310 49.875 80.180 50.105 ;
        RECT 80.950 49.890 84.840 50.350 ;
        RECT 78.310 48.770 78.540 49.875 ;
        RECT 78.710 49.160 79.800 49.640 ;
        RECT 78.330 48.440 78.520 48.770 ;
        RECT 78.310 47.980 78.540 48.440 ;
        RECT 78.710 48.380 79.800 48.860 ;
        RECT 79.950 48.770 80.180 49.875 ;
        RECT 79.970 48.440 80.160 48.770 ;
        RECT 78.330 47.650 78.520 47.980 ;
        RECT 78.310 47.460 78.540 47.650 ;
        RECT 78.700 47.580 79.790 48.060 ;
        RECT 79.950 47.980 80.180 48.440 ;
        RECT 79.970 47.650 80.160 47.980 ;
        RECT 78.060 47.410 78.540 47.460 ;
        RECT 77.890 47.310 78.540 47.410 ;
        RECT 63.180 47.230 64.390 47.280 ;
        RECT 61.530 47.000 64.390 47.230 ;
        RECT 61.530 46.200 61.770 47.000 ;
        RECT 63.180 46.950 64.390 47.000 ;
        RECT 63.180 46.200 64.430 46.950 ;
        RECT 64.580 46.910 65.690 47.280 ;
        RECT 77.490 47.190 78.540 47.310 ;
        RECT 65.840 46.200 66.070 46.950 ;
        RECT 77.490 46.870 78.520 47.190 ;
        RECT 77.890 46.860 78.520 46.870 ;
        RECT 77.890 46.710 78.540 46.860 ;
        RECT 78.700 46.800 79.790 47.280 ;
        RECT 79.950 47.190 80.180 47.650 ;
        RECT 80.960 47.560 83.000 49.890 ;
        RECT 79.970 46.860 80.160 47.190 ;
        RECT 99.970 47.000 100.980 50.580 ;
        RECT 117.070 49.950 147.070 52.030 ;
        RECT 117.070 49.940 140.010 49.950 ;
        RECT 78.310 46.400 78.540 46.710 ;
        RECT 61.530 46.020 66.070 46.200 ;
        RECT 78.330 46.070 78.520 46.400 ;
        RECT 61.530 45.850 61.780 46.020 ;
        RECT 61.530 44.960 61.770 45.850 ;
        RECT 61.530 44.710 61.780 44.960 ;
        RECT 61.530 43.850 61.770 44.710 ;
        RECT 61.950 44.650 62.990 45.010 ;
        RECT 63.180 44.990 64.430 46.020 ;
        RECT 63.190 44.660 64.390 44.990 ;
        RECT 61.530 43.810 61.780 43.850 ;
        RECT 63.180 43.810 64.430 44.660 ;
        RECT 64.630 44.630 65.640 45.030 ;
        RECT 65.840 44.990 66.070 46.020 ;
        RECT 78.310 45.610 78.540 46.070 ;
        RECT 78.690 46.010 79.780 46.490 ;
        RECT 79.950 46.400 80.180 46.860 ;
        RECT 79.970 46.070 80.160 46.400 ;
        RECT 78.330 45.280 78.520 45.610 ;
        RECT 78.310 44.820 78.540 45.280 ;
        RECT 78.700 45.210 79.790 45.690 ;
        RECT 79.950 45.610 80.180 46.070 ;
        RECT 79.970 45.280 80.160 45.610 ;
        RECT 65.840 43.810 66.070 44.660 ;
        RECT 78.330 44.490 78.520 44.820 ;
        RECT 78.310 44.030 78.540 44.490 ;
        RECT 78.720 44.420 79.810 44.900 ;
        RECT 79.950 44.820 80.180 45.280 ;
        RECT 79.970 44.490 80.160 44.820 ;
        RECT 61.530 43.630 66.070 43.810 ;
        RECT 78.330 43.700 78.520 44.030 ;
        RECT 61.530 43.550 61.780 43.630 ;
        RECT 61.530 42.640 61.770 43.550 ;
        RECT 63.180 42.700 64.430 43.630 ;
        RECT 61.975 42.640 62.975 42.650 ;
        RECT 63.180 42.640 64.390 42.700 ;
        RECT 61.530 42.410 64.390 42.640 ;
        RECT 61.530 41.620 61.770 42.410 ;
        RECT 63.180 42.370 64.390 42.410 ;
        RECT 61.530 41.600 61.780 41.620 ;
        RECT 63.180 41.600 64.430 42.370 ;
        RECT 64.580 42.350 65.690 42.720 ;
        RECT 65.840 42.700 66.070 43.630 ;
        RECT 78.310 43.240 78.540 43.700 ;
        RECT 78.710 43.640 79.800 44.120 ;
        RECT 79.950 44.030 80.180 44.490 ;
        RECT 79.970 43.700 80.160 44.030 ;
        RECT 78.330 42.910 78.520 43.240 ;
        RECT 78.310 42.450 78.540 42.910 ;
        RECT 78.720 42.840 79.810 43.320 ;
        RECT 79.950 43.240 80.180 43.700 ;
        RECT 99.930 43.470 100.870 44.560 ;
        RECT 106.985 43.470 108.715 43.500 ;
        RECT 79.970 42.910 80.160 43.240 ;
        RECT 65.840 41.600 66.070 42.370 ;
        RECT 61.530 41.420 66.070 41.600 ;
        RECT 61.530 41.320 61.780 41.420 ;
        RECT 61.530 40.370 61.770 41.320 ;
        RECT 61.530 40.120 61.780 40.370 ;
        RECT 61.530 39.340 61.770 40.120 ;
        RECT 61.960 40.080 63.000 40.440 ;
        RECT 63.180 40.410 64.430 41.420 ;
        RECT 63.190 40.080 64.390 40.410 ;
        RECT 64.620 40.360 65.630 40.460 ;
        RECT 65.840 40.410 66.070 41.420 ;
        RECT 73.170 41.260 73.400 42.070 ;
        RECT 73.560 42.040 74.570 42.400 ;
        RECT 78.330 42.120 78.520 42.450 ;
        RECT 74.720 41.260 74.950 42.070 ;
        RECT 78.310 41.660 78.540 42.120 ;
        RECT 78.710 42.060 79.800 42.540 ;
        RECT 79.950 42.450 80.180 42.910 ;
        RECT 79.970 42.120 80.160 42.450 ;
        RECT 78.330 41.330 78.520 41.660 ;
        RECT 73.170 40.970 74.950 41.260 ;
        RECT 64.620 40.130 65.635 40.360 ;
        RECT 62.020 40.060 62.930 40.080 ;
        RECT 61.530 39.160 61.780 39.340 ;
        RECT 63.180 39.160 64.430 40.080 ;
        RECT 64.620 40.060 65.630 40.130 ;
        RECT 73.170 40.110 73.400 40.970 ;
        RECT 65.840 39.160 66.070 40.080 ;
        RECT 73.190 39.780 73.360 40.110 ;
        RECT 61.530 38.980 66.070 39.160 ;
        RECT 61.530 38.070 61.770 38.980 ;
        RECT 63.180 38.120 64.430 38.980 ;
        RECT 63.180 38.070 64.390 38.120 ;
        RECT 61.530 37.840 64.390 38.070 ;
        RECT 61.530 36.930 61.770 37.840 ;
        RECT 63.180 37.790 64.390 37.840 ;
        RECT 61.530 36.900 61.780 36.930 ;
        RECT 63.180 36.900 64.430 37.790 ;
        RECT 64.580 37.770 65.690 38.140 ;
        RECT 65.840 38.120 66.070 38.980 ;
        RECT 73.170 38.930 73.400 39.780 ;
        RECT 73.540 39.750 74.580 40.140 ;
        RECT 74.720 40.110 74.950 40.970 ;
        RECT 78.310 40.870 78.540 41.330 ;
        RECT 78.720 41.260 79.810 41.740 ;
        RECT 79.950 41.660 80.180 42.120 ;
        RECT 99.930 41.740 108.715 43.470 ;
        RECT 79.970 41.330 80.160 41.660 ;
        RECT 78.330 40.540 78.520 40.870 ;
        RECT 74.760 39.780 74.900 40.110 ;
        RECT 78.310 40.080 78.540 40.540 ;
        RECT 78.710 40.480 79.800 40.960 ;
        RECT 79.950 40.870 80.180 41.330 ;
        RECT 79.970 40.540 80.160 40.870 ;
        RECT 99.930 40.710 100.870 41.740 ;
        RECT 106.985 41.710 108.715 41.740 ;
        RECT 74.720 38.930 74.950 39.780 ;
        RECT 78.330 39.750 78.520 40.080 ;
        RECT 78.310 39.290 78.540 39.750 ;
        RECT 78.700 39.680 79.790 40.160 ;
        RECT 79.950 40.080 80.180 40.540 ;
        RECT 97.370 40.160 103.120 40.710 ;
        RECT 97.340 40.150 103.120 40.160 ;
        RECT 79.970 39.750 80.160 40.080 ;
        RECT 97.340 39.810 103.160 40.150 ;
        RECT 78.330 38.960 78.520 39.290 ;
        RECT 73.170 38.640 74.950 38.930 ;
        RECT 73.170 37.820 73.400 38.640 ;
        RECT 65.840 36.900 66.070 37.790 ;
        RECT 73.190 37.490 73.360 37.820 ;
        RECT 73.550 37.490 74.560 37.850 ;
        RECT 74.720 37.820 74.950 38.640 ;
        RECT 78.310 38.500 78.540 38.960 ;
        RECT 78.710 38.900 79.800 39.380 ;
        RECT 79.950 39.290 80.180 39.750 ;
        RECT 97.340 39.480 98.600 39.810 ;
        RECT 101.900 39.480 103.160 39.810 ;
        RECT 79.970 38.960 80.160 39.290 ;
        RECT 95.790 39.250 100.040 39.480 ;
        RECT 100.370 39.250 104.620 39.480 ;
        RECT 78.330 38.170 78.520 38.500 ;
        RECT 74.760 37.490 74.900 37.820 ;
        RECT 78.310 37.710 78.540 38.170 ;
        RECT 78.710 38.100 79.800 38.580 ;
        RECT 79.950 38.500 80.180 38.960 ;
        RECT 79.970 38.170 80.160 38.500 ;
        RECT 61.530 36.720 66.070 36.900 ;
        RECT 61.530 36.630 61.780 36.720 ;
        RECT 61.530 35.920 61.770 36.630 ;
        RECT 61.530 35.020 61.780 35.920 ;
        RECT 62.020 35.840 62.930 35.850 ;
        RECT 61.980 35.780 62.990 35.840 ;
        RECT 61.975 35.550 62.990 35.780 ;
        RECT 61.980 35.540 62.990 35.550 ;
        RECT 63.180 35.830 64.430 36.720 ;
        RECT 63.180 35.640 64.390 35.830 ;
        RECT 64.640 35.780 65.640 35.840 ;
        RECT 65.840 35.830 66.070 36.720 ;
        RECT 73.170 36.660 73.400 37.490 ;
        RECT 74.720 36.660 74.950 37.490 ;
        RECT 78.330 37.380 78.520 37.710 ;
        RECT 78.310 36.920 78.540 37.380 ;
        RECT 78.710 37.310 79.800 37.790 ;
        RECT 79.950 37.710 80.180 38.170 ;
        RECT 95.060 38.110 96.160 39.110 ;
        RECT 95.510 38.090 95.740 38.110 ;
        RECT 96.620 37.930 99.110 39.250 ;
        RECT 100.090 39.070 100.320 39.090 ;
        RECT 99.640 38.070 100.740 39.070 ;
        RECT 101.220 37.930 103.740 39.250 ;
        RECT 104.190 38.090 105.290 39.090 ;
        RECT 95.790 37.780 100.040 37.930 ;
        RECT 79.970 37.380 80.160 37.710 ;
        RECT 95.790 37.700 97.750 37.780 ;
        RECT 98.080 37.700 100.040 37.780 ;
        RECT 100.370 37.820 104.620 37.930 ;
        RECT 100.370 37.700 102.330 37.820 ;
        RECT 102.660 37.700 104.620 37.820 ;
        RECT 73.170 36.370 74.950 36.660 ;
        RECT 78.330 36.590 78.520 36.920 ;
        RECT 62.020 35.500 62.930 35.540 ;
        RECT 63.180 35.020 63.430 35.640 ;
        RECT 64.635 35.550 65.640 35.780 ;
        RECT 64.640 35.490 65.640 35.550 ;
        RECT 73.170 35.530 73.400 36.370 ;
        RECT 64.670 35.470 65.600 35.490 ;
        RECT 73.190 35.210 73.350 35.530 ;
        RECT 73.190 35.200 73.390 35.210 ;
        RECT 61.530 34.680 63.700 35.020 ;
        RECT 64.710 34.690 65.840 35.110 ;
        RECT 62.570 33.570 63.070 33.860 ;
        RECT 61.940 30.910 62.540 33.420 ;
        RECT 62.680 30.750 62.960 33.570 ;
        RECT 63.310 33.420 63.700 34.680 ;
        RECT 64.500 33.550 65.010 33.850 ;
        RECT 63.100 30.910 63.700 33.420 ;
        RECT 63.870 33.030 64.470 33.410 ;
        RECT 63.840 31.040 64.470 33.030 ;
        RECT 63.870 30.910 64.470 31.040 ;
        RECT 64.610 30.750 64.890 33.550 ;
        RECT 65.250 33.410 65.630 34.690 ;
        RECT 73.170 34.340 73.400 35.200 ;
        RECT 73.540 35.110 74.580 35.620 ;
        RECT 74.720 35.530 74.950 36.370 ;
        RECT 78.310 36.130 78.540 36.590 ;
        RECT 78.720 36.520 79.810 37.000 ;
        RECT 79.950 36.920 80.180 37.380 ;
        RECT 79.970 36.590 80.160 36.920 ;
        RECT 78.330 35.800 78.520 36.130 ;
        RECT 74.760 35.200 74.900 35.530 ;
        RECT 78.310 35.340 78.540 35.800 ;
        RECT 78.710 35.730 79.800 36.210 ;
        RECT 79.950 36.130 80.180 36.590 ;
        RECT 79.970 35.800 80.160 36.130 ;
        RECT 74.720 34.340 74.950 35.200 ;
        RECT 78.330 35.010 78.520 35.340 ;
        RECT 78.310 34.550 78.540 35.010 ;
        RECT 78.720 34.950 79.810 35.430 ;
        RECT 79.950 35.340 80.180 35.800 ;
        RECT 94.870 35.440 106.020 37.020 ;
        RECT 117.070 36.980 123.020 49.940 ;
        RECT 123.760 49.140 125.640 49.940 ;
        RECT 124.140 48.890 125.260 49.140 ;
        RECT 126.430 49.090 128.310 49.940 ;
        RECT 126.860 48.900 127.870 49.090 ;
        RECT 126.865 48.890 127.865 48.900 ;
        RECT 125.440 48.840 126.620 48.870 ;
        RECT 123.770 48.630 124.000 48.840 ;
        RECT 123.770 48.620 124.010 48.630 ;
        RECT 123.760 47.970 124.010 48.620 ;
        RECT 125.410 47.970 126.660 48.840 ;
        RECT 128.070 47.970 128.300 48.840 ;
        RECT 123.760 47.790 128.300 47.970 ;
        RECT 123.760 47.710 124.010 47.790 ;
        RECT 123.760 46.830 124.000 47.710 ;
        RECT 125.410 46.880 126.660 47.790 ;
        RECT 128.070 46.880 128.300 47.790 ;
        RECT 128.940 47.290 140.010 49.940 ;
        RECT 140.540 49.475 142.410 49.705 ;
        RECT 143.180 49.490 147.070 49.950 ;
        RECT 140.540 48.370 140.770 49.475 ;
        RECT 140.940 48.760 142.030 49.240 ;
        RECT 140.560 48.040 140.750 48.370 ;
        RECT 140.540 47.580 140.770 48.040 ;
        RECT 140.940 47.980 142.030 48.460 ;
        RECT 142.180 48.370 142.410 49.475 ;
        RECT 142.200 48.040 142.390 48.370 ;
        RECT 140.560 47.250 140.750 47.580 ;
        RECT 140.540 47.060 140.770 47.250 ;
        RECT 140.930 47.180 142.020 47.660 ;
        RECT 142.180 47.580 142.410 48.040 ;
        RECT 142.200 47.250 142.390 47.580 ;
        RECT 140.290 47.010 140.770 47.060 ;
        RECT 140.120 46.910 140.770 47.010 ;
        RECT 125.410 46.830 126.620 46.880 ;
        RECT 123.760 46.600 126.620 46.830 ;
        RECT 123.760 45.800 124.000 46.600 ;
        RECT 125.410 46.550 126.620 46.600 ;
        RECT 125.410 45.800 126.660 46.550 ;
        RECT 126.810 46.510 127.920 46.880 ;
        RECT 139.720 46.790 140.770 46.910 ;
        RECT 128.070 45.800 128.300 46.550 ;
        RECT 139.720 46.470 140.750 46.790 ;
        RECT 140.120 46.460 140.750 46.470 ;
        RECT 140.120 46.310 140.770 46.460 ;
        RECT 140.930 46.400 142.020 46.880 ;
        RECT 142.180 46.790 142.410 47.250 ;
        RECT 143.190 47.160 145.230 49.490 ;
        RECT 142.200 46.460 142.390 46.790 ;
        RECT 140.540 46.000 140.770 46.310 ;
        RECT 123.760 45.620 128.300 45.800 ;
        RECT 140.560 45.670 140.750 46.000 ;
        RECT 123.760 45.450 124.010 45.620 ;
        RECT 123.760 44.560 124.000 45.450 ;
        RECT 123.760 44.310 124.010 44.560 ;
        RECT 123.760 43.450 124.000 44.310 ;
        RECT 124.180 44.250 125.220 44.610 ;
        RECT 125.410 44.590 126.660 45.620 ;
        RECT 125.420 44.260 126.620 44.590 ;
        RECT 123.760 43.410 124.010 43.450 ;
        RECT 125.410 43.410 126.660 44.260 ;
        RECT 126.860 44.230 127.870 44.630 ;
        RECT 128.070 44.590 128.300 45.620 ;
        RECT 140.540 45.210 140.770 45.670 ;
        RECT 140.920 45.610 142.010 46.090 ;
        RECT 142.180 46.000 142.410 46.460 ;
        RECT 142.200 45.670 142.390 46.000 ;
        RECT 140.560 44.880 140.750 45.210 ;
        RECT 140.540 44.420 140.770 44.880 ;
        RECT 140.930 44.810 142.020 45.290 ;
        RECT 142.180 45.210 142.410 45.670 ;
        RECT 142.200 44.880 142.390 45.210 ;
        RECT 128.070 43.410 128.300 44.260 ;
        RECT 140.560 44.090 140.750 44.420 ;
        RECT 140.540 43.630 140.770 44.090 ;
        RECT 140.950 44.020 142.040 44.500 ;
        RECT 142.180 44.420 142.410 44.880 ;
        RECT 142.200 44.090 142.390 44.420 ;
        RECT 123.760 43.230 128.300 43.410 ;
        RECT 140.560 43.300 140.750 43.630 ;
        RECT 123.760 43.150 124.010 43.230 ;
        RECT 123.760 42.240 124.000 43.150 ;
        RECT 125.410 42.300 126.660 43.230 ;
        RECT 124.205 42.240 125.205 42.250 ;
        RECT 125.410 42.240 126.620 42.300 ;
        RECT 123.760 42.010 126.620 42.240 ;
        RECT 123.760 41.220 124.000 42.010 ;
        RECT 125.410 41.970 126.620 42.010 ;
        RECT 123.760 41.200 124.010 41.220 ;
        RECT 125.410 41.200 126.660 41.970 ;
        RECT 126.810 41.950 127.920 42.320 ;
        RECT 128.070 42.300 128.300 43.230 ;
        RECT 140.540 42.840 140.770 43.300 ;
        RECT 140.940 43.240 142.030 43.720 ;
        RECT 142.180 43.630 142.410 44.090 ;
        RECT 142.200 43.300 142.390 43.630 ;
        RECT 140.560 42.510 140.750 42.840 ;
        RECT 140.540 42.050 140.770 42.510 ;
        RECT 140.950 42.440 142.040 42.920 ;
        RECT 142.180 42.840 142.410 43.300 ;
        RECT 142.200 42.510 142.390 42.840 ;
        RECT 128.070 41.200 128.300 41.970 ;
        RECT 123.760 41.020 128.300 41.200 ;
        RECT 123.760 40.920 124.010 41.020 ;
        RECT 123.760 39.970 124.000 40.920 ;
        RECT 123.760 39.720 124.010 39.970 ;
        RECT 123.760 38.940 124.000 39.720 ;
        RECT 124.190 39.680 125.230 40.040 ;
        RECT 125.410 40.010 126.660 41.020 ;
        RECT 125.420 39.680 126.620 40.010 ;
        RECT 126.850 39.960 127.860 40.060 ;
        RECT 128.070 40.010 128.300 41.020 ;
        RECT 135.400 40.860 135.630 41.670 ;
        RECT 135.790 41.640 136.800 42.000 ;
        RECT 140.560 41.720 140.750 42.050 ;
        RECT 136.950 40.860 137.180 41.670 ;
        RECT 140.540 41.260 140.770 41.720 ;
        RECT 140.940 41.660 142.030 42.140 ;
        RECT 142.180 42.050 142.410 42.510 ;
        RECT 142.200 41.720 142.390 42.050 ;
        RECT 140.560 40.930 140.750 41.260 ;
        RECT 135.400 40.570 137.180 40.860 ;
        RECT 126.850 39.730 127.865 39.960 ;
        RECT 124.250 39.660 125.160 39.680 ;
        RECT 123.760 38.760 124.010 38.940 ;
        RECT 125.410 38.760 126.660 39.680 ;
        RECT 126.850 39.660 127.860 39.730 ;
        RECT 135.400 39.710 135.630 40.570 ;
        RECT 128.070 38.760 128.300 39.680 ;
        RECT 135.420 39.380 135.590 39.710 ;
        RECT 123.760 38.580 128.300 38.760 ;
        RECT 123.760 37.670 124.000 38.580 ;
        RECT 125.410 37.720 126.660 38.580 ;
        RECT 125.410 37.670 126.620 37.720 ;
        RECT 123.760 37.440 126.620 37.670 ;
        RECT 123.760 36.530 124.000 37.440 ;
        RECT 125.410 37.390 126.620 37.440 ;
        RECT 123.760 36.500 124.010 36.530 ;
        RECT 125.410 36.500 126.660 37.390 ;
        RECT 126.810 37.370 127.920 37.740 ;
        RECT 128.070 37.720 128.300 38.580 ;
        RECT 135.400 38.530 135.630 39.380 ;
        RECT 135.770 39.350 136.810 39.740 ;
        RECT 136.950 39.710 137.180 40.570 ;
        RECT 140.540 40.470 140.770 40.930 ;
        RECT 140.950 40.860 142.040 41.340 ;
        RECT 142.180 41.260 142.410 41.720 ;
        RECT 142.200 40.930 142.390 41.260 ;
        RECT 140.560 40.140 140.750 40.470 ;
        RECT 136.990 39.380 137.130 39.710 ;
        RECT 140.540 39.680 140.770 40.140 ;
        RECT 140.940 40.080 142.030 40.560 ;
        RECT 142.180 40.470 142.410 40.930 ;
        RECT 142.200 40.140 142.390 40.470 ;
        RECT 136.950 38.530 137.180 39.380 ;
        RECT 140.560 39.350 140.750 39.680 ;
        RECT 140.540 38.890 140.770 39.350 ;
        RECT 140.930 39.280 142.020 39.760 ;
        RECT 142.180 39.680 142.410 40.140 ;
        RECT 142.200 39.350 142.390 39.680 ;
        RECT 140.560 38.560 140.750 38.890 ;
        RECT 135.400 38.240 137.180 38.530 ;
        RECT 135.400 37.420 135.630 38.240 ;
        RECT 128.070 36.500 128.300 37.390 ;
        RECT 135.420 37.090 135.590 37.420 ;
        RECT 135.780 37.090 136.790 37.450 ;
        RECT 136.950 37.420 137.180 38.240 ;
        RECT 140.540 38.100 140.770 38.560 ;
        RECT 140.940 38.500 142.030 38.980 ;
        RECT 142.180 38.890 142.410 39.350 ;
        RECT 142.200 38.560 142.390 38.890 ;
        RECT 140.560 37.770 140.750 38.100 ;
        RECT 136.990 37.090 137.130 37.420 ;
        RECT 140.540 37.310 140.770 37.770 ;
        RECT 140.940 37.700 142.030 38.180 ;
        RECT 142.180 38.100 142.410 38.560 ;
        RECT 142.200 37.770 142.390 38.100 ;
        RECT 123.760 36.320 128.300 36.500 ;
        RECT 123.760 36.230 124.010 36.320 ;
        RECT 123.760 35.520 124.000 36.230 ;
        RECT 79.970 35.010 80.160 35.340 ;
        RECT 73.170 34.155 74.950 34.340 ;
        RECT 78.330 34.220 78.520 34.550 ;
        RECT 65.030 30.900 65.630 33.410 ;
        RECT 68.025 34.050 74.950 34.155 ;
        RECT 68.025 33.240 73.400 34.050 ;
        RECT 74.720 33.240 74.950 34.050 ;
        RECT 78.310 33.760 78.540 34.220 ;
        RECT 78.710 34.140 79.800 34.620 ;
        RECT 79.950 34.550 80.180 35.010 ;
        RECT 79.970 34.220 80.160 34.550 ;
        RECT 79.950 33.760 80.180 34.220 ;
        RECT 78.330 33.720 78.520 33.760 ;
        RECT 78.710 33.320 79.770 33.760 ;
        RECT 79.970 33.750 80.160 33.760 ;
        RECT 68.025 33.180 73.360 33.240 ;
        RECT 54.870 28.585 56.020 30.450 ;
        RECT 62.570 29.370 63.070 30.750 ;
        RECT 64.500 30.140 65.000 30.750 ;
        RECT 66.615 30.140 67.210 30.260 ;
        RECT 64.500 29.730 67.210 30.140 ;
        RECT 66.615 29.605 67.210 29.730 ;
        RECT 62.570 28.790 64.810 29.370 ;
        RECT 68.025 28.585 69.000 33.180 ;
        RECT 73.190 32.910 73.360 33.180 ;
        RECT 73.540 32.950 74.580 33.210 ;
        RECT 74.760 32.910 74.900 33.240 ;
        RECT 73.170 32.100 73.400 32.910 ;
        RECT 74.720 32.100 74.950 32.910 ;
        RECT 73.170 31.810 74.950 32.100 ;
        RECT 73.170 30.950 73.400 31.810 ;
        RECT 73.190 30.620 73.360 30.950 ;
        RECT 73.170 29.760 73.400 30.620 ;
        RECT 73.540 30.580 74.580 30.970 ;
        RECT 74.720 30.950 74.950 31.810 ;
        RECT 74.760 30.620 74.900 30.950 ;
        RECT 74.720 29.760 74.950 30.620 ;
        RECT 73.170 29.470 74.950 29.760 ;
        RECT 73.170 28.660 73.400 29.470 ;
        RECT 74.720 28.660 74.950 29.470 ;
        RECT 54.870 27.730 69.000 28.585 ;
        RECT 73.190 28.330 73.360 28.660 ;
        RECT 73.540 28.360 74.580 28.630 ;
        RECT 74.760 28.330 74.900 28.660 ;
        RECT 54.880 27.725 69.000 27.730 ;
        RECT 54.880 27.720 68.570 27.725 ;
        RECT 56.260 27.030 57.010 27.720 ;
        RECT 73.170 27.490 73.400 28.330 ;
        RECT 74.720 27.490 74.950 28.330 ;
        RECT 73.170 27.200 74.950 27.490 ;
        RECT 56.260 26.860 63.990 27.030 ;
        RECT 55.850 26.660 64.680 26.860 ;
        RECT 55.850 26.630 57.810 26.660 ;
        RECT 58.140 26.630 60.100 26.660 ;
        RECT 60.430 26.630 62.390 26.660 ;
        RECT 62.720 26.630 64.680 26.660 ;
        RECT 55.490 25.470 55.850 26.470 ;
        RECT 56.630 25.310 57.010 26.630 ;
        RECT 57.790 25.470 58.170 26.470 ;
        RECT 58.940 25.310 59.320 26.630 ;
        RECT 60.070 25.470 60.450 26.470 ;
        RECT 61.180 25.310 61.560 26.630 ;
        RECT 62.360 25.470 62.740 26.470 ;
        RECT 63.520 25.310 63.900 26.630 ;
        RECT 64.660 25.470 65.040 26.470 ;
        RECT 73.170 26.370 73.400 27.200 ;
        RECT 73.540 26.060 74.580 26.400 ;
        RECT 74.720 26.370 74.950 27.200 ;
        RECT 74.760 26.330 74.900 26.370 ;
        RECT 73.560 25.660 74.560 26.060 ;
        RECT 55.850 25.080 57.810 25.310 ;
        RECT 58.140 25.080 60.100 25.310 ;
        RECT 60.430 25.080 62.390 25.310 ;
        RECT 62.720 25.080 64.680 25.310 ;
        RECT 65.530 24.480 84.840 25.660 ;
        RECT 54.840 10.670 84.840 24.480 ;
        RECT 94.300 10.990 106.280 35.440 ;
        RECT 123.760 34.620 124.010 35.520 ;
        RECT 124.250 35.440 125.160 35.450 ;
        RECT 124.210 35.380 125.220 35.440 ;
        RECT 124.205 35.150 125.220 35.380 ;
        RECT 124.210 35.140 125.220 35.150 ;
        RECT 125.410 35.430 126.660 36.320 ;
        RECT 125.410 35.240 126.620 35.430 ;
        RECT 126.870 35.380 127.870 35.440 ;
        RECT 128.070 35.430 128.300 36.320 ;
        RECT 135.400 36.260 135.630 37.090 ;
        RECT 136.950 36.260 137.180 37.090 ;
        RECT 140.560 36.980 140.750 37.310 ;
        RECT 140.540 36.520 140.770 36.980 ;
        RECT 140.940 36.910 142.030 37.390 ;
        RECT 142.180 37.310 142.410 37.770 ;
        RECT 142.200 36.980 142.390 37.310 ;
        RECT 135.400 35.970 137.180 36.260 ;
        RECT 140.560 36.190 140.750 36.520 ;
        RECT 124.250 35.100 125.160 35.140 ;
        RECT 125.410 34.620 125.660 35.240 ;
        RECT 126.865 35.150 127.870 35.380 ;
        RECT 126.870 35.090 127.870 35.150 ;
        RECT 135.400 35.130 135.630 35.970 ;
        RECT 126.900 35.070 127.830 35.090 ;
        RECT 135.420 34.810 135.580 35.130 ;
        RECT 135.420 34.800 135.620 34.810 ;
        RECT 123.760 34.280 125.930 34.620 ;
        RECT 126.940 34.290 128.070 34.710 ;
        RECT 124.800 33.170 125.300 33.460 ;
        RECT 124.170 30.510 124.770 33.020 ;
        RECT 124.910 30.350 125.190 33.170 ;
        RECT 125.540 33.020 125.930 34.280 ;
        RECT 126.730 33.150 127.240 33.450 ;
        RECT 125.330 30.510 125.930 33.020 ;
        RECT 126.100 32.630 126.700 33.010 ;
        RECT 126.070 30.640 126.700 32.630 ;
        RECT 126.100 30.510 126.700 30.640 ;
        RECT 126.840 30.350 127.120 33.150 ;
        RECT 127.480 33.010 127.860 34.290 ;
        RECT 135.400 33.940 135.630 34.800 ;
        RECT 135.770 34.710 136.810 35.220 ;
        RECT 136.950 35.130 137.180 35.970 ;
        RECT 140.540 35.730 140.770 36.190 ;
        RECT 140.950 36.120 142.040 36.600 ;
        RECT 142.180 36.520 142.410 36.980 ;
        RECT 142.200 36.190 142.390 36.520 ;
        RECT 140.560 35.400 140.750 35.730 ;
        RECT 136.990 34.800 137.130 35.130 ;
        RECT 140.540 34.940 140.770 35.400 ;
        RECT 140.940 35.330 142.030 35.810 ;
        RECT 142.180 35.730 142.410 36.190 ;
        RECT 142.200 35.400 142.390 35.730 ;
        RECT 136.950 33.940 137.180 34.800 ;
        RECT 140.560 34.610 140.750 34.940 ;
        RECT 140.540 34.150 140.770 34.610 ;
        RECT 140.950 34.550 142.040 35.030 ;
        RECT 142.180 34.940 142.410 35.400 ;
        RECT 142.200 34.610 142.390 34.940 ;
        RECT 135.400 33.755 137.180 33.940 ;
        RECT 140.560 33.820 140.750 34.150 ;
        RECT 127.260 30.500 127.860 33.010 ;
        RECT 130.255 33.650 137.180 33.755 ;
        RECT 130.255 32.840 135.630 33.650 ;
        RECT 136.950 32.840 137.180 33.650 ;
        RECT 140.540 33.360 140.770 33.820 ;
        RECT 140.940 33.740 142.030 34.220 ;
        RECT 142.180 34.150 142.410 34.610 ;
        RECT 142.200 33.820 142.390 34.150 ;
        RECT 142.180 33.360 142.410 33.820 ;
        RECT 140.560 33.320 140.750 33.360 ;
        RECT 140.940 32.920 142.000 33.360 ;
        RECT 142.200 33.350 142.390 33.360 ;
        RECT 130.255 32.780 135.590 32.840 ;
        RECT 117.100 28.185 118.250 30.050 ;
        RECT 124.800 28.970 125.300 30.350 ;
        RECT 126.730 29.740 127.230 30.350 ;
        RECT 128.845 29.740 129.440 29.860 ;
        RECT 126.730 29.330 129.440 29.740 ;
        RECT 128.845 29.205 129.440 29.330 ;
        RECT 124.800 28.390 127.040 28.970 ;
        RECT 130.255 28.185 131.230 32.780 ;
        RECT 135.420 32.510 135.590 32.780 ;
        RECT 135.770 32.550 136.810 32.810 ;
        RECT 136.990 32.510 137.130 32.840 ;
        RECT 135.400 31.700 135.630 32.510 ;
        RECT 136.950 31.700 137.180 32.510 ;
        RECT 135.400 31.410 137.180 31.700 ;
        RECT 135.400 30.550 135.630 31.410 ;
        RECT 135.420 30.220 135.590 30.550 ;
        RECT 135.400 29.360 135.630 30.220 ;
        RECT 135.770 30.180 136.810 30.570 ;
        RECT 136.950 30.550 137.180 31.410 ;
        RECT 136.990 30.220 137.130 30.550 ;
        RECT 136.950 29.360 137.180 30.220 ;
        RECT 135.400 29.070 137.180 29.360 ;
        RECT 135.400 28.260 135.630 29.070 ;
        RECT 136.950 28.260 137.180 29.070 ;
        RECT 117.100 27.330 131.230 28.185 ;
        RECT 135.420 27.930 135.590 28.260 ;
        RECT 135.770 27.960 136.810 28.230 ;
        RECT 136.990 27.930 137.130 28.260 ;
        RECT 117.110 27.325 131.230 27.330 ;
        RECT 117.110 27.320 130.800 27.325 ;
        RECT 118.490 26.630 119.240 27.320 ;
        RECT 135.400 27.090 135.630 27.930 ;
        RECT 136.950 27.090 137.180 27.930 ;
        RECT 135.400 26.800 137.180 27.090 ;
        RECT 118.490 26.460 126.220 26.630 ;
        RECT 118.080 26.260 126.910 26.460 ;
        RECT 118.080 26.230 120.040 26.260 ;
        RECT 120.370 26.230 122.330 26.260 ;
        RECT 122.660 26.230 124.620 26.260 ;
        RECT 124.950 26.230 126.910 26.260 ;
        RECT 117.720 25.070 118.080 26.070 ;
        RECT 118.860 24.910 119.240 26.230 ;
        RECT 120.020 25.070 120.400 26.070 ;
        RECT 121.170 24.910 121.550 26.230 ;
        RECT 122.300 25.070 122.680 26.070 ;
        RECT 123.410 24.910 123.790 26.230 ;
        RECT 124.590 25.070 124.970 26.070 ;
        RECT 125.750 24.910 126.130 26.230 ;
        RECT 126.890 25.070 127.270 26.070 ;
        RECT 135.400 25.970 135.630 26.800 ;
        RECT 135.770 25.660 136.810 26.000 ;
        RECT 136.950 25.970 137.180 26.800 ;
        RECT 136.990 25.930 137.130 25.970 ;
        RECT 135.790 25.260 136.790 25.660 ;
        RECT 118.080 24.680 120.040 24.910 ;
        RECT 120.370 24.680 122.330 24.910 ;
        RECT 122.660 24.680 124.620 24.910 ;
        RECT 124.950 24.680 126.910 24.910 ;
        RECT 127.760 24.080 147.070 25.260 ;
        RECT 117.070 23.460 147.070 24.080 ;
        RECT 117.070 22.030 147.050 23.460 ;
        RECT 117.100 12.950 146.870 22.030 ;
        RECT 117.100 12.940 127.920 12.950 ;
      LAYER via ;
        RECT 27.770 213.500 28.030 213.760 ;
        RECT 28.090 213.500 28.350 213.760 ;
        RECT 28.410 213.500 28.670 213.760 ;
        RECT 28.730 213.500 28.990 213.760 ;
        RECT 29.050 213.500 29.310 213.760 ;
        RECT 62.615 213.500 62.875 213.760 ;
        RECT 62.935 213.500 63.195 213.760 ;
        RECT 63.255 213.500 63.515 213.760 ;
        RECT 63.575 213.500 63.835 213.760 ;
        RECT 63.895 213.500 64.155 213.760 ;
        RECT 97.460 213.500 97.720 213.760 ;
        RECT 97.780 213.500 98.040 213.760 ;
        RECT 98.100 213.500 98.360 213.760 ;
        RECT 98.420 213.500 98.680 213.760 ;
        RECT 98.740 213.500 99.000 213.760 ;
        RECT 132.305 213.500 132.565 213.760 ;
        RECT 132.625 213.500 132.885 213.760 ;
        RECT 132.945 213.500 133.205 213.760 ;
        RECT 133.265 213.500 133.525 213.760 ;
        RECT 133.585 213.500 133.845 213.760 ;
        RECT 65.500 212.990 65.760 213.250 ;
        RECT 105.980 212.990 106.240 213.250 ;
        RECT 64.120 211.970 64.380 212.230 ;
        RECT 86.660 211.970 86.920 212.230 ;
        RECT 95.860 211.970 96.120 212.230 ;
        RECT 104.600 211.970 104.860 212.230 ;
        RECT 89.420 211.290 89.680 211.550 ;
        RECT 99.080 211.290 99.340 211.550 ;
        RECT 107.820 211.290 108.080 211.550 ;
        RECT 108.740 211.290 109.000 211.550 ;
        RECT 116.100 211.970 116.360 212.230 ;
        RECT 126.220 211.970 126.480 212.230 ;
        RECT 136.340 211.970 136.600 212.230 ;
        RECT 116.560 211.290 116.820 211.550 ;
        RECT 127.600 211.290 127.860 211.550 ;
        RECT 137.720 211.290 137.980 211.550 ;
        RECT 45.190 210.780 45.450 211.040 ;
        RECT 45.510 210.780 45.770 211.040 ;
        RECT 45.830 210.780 46.090 211.040 ;
        RECT 46.150 210.780 46.410 211.040 ;
        RECT 46.470 210.780 46.730 211.040 ;
        RECT 80.035 210.780 80.295 211.040 ;
        RECT 80.355 210.780 80.615 211.040 ;
        RECT 80.675 210.780 80.935 211.040 ;
        RECT 80.995 210.780 81.255 211.040 ;
        RECT 81.315 210.780 81.575 211.040 ;
        RECT 114.880 210.780 115.140 211.040 ;
        RECT 115.200 210.780 115.460 211.040 ;
        RECT 115.520 210.780 115.780 211.040 ;
        RECT 115.840 210.780 116.100 211.040 ;
        RECT 116.160 210.780 116.420 211.040 ;
        RECT 149.725 210.780 149.985 211.040 ;
        RECT 150.045 210.780 150.305 211.040 ;
        RECT 150.365 210.780 150.625 211.040 ;
        RECT 150.685 210.780 150.945 211.040 ;
        RECT 151.005 210.780 151.265 211.040 ;
        RECT 14.900 209.930 15.160 210.190 ;
        RECT 25.020 209.930 25.280 210.190 ;
        RECT 35.140 209.930 35.400 210.190 ;
        RECT 19.500 209.590 19.760 209.850 ;
        RECT 21.340 209.590 21.600 209.850 ;
        RECT 19.960 209.250 20.220 209.510 ;
        RECT 30.080 209.250 30.340 209.510 ;
        RECT 32.840 209.590 33.100 209.850 ;
        RECT 36.060 209.590 36.320 209.850 ;
        RECT 37.900 209.590 38.160 209.850 ;
        RECT 43.420 209.590 43.680 209.850 ;
        RECT 38.820 209.250 39.080 209.510 ;
        RECT 42.960 208.910 43.220 209.170 ;
        RECT 44.800 208.910 45.060 209.170 ;
        RECT 48.020 209.590 48.280 209.850 ;
        RECT 53.080 209.590 53.340 209.850 ;
        RECT 55.840 209.590 56.100 209.850 ;
        RECT 58.140 209.590 58.400 209.850 ;
        RECT 64.580 209.590 64.840 209.850 ;
        RECT 47.560 209.250 47.820 209.510 ;
        RECT 64.120 208.910 64.380 209.170 ;
        RECT 74.700 209.590 74.960 209.850 ;
        RECT 83.440 209.930 83.700 210.190 ;
        RECT 86.660 210.270 86.920 210.530 ;
        RECT 104.600 210.270 104.860 210.530 ;
        RECT 116.560 210.270 116.820 210.530 ;
        RECT 85.740 209.930 86.000 210.190 ;
        RECT 84.360 209.590 84.620 209.850 ;
        RECT 89.420 209.590 89.680 209.850 ;
        RECT 107.820 209.930 108.080 210.190 ;
        RECT 100.000 209.590 100.260 209.850 ;
        RECT 88.960 209.250 89.220 209.510 ;
        RECT 79.300 208.910 79.560 209.170 ;
        RECT 26.860 208.570 27.120 208.830 ;
        RECT 30.540 208.570 30.800 208.830 ;
        RECT 33.300 208.570 33.560 208.830 ;
        RECT 38.360 208.570 38.620 208.830 ;
        RECT 45.720 208.570 45.980 208.830 ;
        RECT 61.820 208.570 62.080 208.830 ;
        RECT 75.620 208.570 75.880 208.830 ;
        RECT 82.520 208.570 82.780 208.830 ;
        RECT 83.900 208.570 84.160 208.830 ;
        RECT 122.540 209.590 122.800 209.850 ;
        RECT 124.840 209.590 125.100 209.850 ;
        RECT 111.500 208.910 111.760 209.170 ;
        RECT 105.520 208.570 105.780 208.830 ;
        RECT 111.960 208.570 112.220 208.830 ;
        RECT 112.880 208.570 113.140 208.830 ;
        RECT 123.000 208.570 123.260 208.830 ;
        RECT 130.360 208.570 130.620 208.830 ;
        RECT 27.770 208.060 28.030 208.320 ;
        RECT 28.090 208.060 28.350 208.320 ;
        RECT 28.410 208.060 28.670 208.320 ;
        RECT 28.730 208.060 28.990 208.320 ;
        RECT 29.050 208.060 29.310 208.320 ;
        RECT 62.615 208.060 62.875 208.320 ;
        RECT 62.935 208.060 63.195 208.320 ;
        RECT 63.255 208.060 63.515 208.320 ;
        RECT 63.575 208.060 63.835 208.320 ;
        RECT 63.895 208.060 64.155 208.320 ;
        RECT 97.460 208.060 97.720 208.320 ;
        RECT 97.780 208.060 98.040 208.320 ;
        RECT 98.100 208.060 98.360 208.320 ;
        RECT 98.420 208.060 98.680 208.320 ;
        RECT 98.740 208.060 99.000 208.320 ;
        RECT 132.305 208.060 132.565 208.320 ;
        RECT 132.625 208.060 132.885 208.320 ;
        RECT 132.945 208.060 133.205 208.320 ;
        RECT 133.265 208.060 133.525 208.320 ;
        RECT 133.585 208.060 133.845 208.320 ;
        RECT 21.340 207.550 21.600 207.810 ;
        RECT 31.000 207.550 31.260 207.810 ;
        RECT 47.560 207.550 47.820 207.810 ;
        RECT 55.380 207.550 55.640 207.810 ;
        RECT 61.820 207.550 62.080 207.810 ;
        RECT 26.860 207.210 27.120 207.470 ;
        RECT 26.860 206.530 27.120 206.790 ;
        RECT 32.840 207.210 33.100 207.470 ;
        RECT 47.100 207.210 47.360 207.470 ;
        RECT 38.360 206.530 38.620 206.790 ;
        RECT 39.740 206.530 40.000 206.790 ;
        RECT 52.160 206.530 52.420 206.790 ;
        RECT 74.700 207.550 74.960 207.810 ;
        RECT 83.440 207.550 83.700 207.810 ;
        RECT 100.000 207.550 100.260 207.810 ;
        RECT 92.180 207.210 92.440 207.470 ;
        RECT 64.120 206.870 64.380 207.130 ;
        RECT 44.800 206.190 45.060 206.450 ;
        RECT 70.560 206.530 70.820 206.790 ;
        RECT 84.360 206.870 84.620 207.130 ;
        RECT 72.400 206.530 72.660 206.790 ;
        RECT 82.060 206.530 82.320 206.790 ;
        RECT 84.820 206.530 85.080 206.790 ;
        RECT 91.720 206.530 91.980 206.790 ;
        RECT 99.080 206.530 99.340 206.790 ;
        RECT 110.580 206.530 110.840 206.790 ;
        RECT 112.880 206.530 113.140 206.790 ;
        RECT 29.620 205.850 29.880 206.110 ;
        RECT 30.080 205.850 30.340 206.110 ;
        RECT 45.720 205.850 45.980 206.110 ;
        RECT 65.500 205.850 65.760 206.110 ;
        RECT 68.260 205.850 68.520 206.110 ;
        RECT 71.480 205.850 71.740 206.110 ;
        RECT 77.920 205.850 78.180 206.110 ;
        RECT 83.900 205.850 84.160 206.110 ;
        RECT 93.100 205.850 93.360 206.110 ;
        RECT 99.080 205.850 99.340 206.110 ;
        RECT 105.520 206.190 105.780 206.450 ;
        RECT 108.740 206.190 109.000 206.450 ;
        RECT 122.540 207.550 122.800 207.810 ;
        RECT 124.840 207.550 125.100 207.810 ;
        RECT 130.360 207.550 130.620 207.810 ;
        RECT 127.600 206.530 127.860 206.790 ;
        RECT 127.140 206.190 127.400 206.450 ;
        RECT 137.720 206.190 137.980 206.450 ;
        RECT 110.120 205.850 110.380 206.110 ;
        RECT 129.440 205.850 129.700 206.110 ;
        RECT 45.190 205.340 45.450 205.600 ;
        RECT 45.510 205.340 45.770 205.600 ;
        RECT 45.830 205.340 46.090 205.600 ;
        RECT 46.150 205.340 46.410 205.600 ;
        RECT 46.470 205.340 46.730 205.600 ;
        RECT 80.035 205.340 80.295 205.600 ;
        RECT 80.355 205.340 80.615 205.600 ;
        RECT 80.675 205.340 80.935 205.600 ;
        RECT 80.995 205.340 81.255 205.600 ;
        RECT 81.315 205.340 81.575 205.600 ;
        RECT 114.880 205.340 115.140 205.600 ;
        RECT 115.200 205.340 115.460 205.600 ;
        RECT 115.520 205.340 115.780 205.600 ;
        RECT 115.840 205.340 116.100 205.600 ;
        RECT 116.160 205.340 116.420 205.600 ;
        RECT 149.725 205.340 149.985 205.600 ;
        RECT 150.045 205.340 150.305 205.600 ;
        RECT 150.365 205.340 150.625 205.600 ;
        RECT 150.685 205.340 150.945 205.600 ;
        RECT 151.005 205.340 151.265 205.600 ;
        RECT 33.300 204.830 33.560 205.090 ;
        RECT 38.820 204.830 39.080 205.090 ;
        RECT 44.800 204.830 45.060 205.090 ;
        RECT 46.180 204.830 46.440 205.090 ;
        RECT 47.100 204.830 47.360 205.090 ;
        RECT 42.500 204.150 42.760 204.410 ;
        RECT 31.000 203.810 31.260 204.070 ;
        RECT 37.900 203.810 38.160 204.070 ;
        RECT 41.120 203.810 41.380 204.070 ;
        RECT 46.180 204.150 46.440 204.410 ;
        RECT 47.560 204.150 47.820 204.410 ;
        RECT 58.600 204.150 58.860 204.410 ;
        RECT 40.200 203.470 40.460 203.730 ;
        RECT 30.540 203.130 30.800 203.390 ;
        RECT 64.120 204.830 64.380 205.090 ;
        RECT 68.260 204.830 68.520 205.090 ;
        RECT 72.400 204.830 72.660 205.090 ;
        RECT 79.300 204.830 79.560 205.090 ;
        RECT 82.060 204.830 82.320 205.090 ;
        RECT 84.820 204.830 85.080 205.090 ;
        RECT 93.100 204.830 93.360 205.090 ;
        RECT 69.640 204.150 69.900 204.410 ;
        RECT 70.100 204.150 70.360 204.410 ;
        RECT 71.020 204.150 71.280 204.410 ;
        RECT 71.480 204.150 71.740 204.410 ;
        RECT 66.420 203.470 66.680 203.730 ;
        RECT 67.340 203.470 67.600 203.730 ;
        RECT 77.920 204.490 78.180 204.750 ;
        RECT 73.780 203.470 74.040 203.730 ;
        RECT 78.380 203.130 78.640 203.390 ;
        RECT 82.060 203.810 82.320 204.070 ;
        RECT 88.960 204.150 89.220 204.410 ;
        RECT 91.260 204.150 91.520 204.410 ;
        RECT 112.420 204.150 112.680 204.410 ;
        RECT 84.360 203.810 84.620 204.070 ;
        RECT 92.180 203.130 92.440 203.390 ;
        RECT 92.640 203.130 92.900 203.390 ;
        RECT 106.900 203.470 107.160 203.730 ;
        RECT 99.540 203.130 99.800 203.390 ;
        RECT 110.580 203.130 110.840 203.390 ;
        RECT 27.770 202.620 28.030 202.880 ;
        RECT 28.090 202.620 28.350 202.880 ;
        RECT 28.410 202.620 28.670 202.880 ;
        RECT 28.730 202.620 28.990 202.880 ;
        RECT 29.050 202.620 29.310 202.880 ;
        RECT 62.615 202.620 62.875 202.880 ;
        RECT 62.935 202.620 63.195 202.880 ;
        RECT 63.255 202.620 63.515 202.880 ;
        RECT 63.575 202.620 63.835 202.880 ;
        RECT 63.895 202.620 64.155 202.880 ;
        RECT 97.460 202.620 97.720 202.880 ;
        RECT 97.780 202.620 98.040 202.880 ;
        RECT 98.100 202.620 98.360 202.880 ;
        RECT 98.420 202.620 98.680 202.880 ;
        RECT 98.740 202.620 99.000 202.880 ;
        RECT 132.305 202.620 132.565 202.880 ;
        RECT 132.625 202.620 132.885 202.880 ;
        RECT 132.945 202.620 133.205 202.880 ;
        RECT 133.265 202.620 133.525 202.880 ;
        RECT 133.585 202.620 133.845 202.880 ;
        RECT 15.360 201.090 15.620 201.350 ;
        RECT 19.960 201.090 20.220 201.350 ;
        RECT 20.420 200.750 20.680 201.010 ;
        RECT 38.360 202.110 38.620 202.370 ;
        RECT 41.120 202.110 41.380 202.370 ;
        RECT 48.020 202.110 48.280 202.370 ;
        RECT 31.920 200.750 32.180 201.010 ;
        RECT 39.740 201.090 40.000 201.350 ;
        RECT 42.040 201.770 42.300 202.030 ;
        RECT 43.420 201.770 43.680 202.030 ;
        RECT 65.040 201.770 65.300 202.030 ;
        RECT 71.020 202.110 71.280 202.370 ;
        RECT 73.780 202.110 74.040 202.370 ;
        RECT 77.920 201.770 78.180 202.030 ;
        RECT 48.020 201.090 48.280 201.350 ;
        RECT 51.700 201.090 51.960 201.350 ;
        RECT 42.500 200.750 42.760 201.010 ;
        RECT 47.100 200.750 47.360 201.010 ;
        RECT 69.640 201.090 69.900 201.350 ;
        RECT 24.100 200.410 24.360 200.670 ;
        RECT 38.360 200.410 38.620 200.670 ;
        RECT 40.200 200.410 40.460 200.670 ;
        RECT 52.160 200.410 52.420 200.670 ;
        RECT 67.800 200.410 68.060 200.670 ;
        RECT 82.520 201.430 82.780 201.690 ;
        RECT 91.260 202.110 91.520 202.370 ;
        RECT 112.420 202.110 112.680 202.370 ;
        RECT 71.480 200.750 71.740 201.010 ;
        RECT 71.940 200.750 72.200 201.010 ;
        RECT 78.380 201.090 78.640 201.350 ;
        RECT 82.980 201.090 83.240 201.350 ;
        RECT 99.080 201.770 99.340 202.030 ;
        RECT 100.460 201.090 100.720 201.350 ;
        RECT 108.280 201.090 108.540 201.350 ;
        RECT 110.580 201.430 110.840 201.690 ;
        RECT 110.120 201.090 110.380 201.350 ;
        RECT 123.000 201.090 123.260 201.350 ;
        RECT 127.600 201.090 127.860 201.350 ;
        RECT 84.820 200.410 85.080 200.670 ;
        RECT 117.020 200.750 117.280 201.010 ;
        RECT 101.840 200.410 102.100 200.670 ;
        RECT 121.620 200.410 121.880 200.670 ;
        RECT 45.190 199.900 45.450 200.160 ;
        RECT 45.510 199.900 45.770 200.160 ;
        RECT 45.830 199.900 46.090 200.160 ;
        RECT 46.150 199.900 46.410 200.160 ;
        RECT 46.470 199.900 46.730 200.160 ;
        RECT 80.035 199.900 80.295 200.160 ;
        RECT 80.355 199.900 80.615 200.160 ;
        RECT 80.675 199.900 80.935 200.160 ;
        RECT 80.995 199.900 81.255 200.160 ;
        RECT 81.315 199.900 81.575 200.160 ;
        RECT 114.880 199.900 115.140 200.160 ;
        RECT 115.200 199.900 115.460 200.160 ;
        RECT 115.520 199.900 115.780 200.160 ;
        RECT 115.840 199.900 116.100 200.160 ;
        RECT 116.160 199.900 116.420 200.160 ;
        RECT 149.725 199.900 149.985 200.160 ;
        RECT 150.045 199.900 150.305 200.160 ;
        RECT 150.365 199.900 150.625 200.160 ;
        RECT 150.685 199.900 150.945 200.160 ;
        RECT 151.005 199.900 151.265 200.160 ;
        RECT 20.420 199.390 20.680 199.650 ;
        RECT 24.100 199.390 24.360 199.650 ;
        RECT 26.860 199.390 27.120 199.650 ;
        RECT 30.080 199.390 30.340 199.650 ;
        RECT 25.020 198.710 25.280 198.970 ;
        RECT 31.920 199.390 32.180 199.650 ;
        RECT 48.020 199.390 48.280 199.650 ;
        RECT 51.700 199.390 51.960 199.650 ;
        RECT 52.160 199.390 52.420 199.650 ;
        RECT 53.080 199.390 53.340 199.650 ;
        RECT 69.640 199.390 69.900 199.650 ;
        RECT 32.840 198.710 33.100 198.970 ;
        RECT 35.600 198.710 35.860 198.970 ;
        RECT 27.320 198.370 27.580 198.630 ;
        RECT 41.580 198.370 41.840 198.630 ;
        RECT 49.860 198.710 50.120 198.970 ;
        RECT 66.420 199.050 66.680 199.310 ;
        RECT 78.380 199.050 78.640 199.310 ;
        RECT 80.220 199.390 80.480 199.650 ;
        RECT 82.520 199.390 82.780 199.650 ;
        RECT 84.820 199.390 85.080 199.650 ;
        RECT 100.460 199.390 100.720 199.650 ;
        RECT 117.020 199.390 117.280 199.650 ;
        RECT 77.000 198.710 77.260 198.970 ;
        RECT 51.700 198.370 51.960 198.630 ;
        RECT 71.020 198.370 71.280 198.630 ;
        RECT 92.640 199.050 92.900 199.310 ;
        RECT 92.180 198.710 92.440 198.970 ;
        RECT 100.000 199.050 100.260 199.310 ;
        RECT 101.380 199.050 101.640 199.310 ;
        RECT 106.440 198.710 106.700 198.970 ;
        RECT 127.600 199.050 127.860 199.310 ;
        RECT 30.080 197.690 30.340 197.950 ;
        RECT 35.140 197.690 35.400 197.950 ;
        RECT 35.600 197.690 35.860 197.950 ;
        RECT 56.300 197.690 56.560 197.950 ;
        RECT 71.940 197.690 72.200 197.950 ;
        RECT 73.780 197.690 74.040 197.950 ;
        RECT 81.140 198.370 81.400 198.630 ;
        RECT 82.980 198.370 83.240 198.630 ;
        RECT 101.840 198.370 102.100 198.630 ;
        RECT 115.640 198.710 115.900 198.970 ;
        RECT 129.440 198.710 129.700 198.970 ;
        RECT 78.840 197.690 79.100 197.950 ;
        RECT 94.020 197.690 94.280 197.950 ;
        RECT 99.080 197.690 99.340 197.950 ;
        RECT 124.380 198.370 124.640 198.630 ;
        RECT 108.280 197.690 108.540 197.950 ;
        RECT 113.340 197.690 113.600 197.950 ;
        RECT 123.000 197.690 123.260 197.950 ;
        RECT 27.770 197.180 28.030 197.440 ;
        RECT 28.090 197.180 28.350 197.440 ;
        RECT 28.410 197.180 28.670 197.440 ;
        RECT 28.730 197.180 28.990 197.440 ;
        RECT 29.050 197.180 29.310 197.440 ;
        RECT 62.615 197.180 62.875 197.440 ;
        RECT 62.935 197.180 63.195 197.440 ;
        RECT 63.255 197.180 63.515 197.440 ;
        RECT 63.575 197.180 63.835 197.440 ;
        RECT 63.895 197.180 64.155 197.440 ;
        RECT 97.460 197.180 97.720 197.440 ;
        RECT 97.780 197.180 98.040 197.440 ;
        RECT 98.100 197.180 98.360 197.440 ;
        RECT 98.420 197.180 98.680 197.440 ;
        RECT 98.740 197.180 99.000 197.440 ;
        RECT 132.305 197.180 132.565 197.440 ;
        RECT 132.625 197.180 132.885 197.440 ;
        RECT 132.945 197.180 133.205 197.440 ;
        RECT 133.265 197.180 133.525 197.440 ;
        RECT 133.585 197.180 133.845 197.440 ;
        RECT 27.320 196.330 27.580 196.590 ;
        RECT 41.580 196.670 41.840 196.930 ;
        RECT 43.420 196.670 43.680 196.930 ;
        RECT 57.680 196.670 57.940 196.930 ;
        RECT 67.800 196.670 68.060 196.930 ;
        RECT 71.020 196.670 71.280 196.930 ;
        RECT 79.300 196.670 79.560 196.930 ;
        RECT 82.060 196.670 82.320 196.930 ;
        RECT 100.000 196.670 100.260 196.930 ;
        RECT 104.600 196.670 104.860 196.930 ;
        RECT 106.440 196.670 106.700 196.930 ;
        RECT 115.640 196.670 115.900 196.930 ;
        RECT 121.620 196.670 121.880 196.930 ;
        RECT 66.880 196.330 67.140 196.590 ;
        RECT 70.100 195.990 70.360 196.250 ;
        RECT 82.520 196.330 82.780 196.590 ;
        RECT 37.900 195.310 38.160 195.570 ;
        RECT 44.800 194.970 45.060 195.230 ;
        RECT 55.840 195.650 56.100 195.910 ;
        RECT 56.300 195.650 56.560 195.910 ;
        RECT 63.660 195.650 63.920 195.910 ;
        RECT 71.480 195.650 71.740 195.910 ;
        RECT 71.940 195.650 72.200 195.910 ;
        RECT 77.920 195.650 78.180 195.910 ;
        RECT 78.380 195.650 78.640 195.910 ;
        RECT 61.360 195.310 61.620 195.570 ;
        RECT 62.280 195.310 62.540 195.570 ;
        RECT 78.840 195.310 79.100 195.570 ;
        RECT 81.140 195.310 81.400 195.570 ;
        RECT 88.960 195.990 89.220 196.250 ;
        RECT 112.420 195.990 112.680 196.250 ;
        RECT 118.400 195.990 118.660 196.250 ;
        RECT 60.440 194.970 60.700 195.230 ;
        RECT 63.200 194.970 63.460 195.230 ;
        RECT 66.880 194.970 67.140 195.230 ;
        RECT 79.300 194.970 79.560 195.230 ;
        RECT 99.080 195.310 99.340 195.570 ;
        RECT 100.920 194.970 101.180 195.230 ;
        RECT 102.300 194.970 102.560 195.230 ;
        RECT 117.480 195.650 117.740 195.910 ;
        RECT 104.600 194.970 104.860 195.230 ;
        RECT 106.440 195.310 106.700 195.570 ;
        RECT 105.520 194.970 105.780 195.230 ;
        RECT 111.500 194.970 111.760 195.230 ;
        RECT 113.800 194.970 114.060 195.230 ;
        RECT 121.620 194.970 121.880 195.230 ;
        RECT 45.190 194.460 45.450 194.720 ;
        RECT 45.510 194.460 45.770 194.720 ;
        RECT 45.830 194.460 46.090 194.720 ;
        RECT 46.150 194.460 46.410 194.720 ;
        RECT 46.470 194.460 46.730 194.720 ;
        RECT 80.035 194.460 80.295 194.720 ;
        RECT 80.355 194.460 80.615 194.720 ;
        RECT 80.675 194.460 80.935 194.720 ;
        RECT 80.995 194.460 81.255 194.720 ;
        RECT 81.315 194.460 81.575 194.720 ;
        RECT 114.880 194.460 115.140 194.720 ;
        RECT 115.200 194.460 115.460 194.720 ;
        RECT 115.520 194.460 115.780 194.720 ;
        RECT 115.840 194.460 116.100 194.720 ;
        RECT 116.160 194.460 116.420 194.720 ;
        RECT 149.725 194.460 149.985 194.720 ;
        RECT 150.045 194.460 150.305 194.720 ;
        RECT 150.365 194.460 150.625 194.720 ;
        RECT 150.685 194.460 150.945 194.720 ;
        RECT 151.005 194.460 151.265 194.720 ;
        RECT 14.900 193.270 15.160 193.530 ;
        RECT 15.360 192.930 15.620 193.190 ;
        RECT 19.040 193.270 19.300 193.530 ;
        RECT 25.940 193.270 26.200 193.530 ;
        RECT 26.860 193.270 27.120 193.530 ;
        RECT 35.140 193.950 35.400 194.210 ;
        RECT 47.100 193.950 47.360 194.210 ;
        RECT 51.700 193.950 51.960 194.210 ;
        RECT 54.460 193.950 54.720 194.210 ;
        RECT 60.440 193.950 60.700 194.210 ;
        RECT 61.360 193.950 61.620 194.210 ;
        RECT 62.280 193.950 62.540 194.210 ;
        RECT 35.140 192.930 35.400 193.190 ;
        RECT 37.900 192.930 38.160 193.190 ;
        RECT 40.200 193.270 40.460 193.530 ;
        RECT 13.980 192.250 14.240 192.510 ;
        RECT 29.620 192.250 29.880 192.510 ;
        RECT 39.280 192.590 39.540 192.850 ;
        RECT 47.100 193.270 47.360 193.530 ;
        RECT 64.120 193.950 64.380 194.210 ;
        RECT 73.320 193.950 73.580 194.210 ;
        RECT 77.920 193.950 78.180 194.210 ;
        RECT 78.380 193.950 78.640 194.210 ;
        RECT 34.680 192.250 34.940 192.510 ;
        RECT 35.140 192.250 35.400 192.510 ;
        RECT 37.440 192.250 37.700 192.510 ;
        RECT 38.360 192.250 38.620 192.510 ;
        RECT 38.820 192.250 39.080 192.510 ;
        RECT 40.660 192.250 40.920 192.510 ;
        RECT 44.800 192.590 45.060 192.850 ;
        RECT 66.420 193.270 66.680 193.530 ;
        RECT 63.200 192.930 63.460 193.190 ;
        RECT 63.660 192.930 63.920 193.190 ;
        RECT 64.120 192.930 64.380 193.190 ;
        RECT 67.340 193.270 67.600 193.530 ;
        RECT 73.780 193.270 74.040 193.530 ;
        RECT 79.300 193.950 79.560 194.210 ;
        RECT 86.200 193.950 86.460 194.210 ;
        RECT 47.100 192.250 47.360 192.510 ;
        RECT 53.540 192.250 53.800 192.510 ;
        RECT 56.300 192.590 56.560 192.850 ;
        RECT 57.220 192.250 57.480 192.510 ;
        RECT 61.820 192.250 62.080 192.510 ;
        RECT 68.720 192.930 68.980 193.190 ;
        RECT 72.400 192.930 72.660 193.190 ;
        RECT 78.840 192.930 79.100 193.190 ;
        RECT 66.880 192.590 67.140 192.850 ;
        RECT 67.340 192.250 67.600 192.510 ;
        RECT 77.920 192.250 78.180 192.510 ;
        RECT 81.600 192.250 81.860 192.510 ;
        RECT 88.960 193.270 89.220 193.530 ;
        RECT 98.620 193.270 98.880 193.530 ;
        RECT 100.920 193.270 101.180 193.530 ;
        RECT 101.380 193.270 101.640 193.530 ;
        RECT 102.300 193.950 102.560 194.210 ;
        RECT 120.700 193.950 120.960 194.210 ;
        RECT 121.620 193.950 121.880 194.210 ;
        RECT 110.120 193.270 110.380 193.530 ;
        RECT 116.560 193.270 116.820 193.530 ;
        RECT 102.300 192.930 102.560 193.190 ;
        RECT 106.440 192.930 106.700 193.190 ;
        RECT 111.040 192.930 111.300 193.190 ;
        RECT 113.340 192.590 113.600 192.850 ;
        RECT 117.480 192.590 117.740 192.850 ;
        RECT 121.160 193.270 121.420 193.530 ;
        RECT 124.380 193.270 124.640 193.530 ;
        RECT 119.320 192.930 119.580 193.190 ;
        RECT 93.560 192.250 93.820 192.510 ;
        RECT 96.780 192.250 97.040 192.510 ;
        RECT 100.000 192.250 100.260 192.510 ;
        RECT 100.460 192.250 100.720 192.510 ;
        RECT 120.700 192.250 120.960 192.510 ;
        RECT 123.920 192.590 124.180 192.850 ;
        RECT 126.220 193.270 126.480 193.530 ;
        RECT 130.820 193.270 131.080 193.530 ;
        RECT 127.600 192.930 127.860 193.190 ;
        RECT 124.380 192.250 124.640 192.510 ;
        RECT 129.440 192.250 129.700 192.510 ;
        RECT 131.280 192.250 131.540 192.510 ;
        RECT 27.770 191.740 28.030 192.000 ;
        RECT 28.090 191.740 28.350 192.000 ;
        RECT 28.410 191.740 28.670 192.000 ;
        RECT 28.730 191.740 28.990 192.000 ;
        RECT 29.050 191.740 29.310 192.000 ;
        RECT 62.615 191.740 62.875 192.000 ;
        RECT 62.935 191.740 63.195 192.000 ;
        RECT 63.255 191.740 63.515 192.000 ;
        RECT 63.575 191.740 63.835 192.000 ;
        RECT 63.895 191.740 64.155 192.000 ;
        RECT 97.460 191.740 97.720 192.000 ;
        RECT 97.780 191.740 98.040 192.000 ;
        RECT 98.100 191.740 98.360 192.000 ;
        RECT 98.420 191.740 98.680 192.000 ;
        RECT 98.740 191.740 99.000 192.000 ;
        RECT 132.305 191.740 132.565 192.000 ;
        RECT 132.625 191.740 132.885 192.000 ;
        RECT 132.945 191.740 133.205 192.000 ;
        RECT 133.265 191.740 133.525 192.000 ;
        RECT 133.585 191.740 133.845 192.000 ;
        RECT 19.040 191.230 19.300 191.490 ;
        RECT 26.860 191.230 27.120 191.490 ;
        RECT 29.620 191.230 29.880 191.490 ;
        RECT 32.840 191.230 33.100 191.490 ;
        RECT 37.440 191.230 37.700 191.490 ;
        RECT 38.820 191.230 39.080 191.490 ;
        RECT 44.800 191.230 45.060 191.490 ;
        RECT 53.540 191.230 53.800 191.490 ;
        RECT 54.000 191.230 54.260 191.490 ;
        RECT 65.960 191.230 66.220 191.490 ;
        RECT 71.940 191.230 72.200 191.490 ;
        RECT 78.840 191.230 79.100 191.490 ;
        RECT 86.660 191.230 86.920 191.490 ;
        RECT 88.960 191.230 89.220 191.490 ;
        RECT 108.280 191.230 108.540 191.490 ;
        RECT 111.040 191.230 111.300 191.490 ;
        RECT 126.220 191.230 126.480 191.490 ;
        RECT 129.440 191.230 129.700 191.490 ;
        RECT 130.820 191.230 131.080 191.490 ;
        RECT 54.460 190.890 54.720 191.150 ;
        RECT 86.200 190.890 86.460 191.150 ;
        RECT 92.180 190.890 92.440 191.150 ;
        RECT 96.780 190.890 97.040 191.150 ;
        RECT 13.980 189.870 14.240 190.130 ;
        RECT 15.360 190.210 15.620 190.470 ;
        RECT 22.720 190.210 22.980 190.470 ;
        RECT 29.620 190.210 29.880 190.470 ;
        RECT 26.860 189.870 27.120 190.130 ;
        RECT 34.680 190.210 34.940 190.470 ;
        RECT 40.660 190.210 40.920 190.470 ;
        RECT 53.540 190.210 53.800 190.470 ;
        RECT 57.220 190.550 57.480 190.810 ;
        RECT 73.320 190.550 73.580 190.810 ;
        RECT 77.460 190.550 77.720 190.810 ;
        RECT 54.460 190.210 54.720 190.470 ;
        RECT 55.380 190.210 55.640 190.470 ;
        RECT 14.440 189.530 14.700 189.790 ;
        RECT 20.420 189.530 20.680 189.790 ;
        RECT 26.400 189.530 26.660 189.790 ;
        RECT 47.560 189.870 47.820 190.130 ;
        RECT 73.780 190.210 74.040 190.470 ;
        RECT 72.400 189.870 72.660 190.130 ;
        RECT 73.320 189.870 73.580 190.130 ;
        RECT 92.640 189.870 92.900 190.130 ;
        RECT 94.020 190.210 94.280 190.470 ;
        RECT 102.300 190.550 102.560 190.810 ;
        RECT 112.420 190.550 112.680 190.810 ;
        RECT 116.560 190.550 116.820 190.810 ;
        RECT 103.220 190.210 103.480 190.470 ;
        RECT 113.340 190.210 113.600 190.470 ;
        RECT 117.940 190.210 118.200 190.470 ;
        RECT 120.700 190.550 120.960 190.810 ;
        RECT 95.400 189.870 95.660 190.130 ;
        RECT 97.700 189.870 97.960 190.130 ;
        RECT 120.240 190.210 120.500 190.470 ;
        RECT 124.380 190.210 124.640 190.470 ;
        RECT 125.300 190.210 125.560 190.470 ;
        RECT 52.620 189.530 52.880 189.790 ;
        RECT 53.080 189.530 53.340 189.790 ;
        RECT 56.760 189.530 57.020 189.790 ;
        RECT 66.420 189.530 66.680 189.790 ;
        RECT 69.640 189.530 69.900 189.790 ;
        RECT 71.020 189.530 71.280 189.790 ;
        RECT 76.540 189.530 76.800 189.790 ;
        RECT 79.300 189.530 79.560 189.790 ;
        RECT 99.080 189.530 99.340 189.790 ;
        RECT 121.160 189.530 121.420 189.790 ;
        RECT 121.620 189.530 121.880 189.790 ;
        RECT 130.360 190.210 130.620 190.470 ;
        RECT 131.280 190.210 131.540 190.470 ;
        RECT 45.190 189.020 45.450 189.280 ;
        RECT 45.510 189.020 45.770 189.280 ;
        RECT 45.830 189.020 46.090 189.280 ;
        RECT 46.150 189.020 46.410 189.280 ;
        RECT 46.470 189.020 46.730 189.280 ;
        RECT 80.035 189.020 80.295 189.280 ;
        RECT 80.355 189.020 80.615 189.280 ;
        RECT 80.675 189.020 80.935 189.280 ;
        RECT 80.995 189.020 81.255 189.280 ;
        RECT 81.315 189.020 81.575 189.280 ;
        RECT 114.880 189.020 115.140 189.280 ;
        RECT 115.200 189.020 115.460 189.280 ;
        RECT 115.520 189.020 115.780 189.280 ;
        RECT 115.840 189.020 116.100 189.280 ;
        RECT 116.160 189.020 116.420 189.280 ;
        RECT 149.725 189.020 149.985 189.280 ;
        RECT 150.045 189.020 150.305 189.280 ;
        RECT 150.365 189.020 150.625 189.280 ;
        RECT 150.685 189.020 150.945 189.280 ;
        RECT 151.005 189.020 151.265 189.280 ;
        RECT 14.900 188.510 15.160 188.770 ;
        RECT 17.200 188.170 17.460 188.430 ;
        RECT 19.040 188.170 19.300 188.430 ;
        RECT 20.420 187.490 20.680 187.750 ;
        RECT 24.560 188.170 24.820 188.430 ;
        RECT 25.940 188.510 26.200 188.770 ;
        RECT 55.380 188.510 55.640 188.770 ;
        RECT 31.000 188.170 31.260 188.430 ;
        RECT 52.160 188.170 52.420 188.430 ;
        RECT 53.540 188.170 53.800 188.430 ;
        RECT 30.540 187.830 30.800 188.090 ;
        RECT 31.460 187.830 31.720 188.090 ;
        RECT 35.140 187.830 35.400 188.090 ;
        RECT 41.580 187.830 41.840 188.090 ;
        RECT 47.560 187.830 47.820 188.090 ;
        RECT 51.700 187.830 51.960 188.090 ;
        RECT 42.040 187.490 42.300 187.750 ;
        RECT 49.860 187.490 50.120 187.750 ;
        RECT 56.760 188.170 57.020 188.430 ;
        RECT 55.840 187.830 56.100 188.090 ;
        RECT 61.820 188.510 62.080 188.770 ;
        RECT 65.040 188.510 65.300 188.770 ;
        RECT 67.800 188.510 68.060 188.770 ;
        RECT 73.320 188.510 73.580 188.770 ;
        RECT 77.460 188.510 77.720 188.770 ;
        RECT 78.380 188.510 78.640 188.770 ;
        RECT 78.840 188.510 79.100 188.770 ;
        RECT 67.340 187.830 67.600 188.090 ;
        RECT 69.180 187.830 69.440 188.090 ;
        RECT 69.640 187.830 69.900 188.090 ;
        RECT 70.100 187.830 70.360 188.090 ;
        RECT 71.020 187.830 71.280 188.090 ;
        RECT 65.040 187.490 65.300 187.750 ;
        RECT 66.880 187.490 67.140 187.750 ;
        RECT 72.860 187.830 73.120 188.090 ;
        RECT 73.780 187.830 74.040 188.090 ;
        RECT 75.160 187.830 75.420 188.090 ;
        RECT 83.440 188.170 83.700 188.430 ;
        RECT 84.820 188.170 85.080 188.430 ;
        RECT 86.200 188.170 86.460 188.430 ;
        RECT 97.700 188.510 97.960 188.770 ;
        RECT 113.340 188.510 113.600 188.770 ;
        RECT 116.560 188.510 116.820 188.770 ;
        RECT 82.520 187.830 82.780 188.090 ;
        RECT 22.720 187.150 22.980 187.410 ;
        RECT 16.740 186.810 17.000 187.070 ;
        RECT 27.320 186.810 27.580 187.070 ;
        RECT 31.000 186.810 31.260 187.070 ;
        RECT 53.080 186.810 53.340 187.070 ;
        RECT 58.600 186.810 58.860 187.070 ;
        RECT 61.820 186.810 62.080 187.070 ;
        RECT 66.420 186.810 66.680 187.070 ;
        RECT 71.480 187.150 71.740 187.410 ;
        RECT 74.240 187.150 74.500 187.410 ;
        RECT 82.060 187.490 82.320 187.750 ;
        RECT 78.380 187.150 78.640 187.410 ;
        RECT 92.180 187.830 92.440 188.090 ;
        RECT 92.640 187.830 92.900 188.090 ;
        RECT 94.480 187.830 94.740 188.090 ;
        RECT 94.940 187.830 95.200 188.090 ;
        RECT 100.000 187.830 100.260 188.090 ;
        RECT 100.460 187.830 100.720 188.090 ;
        RECT 101.840 187.830 102.100 188.090 ;
        RECT 102.300 187.830 102.560 188.090 ;
        RECT 102.760 187.830 103.020 188.090 ;
        RECT 103.680 187.830 103.940 188.090 ;
        RECT 117.940 188.170 118.200 188.430 ;
        RECT 98.620 187.490 98.880 187.750 ;
        RECT 76.540 186.810 76.800 187.070 ;
        RECT 77.000 186.810 77.260 187.070 ;
        RECT 80.680 186.810 80.940 187.070 ;
        RECT 117.020 187.150 117.280 187.410 ;
        RECT 83.900 186.810 84.160 187.070 ;
        RECT 87.580 186.810 87.840 187.070 ;
        RECT 92.640 186.810 92.900 187.070 ;
        RECT 96.320 186.810 96.580 187.070 ;
        RECT 99.080 186.810 99.340 187.070 ;
        RECT 103.220 186.810 103.480 187.070 ;
        RECT 104.140 186.810 104.400 187.070 ;
        RECT 117.480 186.810 117.740 187.070 ;
        RECT 27.770 186.300 28.030 186.560 ;
        RECT 28.090 186.300 28.350 186.560 ;
        RECT 28.410 186.300 28.670 186.560 ;
        RECT 28.730 186.300 28.990 186.560 ;
        RECT 29.050 186.300 29.310 186.560 ;
        RECT 62.615 186.300 62.875 186.560 ;
        RECT 62.935 186.300 63.195 186.560 ;
        RECT 63.255 186.300 63.515 186.560 ;
        RECT 63.575 186.300 63.835 186.560 ;
        RECT 63.895 186.300 64.155 186.560 ;
        RECT 97.460 186.300 97.720 186.560 ;
        RECT 97.780 186.300 98.040 186.560 ;
        RECT 98.100 186.300 98.360 186.560 ;
        RECT 98.420 186.300 98.680 186.560 ;
        RECT 98.740 186.300 99.000 186.560 ;
        RECT 132.305 186.300 132.565 186.560 ;
        RECT 132.625 186.300 132.885 186.560 ;
        RECT 132.945 186.300 133.205 186.560 ;
        RECT 133.265 186.300 133.525 186.560 ;
        RECT 133.585 186.300 133.845 186.560 ;
        RECT 17.200 185.790 17.460 186.050 ;
        RECT 19.040 185.790 19.300 186.050 ;
        RECT 24.560 185.790 24.820 186.050 ;
        RECT 26.860 185.790 27.120 186.050 ;
        RECT 27.320 185.790 27.580 186.050 ;
        RECT 31.000 185.790 31.260 186.050 ;
        RECT 20.420 184.770 20.680 185.030 ;
        RECT 25.480 184.770 25.740 185.030 ;
        RECT 38.360 185.790 38.620 186.050 ;
        RECT 39.280 185.790 39.540 186.050 ;
        RECT 42.960 185.790 43.220 186.050 ;
        RECT 53.080 185.790 53.340 186.050 ;
        RECT 57.680 185.790 57.940 186.050 ;
        RECT 60.440 185.790 60.700 186.050 ;
        RECT 65.500 185.790 65.760 186.050 ;
        RECT 67.340 185.790 67.600 186.050 ;
        RECT 67.800 185.790 68.060 186.050 ;
        RECT 69.180 185.790 69.440 186.050 ;
        RECT 71.480 185.790 71.740 186.050 ;
        RECT 41.120 185.450 41.380 185.710 ;
        RECT 26.400 184.430 26.660 184.690 ;
        RECT 25.480 184.090 25.740 184.350 ;
        RECT 30.080 184.430 30.340 184.690 ;
        RECT 32.840 184.770 33.100 185.030 ;
        RECT 35.140 184.770 35.400 185.030 ;
        RECT 40.200 185.110 40.460 185.370 ;
        RECT 40.660 185.110 40.920 185.370 ;
        RECT 66.420 185.450 66.680 185.710 ;
        RECT 48.480 184.770 48.740 185.030 ;
        RECT 52.160 185.110 52.420 185.370 ;
        RECT 42.040 184.430 42.300 184.690 ;
        RECT 47.100 184.430 47.360 184.690 ;
        RECT 49.860 184.430 50.120 184.690 ;
        RECT 56.760 184.770 57.020 185.030 ;
        RECT 61.820 184.770 62.080 185.030 ;
        RECT 71.940 185.110 72.200 185.370 ;
        RECT 76.540 185.450 76.800 185.710 ;
        RECT 78.380 185.450 78.640 185.710 ;
        RECT 90.340 185.790 90.600 186.050 ;
        RECT 103.680 185.790 103.940 186.050 ;
        RECT 84.820 185.450 85.080 185.710 ;
        RECT 31.460 184.090 31.720 184.350 ;
        RECT 37.440 184.090 37.700 184.350 ;
        RECT 38.360 184.090 38.620 184.350 ;
        RECT 52.160 184.090 52.420 184.350 ;
        RECT 53.080 184.090 53.340 184.350 ;
        RECT 72.400 184.770 72.660 185.030 ;
        RECT 66.880 184.430 67.140 184.690 ;
        RECT 71.020 184.090 71.280 184.350 ;
        RECT 75.160 184.430 75.420 184.690 ;
        RECT 103.220 185.450 103.480 185.710 ;
        RECT 112.420 185.790 112.680 186.050 ;
        RECT 120.240 185.790 120.500 186.050 ;
        RECT 105.060 185.450 105.320 185.710 ;
        RECT 109.660 185.450 109.920 185.710 ;
        RECT 87.580 185.110 87.840 185.370 ;
        RECT 99.540 185.110 99.800 185.370 ;
        RECT 104.140 185.110 104.400 185.370 ;
        RECT 111.960 185.450 112.220 185.710 ;
        RECT 114.260 185.450 114.520 185.710 ;
        RECT 79.300 184.770 79.560 185.030 ;
        RECT 82.520 184.770 82.780 185.030 ;
        RECT 80.680 184.430 80.940 184.690 ;
        RECT 72.860 184.090 73.120 184.350 ;
        RECT 103.680 184.770 103.940 185.030 ;
        RECT 99.080 184.430 99.340 184.690 ;
        RECT 90.800 184.090 91.060 184.350 ;
        RECT 111.040 184.770 111.300 185.030 ;
        RECT 109.660 184.430 109.920 184.690 ;
        RECT 113.340 184.770 113.600 185.030 ;
        RECT 119.320 185.110 119.580 185.370 ;
        RECT 121.620 185.110 121.880 185.370 ;
        RECT 124.840 185.110 125.100 185.370 ;
        RECT 127.600 185.110 127.860 185.370 ;
        RECT 121.160 184.770 121.420 185.030 ;
        RECT 125.760 184.770 126.020 185.030 ;
        RECT 123.920 184.430 124.180 184.690 ;
        RECT 129.900 184.430 130.160 184.690 ;
        RECT 111.040 184.090 111.300 184.350 ;
        RECT 116.560 184.090 116.820 184.350 ;
        RECT 118.860 184.090 119.120 184.350 ;
        RECT 119.780 184.090 120.040 184.350 ;
        RECT 126.680 184.090 126.940 184.350 ;
        RECT 134.500 184.090 134.760 184.350 ;
        RECT 45.190 183.580 45.450 183.840 ;
        RECT 45.510 183.580 45.770 183.840 ;
        RECT 45.830 183.580 46.090 183.840 ;
        RECT 46.150 183.580 46.410 183.840 ;
        RECT 46.470 183.580 46.730 183.840 ;
        RECT 80.035 183.580 80.295 183.840 ;
        RECT 80.355 183.580 80.615 183.840 ;
        RECT 80.675 183.580 80.935 183.840 ;
        RECT 80.995 183.580 81.255 183.840 ;
        RECT 81.315 183.580 81.575 183.840 ;
        RECT 114.880 183.580 115.140 183.840 ;
        RECT 115.200 183.580 115.460 183.840 ;
        RECT 115.520 183.580 115.780 183.840 ;
        RECT 115.840 183.580 116.100 183.840 ;
        RECT 116.160 183.580 116.420 183.840 ;
        RECT 149.725 183.580 149.985 183.840 ;
        RECT 150.045 183.580 150.305 183.840 ;
        RECT 150.365 183.580 150.625 183.840 ;
        RECT 150.685 183.580 150.945 183.840 ;
        RECT 151.005 183.580 151.265 183.840 ;
        RECT 32.840 183.070 33.100 183.330 ;
        RECT 37.440 183.070 37.700 183.330 ;
        RECT 40.660 183.070 40.920 183.330 ;
        RECT 53.080 183.070 53.340 183.330 ;
        RECT 30.540 182.730 30.800 182.990 ;
        RECT 35.140 182.730 35.400 182.990 ;
        RECT 15.820 182.390 16.080 182.650 ;
        RECT 17.660 182.390 17.920 182.650 ;
        RECT 25.480 182.050 25.740 182.310 ;
        RECT 42.040 182.390 42.300 182.650 ;
        RECT 50.780 182.390 51.040 182.650 ;
        RECT 56.760 182.730 57.020 182.990 ;
        RECT 61.360 182.730 61.620 182.990 ;
        RECT 56.300 182.390 56.560 182.650 ;
        RECT 60.900 182.390 61.160 182.650 ;
        RECT 63.660 182.390 63.920 182.650 ;
        RECT 69.640 182.730 69.900 182.990 ;
        RECT 75.160 182.730 75.420 182.990 ;
        RECT 76.540 182.730 76.800 182.990 ;
        RECT 88.960 182.730 89.220 182.990 ;
        RECT 94.480 182.730 94.740 182.990 ;
        RECT 82.060 182.390 82.320 182.650 ;
        RECT 40.660 181.710 40.920 181.970 ;
        RECT 17.200 181.370 17.460 181.630 ;
        RECT 18.580 181.370 18.840 181.630 ;
        RECT 20.420 181.370 20.680 181.630 ;
        RECT 41.580 181.370 41.840 181.630 ;
        RECT 49.860 181.370 50.120 181.630 ;
        RECT 70.560 182.050 70.820 182.310 ;
        RECT 71.480 182.050 71.740 182.310 ;
        RECT 83.900 182.050 84.160 182.310 ;
        RECT 90.800 182.050 91.060 182.310 ;
        RECT 58.140 181.710 58.400 181.970 ;
        RECT 64.120 181.710 64.380 181.970 ;
        RECT 68.260 181.710 68.520 181.970 ;
        RECT 102.760 182.730 103.020 182.990 ;
        RECT 106.900 183.070 107.160 183.330 ;
        RECT 113.340 183.070 113.600 183.330 ;
        RECT 121.160 183.070 121.420 183.330 ;
        RECT 117.020 182.730 117.280 182.990 ;
        RECT 105.520 182.390 105.780 182.650 ;
        RECT 102.300 182.050 102.560 182.310 ;
        RECT 109.660 182.390 109.920 182.650 ;
        RECT 111.040 182.390 111.300 182.650 ;
        RECT 118.860 182.730 119.120 182.990 ;
        RECT 119.780 182.730 120.040 182.990 ;
        RECT 126.680 183.070 126.940 183.330 ;
        RECT 129.900 183.070 130.160 183.330 ;
        RECT 121.620 182.390 121.880 182.650 ;
        RECT 123.000 182.390 123.260 182.650 ;
        RECT 113.340 182.050 113.600 182.310 ;
        RECT 110.120 181.710 110.380 181.970 ;
        RECT 116.560 181.710 116.820 181.970 ;
        RECT 120.700 182.050 120.960 182.310 ;
        RECT 125.760 182.390 126.020 182.650 ;
        RECT 126.220 181.710 126.480 181.970 ;
        RECT 51.700 181.370 51.960 181.630 ;
        RECT 53.540 181.370 53.800 181.630 ;
        RECT 54.920 181.370 55.180 181.630 ;
        RECT 57.680 181.370 57.940 181.630 ;
        RECT 65.500 181.370 65.760 181.630 ;
        RECT 83.900 181.370 84.160 181.630 ;
        RECT 91.720 181.370 91.980 181.630 ;
        RECT 96.780 181.370 97.040 181.630 ;
        RECT 109.660 181.370 109.920 181.630 ;
        RECT 117.020 181.370 117.280 181.630 ;
        RECT 123.000 181.370 123.260 181.630 ;
        RECT 27.770 180.860 28.030 181.120 ;
        RECT 28.090 180.860 28.350 181.120 ;
        RECT 28.410 180.860 28.670 181.120 ;
        RECT 28.730 180.860 28.990 181.120 ;
        RECT 29.050 180.860 29.310 181.120 ;
        RECT 62.615 180.860 62.875 181.120 ;
        RECT 62.935 180.860 63.195 181.120 ;
        RECT 63.255 180.860 63.515 181.120 ;
        RECT 63.575 180.860 63.835 181.120 ;
        RECT 63.895 180.860 64.155 181.120 ;
        RECT 97.460 180.860 97.720 181.120 ;
        RECT 97.780 180.860 98.040 181.120 ;
        RECT 98.100 180.860 98.360 181.120 ;
        RECT 98.420 180.860 98.680 181.120 ;
        RECT 98.740 180.860 99.000 181.120 ;
        RECT 132.305 180.860 132.565 181.120 ;
        RECT 132.625 180.860 132.885 181.120 ;
        RECT 132.945 180.860 133.205 181.120 ;
        RECT 133.265 180.860 133.525 181.120 ;
        RECT 133.585 180.860 133.845 181.120 ;
        RECT 20.420 180.350 20.680 180.610 ;
        RECT 42.960 180.350 43.220 180.610 ;
        RECT 13.980 179.330 14.240 179.590 ;
        RECT 17.200 179.330 17.460 179.590 ;
        RECT 34.220 180.010 34.480 180.270 ;
        RECT 35.140 180.010 35.400 180.270 ;
        RECT 36.060 179.670 36.320 179.930 ;
        RECT 22.720 178.650 22.980 178.910 ;
        RECT 23.640 178.990 23.900 179.250 ;
        RECT 35.140 179.330 35.400 179.590 ;
        RECT 43.420 179.330 43.680 179.590 ;
        RECT 43.880 179.330 44.140 179.590 ;
        RECT 49.860 180.350 50.120 180.610 ;
        RECT 54.920 180.350 55.180 180.610 ;
        RECT 56.300 180.350 56.560 180.610 ;
        RECT 78.380 180.350 78.640 180.610 ;
        RECT 48.480 179.670 48.740 179.930 ;
        RECT 47.100 179.330 47.360 179.590 ;
        RECT 25.020 178.650 25.280 178.910 ;
        RECT 37.440 178.990 37.700 179.250 ;
        RECT 32.380 178.650 32.640 178.910 ;
        RECT 42.040 178.650 42.300 178.910 ;
        RECT 50.320 179.330 50.580 179.590 ;
        RECT 51.700 179.330 51.960 179.590 ;
        RECT 54.920 179.670 55.180 179.930 ;
        RECT 53.540 179.330 53.800 179.590 ;
        RECT 57.680 179.670 57.940 179.930 ;
        RECT 58.600 179.330 58.860 179.590 ;
        RECT 60.900 179.330 61.160 179.590 ;
        RECT 56.300 178.650 56.560 178.910 ;
        RECT 59.520 178.990 59.780 179.250 ;
        RECT 59.980 178.650 60.240 178.910 ;
        RECT 67.800 180.010 68.060 180.270 ;
        RECT 68.720 179.670 68.980 179.930 ;
        RECT 86.660 180.350 86.920 180.610 ;
        RECT 87.580 180.350 87.840 180.610 ;
        RECT 94.480 180.350 94.740 180.610 ;
        RECT 102.760 180.350 103.020 180.610 ;
        RECT 113.800 180.350 114.060 180.610 ;
        RECT 122.080 180.350 122.340 180.610 ;
        RECT 122.540 180.350 122.800 180.610 ;
        RECT 71.940 179.330 72.200 179.590 ;
        RECT 67.340 178.650 67.600 178.910 ;
        RECT 78.840 178.990 79.100 179.250 ;
        RECT 83.440 179.330 83.700 179.590 ;
        RECT 82.520 178.990 82.780 179.250 ;
        RECT 119.780 180.010 120.040 180.270 ;
        RECT 96.780 179.670 97.040 179.930 ;
        RECT 89.880 179.330 90.140 179.590 ;
        RECT 87.580 178.650 87.840 178.910 ;
        RECT 94.480 179.330 94.740 179.590 ;
        RECT 96.320 179.330 96.580 179.590 ;
        RECT 98.620 179.330 98.880 179.590 ;
        RECT 111.960 179.670 112.220 179.930 ;
        RECT 103.220 179.330 103.480 179.590 ;
        RECT 105.060 179.330 105.320 179.590 ;
        RECT 92.180 178.650 92.440 178.910 ;
        RECT 110.120 179.330 110.380 179.590 ;
        RECT 106.900 178.990 107.160 179.250 ;
        RECT 108.280 178.990 108.540 179.250 ;
        RECT 113.340 179.330 113.600 179.590 ;
        RECT 121.620 179.670 121.880 179.930 ;
        RECT 123.000 179.670 123.260 179.930 ;
        RECT 116.560 179.330 116.820 179.590 ;
        RECT 119.320 179.330 119.580 179.590 ;
        RECT 129.900 179.670 130.160 179.930 ;
        RECT 134.500 179.330 134.760 179.590 ;
        RECT 105.980 178.650 106.240 178.910 ;
        RECT 109.660 178.650 109.920 178.910 ;
        RECT 117.940 178.650 118.200 178.910 ;
        RECT 123.460 178.650 123.720 178.910 ;
        RECT 127.600 178.650 127.860 178.910 ;
        RECT 45.190 178.140 45.450 178.400 ;
        RECT 45.510 178.140 45.770 178.400 ;
        RECT 45.830 178.140 46.090 178.400 ;
        RECT 46.150 178.140 46.410 178.400 ;
        RECT 46.470 178.140 46.730 178.400 ;
        RECT 80.035 178.140 80.295 178.400 ;
        RECT 80.355 178.140 80.615 178.400 ;
        RECT 80.675 178.140 80.935 178.400 ;
        RECT 80.995 178.140 81.255 178.400 ;
        RECT 81.315 178.140 81.575 178.400 ;
        RECT 114.880 178.140 115.140 178.400 ;
        RECT 115.200 178.140 115.460 178.400 ;
        RECT 115.520 178.140 115.780 178.400 ;
        RECT 115.840 178.140 116.100 178.400 ;
        RECT 116.160 178.140 116.420 178.400 ;
        RECT 149.725 178.140 149.985 178.400 ;
        RECT 150.045 178.140 150.305 178.400 ;
        RECT 150.365 178.140 150.625 178.400 ;
        RECT 150.685 178.140 150.945 178.400 ;
        RECT 151.005 178.140 151.265 178.400 ;
        RECT 17.660 177.630 17.920 177.890 ;
        RECT 23.640 177.630 23.900 177.890 ;
        RECT 34.680 177.630 34.940 177.890 ;
        RECT 36.060 177.630 36.320 177.890 ;
        RECT 55.840 177.630 56.100 177.890 ;
        RECT 57.220 177.630 57.480 177.890 ;
        RECT 59.980 177.630 60.240 177.890 ;
        RECT 16.740 176.950 17.000 177.210 ;
        RECT 18.580 176.950 18.840 177.210 ;
        RECT 22.720 176.950 22.980 177.210 ;
        RECT 32.380 176.950 32.640 177.210 ;
        RECT 33.300 176.950 33.560 177.210 ;
        RECT 56.760 177.290 57.020 177.550 ;
        RECT 71.020 177.630 71.280 177.890 ;
        RECT 76.080 177.630 76.340 177.890 ;
        RECT 65.960 177.290 66.220 177.550 ;
        RECT 68.260 177.290 68.520 177.550 ;
        RECT 15.820 175.930 16.080 176.190 ;
        RECT 33.760 176.610 34.020 176.870 ;
        RECT 35.600 176.950 35.860 177.210 ;
        RECT 39.740 176.950 40.000 177.210 ;
        RECT 49.400 176.950 49.660 177.210 ;
        RECT 59.520 176.950 59.780 177.210 ;
        RECT 77.920 177.290 78.180 177.550 ;
        RECT 36.060 176.610 36.320 176.870 ;
        RECT 57.680 176.610 57.940 176.870 ;
        RECT 58.140 176.610 58.400 176.870 ;
        RECT 58.600 176.610 58.860 176.870 ;
        RECT 25.020 176.270 25.280 176.530 ;
        RECT 38.820 176.270 39.080 176.530 ;
        RECT 66.880 176.610 67.140 176.870 ;
        RECT 68.260 176.610 68.520 176.870 ;
        RECT 72.400 176.950 72.660 177.210 ;
        RECT 64.580 176.270 64.840 176.530 ;
        RECT 26.860 175.930 27.120 176.190 ;
        RECT 36.520 175.930 36.780 176.190 ;
        RECT 38.360 175.930 38.620 176.190 ;
        RECT 79.300 176.950 79.560 177.210 ;
        RECT 82.520 177.630 82.780 177.890 ;
        RECT 87.580 177.630 87.840 177.890 ;
        RECT 90.800 177.630 91.060 177.890 ;
        RECT 83.440 176.950 83.700 177.210 ;
        RECT 94.020 176.950 94.280 177.210 ;
        RECT 96.320 176.950 96.580 177.210 ;
        RECT 96.780 176.950 97.040 177.210 ;
        RECT 103.220 177.630 103.480 177.890 ;
        RECT 112.420 177.630 112.680 177.890 ;
        RECT 122.080 177.630 122.340 177.890 ;
        RECT 127.600 177.630 127.860 177.890 ;
        RECT 105.980 177.290 106.240 177.550 ;
        RECT 108.280 177.290 108.540 177.550 ;
        RECT 117.020 177.290 117.280 177.550 ;
        RECT 92.180 176.610 92.440 176.870 ;
        RECT 103.220 176.610 103.480 176.870 ;
        RECT 106.900 176.950 107.160 177.210 ;
        RECT 105.520 176.610 105.780 176.870 ;
        RECT 108.740 176.950 109.000 177.210 ;
        RECT 109.660 176.950 109.920 177.210 ;
        RECT 117.480 176.950 117.740 177.210 ;
        RECT 122.540 177.290 122.800 177.550 ;
        RECT 123.460 176.950 123.720 177.210 ;
        RECT 120.700 176.270 120.960 176.530 ;
        RECT 130.360 176.270 130.620 176.530 ;
        RECT 78.840 175.930 79.100 176.190 ;
        RECT 82.060 175.930 82.320 176.190 ;
        RECT 94.480 175.930 94.740 176.190 ;
        RECT 104.600 175.930 104.860 176.190 ;
        RECT 108.740 175.930 109.000 176.190 ;
        RECT 112.880 175.930 113.140 176.190 ;
        RECT 119.320 175.930 119.580 176.190 ;
        RECT 125.300 175.930 125.560 176.190 ;
        RECT 27.770 175.420 28.030 175.680 ;
        RECT 28.090 175.420 28.350 175.680 ;
        RECT 28.410 175.420 28.670 175.680 ;
        RECT 28.730 175.420 28.990 175.680 ;
        RECT 29.050 175.420 29.310 175.680 ;
        RECT 62.615 175.420 62.875 175.680 ;
        RECT 62.935 175.420 63.195 175.680 ;
        RECT 63.255 175.420 63.515 175.680 ;
        RECT 63.575 175.420 63.835 175.680 ;
        RECT 63.895 175.420 64.155 175.680 ;
        RECT 97.460 175.420 97.720 175.680 ;
        RECT 97.780 175.420 98.040 175.680 ;
        RECT 98.100 175.420 98.360 175.680 ;
        RECT 98.420 175.420 98.680 175.680 ;
        RECT 98.740 175.420 99.000 175.680 ;
        RECT 132.305 175.420 132.565 175.680 ;
        RECT 132.625 175.420 132.885 175.680 ;
        RECT 132.945 175.420 133.205 175.680 ;
        RECT 133.265 175.420 133.525 175.680 ;
        RECT 133.585 175.420 133.845 175.680 ;
        RECT 37.440 174.910 37.700 175.170 ;
        RECT 42.500 174.910 42.760 175.170 ;
        RECT 58.140 174.910 58.400 175.170 ;
        RECT 63.660 174.910 63.920 175.170 ;
        RECT 72.400 174.910 72.660 175.170 ;
        RECT 89.880 174.910 90.140 175.170 ;
        RECT 90.340 174.910 90.600 175.170 ;
        RECT 105.060 174.910 105.320 175.170 ;
        RECT 105.980 174.910 106.240 175.170 ;
        RECT 112.880 174.910 113.140 175.170 ;
        RECT 114.260 174.910 114.520 175.170 ;
        RECT 117.480 174.910 117.740 175.170 ;
        RECT 119.320 174.910 119.580 175.170 ;
        RECT 125.300 174.910 125.560 175.170 ;
        RECT 42.040 174.570 42.300 174.830 ;
        RECT 38.820 174.230 39.080 174.490 ;
        RECT 44.340 174.230 44.600 174.490 ;
        RECT 44.800 174.230 45.060 174.490 ;
        RECT 50.320 174.230 50.580 174.490 ;
        RECT 50.780 174.230 51.040 174.490 ;
        RECT 71.940 174.570 72.200 174.830 ;
        RECT 18.120 173.890 18.380 174.150 ;
        RECT 36.520 173.890 36.780 174.150 ;
        RECT 38.360 173.890 38.620 174.150 ;
        RECT 42.960 173.890 43.220 174.150 ;
        RECT 43.880 173.890 44.140 174.150 ;
        RECT 56.300 174.230 56.560 174.490 ;
        RECT 35.140 173.550 35.400 173.810 ;
        RECT 36.980 173.550 37.240 173.810 ;
        RECT 42.040 173.550 42.300 173.810 ;
        RECT 54.920 173.890 55.180 174.150 ;
        RECT 64.580 173.890 64.840 174.150 ;
        RECT 71.480 174.230 71.740 174.490 ;
        RECT 68.260 173.890 68.520 174.150 ;
        RECT 73.320 173.890 73.580 174.150 ;
        RECT 78.380 174.230 78.640 174.490 ;
        RECT 82.060 174.230 82.320 174.490 ;
        RECT 85.280 174.230 85.540 174.490 ;
        RECT 74.240 173.890 74.500 174.150 ;
        RECT 76.540 173.890 76.800 174.150 ;
        RECT 65.500 173.550 65.760 173.810 ;
        RECT 16.280 173.210 16.540 173.470 ;
        RECT 33.300 173.210 33.560 173.470 ;
        RECT 38.820 173.210 39.080 173.470 ;
        RECT 43.420 173.210 43.680 173.470 ;
        RECT 44.340 173.210 44.600 173.470 ;
        RECT 65.040 173.210 65.300 173.470 ;
        RECT 69.180 173.550 69.440 173.810 ;
        RECT 92.180 174.230 92.440 174.490 ;
        RECT 93.100 174.230 93.360 174.490 ;
        RECT 94.020 174.230 94.280 174.490 ;
        RECT 91.260 173.890 91.520 174.150 ;
        RECT 103.220 173.550 103.480 173.810 ;
        RECT 111.040 173.890 111.300 174.150 ;
        RECT 113.340 173.890 113.600 174.150 ;
        RECT 117.020 173.890 117.280 174.150 ;
        RECT 118.860 173.890 119.120 174.150 ;
        RECT 120.700 173.890 120.960 174.150 ;
        RECT 125.760 173.890 126.020 174.150 ;
        RECT 70.100 173.210 70.360 173.470 ;
        RECT 72.860 173.210 73.120 173.470 ;
        RECT 74.240 173.210 74.500 173.470 ;
        RECT 82.520 173.210 82.780 173.470 ;
        RECT 94.480 173.210 94.740 173.470 ;
        RECT 99.080 173.210 99.340 173.470 ;
        RECT 116.560 173.210 116.820 173.470 ;
        RECT 122.540 173.210 122.800 173.470 ;
        RECT 45.190 172.700 45.450 172.960 ;
        RECT 45.510 172.700 45.770 172.960 ;
        RECT 45.830 172.700 46.090 172.960 ;
        RECT 46.150 172.700 46.410 172.960 ;
        RECT 46.470 172.700 46.730 172.960 ;
        RECT 80.035 172.700 80.295 172.960 ;
        RECT 80.355 172.700 80.615 172.960 ;
        RECT 80.675 172.700 80.935 172.960 ;
        RECT 80.995 172.700 81.255 172.960 ;
        RECT 81.315 172.700 81.575 172.960 ;
        RECT 114.880 172.700 115.140 172.960 ;
        RECT 115.200 172.700 115.460 172.960 ;
        RECT 115.520 172.700 115.780 172.960 ;
        RECT 115.840 172.700 116.100 172.960 ;
        RECT 116.160 172.700 116.420 172.960 ;
        RECT 149.725 172.700 149.985 172.960 ;
        RECT 150.045 172.700 150.305 172.960 ;
        RECT 150.365 172.700 150.625 172.960 ;
        RECT 150.685 172.700 150.945 172.960 ;
        RECT 151.005 172.700 151.265 172.960 ;
        RECT 16.280 171.850 16.540 172.110 ;
        RECT 13.980 171.510 14.240 171.770 ;
        RECT 15.820 170.490 16.080 170.750 ;
        RECT 22.720 170.490 22.980 170.750 ;
        RECT 26.400 171.850 26.660 172.110 ;
        RECT 43.420 172.190 43.680 172.450 ;
        RECT 32.380 171.510 32.640 171.770 ;
        RECT 33.300 171.170 33.560 171.430 ;
        RECT 33.760 171.170 34.020 171.430 ;
        RECT 36.980 171.170 37.240 171.430 ;
        RECT 39.280 171.510 39.540 171.770 ;
        RECT 42.040 171.510 42.300 171.770 ;
        RECT 42.960 171.510 43.220 171.770 ;
        RECT 45.260 171.850 45.520 172.110 ;
        RECT 53.540 172.190 53.800 172.450 ;
        RECT 54.920 172.190 55.180 172.450 ;
        RECT 65.040 172.190 65.300 172.450 ;
        RECT 68.260 172.190 68.520 172.450 ;
        RECT 73.320 172.190 73.580 172.450 ;
        RECT 74.700 172.190 74.960 172.450 ;
        RECT 76.080 172.190 76.340 172.450 ;
        RECT 76.540 172.190 76.800 172.450 ;
        RECT 82.060 172.190 82.320 172.450 ;
        RECT 82.980 172.190 83.240 172.450 ;
        RECT 85.280 172.190 85.540 172.450 ;
        RECT 90.340 172.190 90.600 172.450 ;
        RECT 92.180 172.190 92.440 172.450 ;
        RECT 94.480 172.190 94.740 172.450 ;
        RECT 113.340 172.190 113.600 172.450 ;
        RECT 51.240 171.850 51.500 172.110 ;
        RECT 48.940 171.510 49.200 171.770 ;
        RECT 44.800 171.170 45.060 171.430 ;
        RECT 57.220 171.510 57.480 171.770 ;
        RECT 58.140 171.510 58.400 171.770 ;
        RECT 72.400 171.510 72.660 171.770 ;
        RECT 88.960 171.850 89.220 172.110 ;
        RECT 118.860 172.190 119.120 172.450 ;
        RECT 123.460 172.190 123.720 172.450 ;
        RECT 129.900 172.190 130.160 172.450 ;
        RECT 74.240 171.510 74.500 171.770 ;
        RECT 77.460 171.510 77.720 171.770 ;
        RECT 77.920 171.510 78.180 171.770 ;
        RECT 79.300 171.510 79.560 171.770 ;
        RECT 27.320 170.830 27.580 171.090 ;
        RECT 30.540 170.490 30.800 170.750 ;
        RECT 31.000 170.490 31.260 170.750 ;
        RECT 36.060 170.490 36.320 170.750 ;
        RECT 40.660 170.490 40.920 170.750 ;
        RECT 41.580 170.490 41.840 170.750 ;
        RECT 48.480 170.490 48.740 170.750 ;
        RECT 59.520 170.490 59.780 170.750 ;
        RECT 59.980 170.490 60.240 170.750 ;
        RECT 72.860 171.170 73.120 171.430 ;
        RECT 76.540 171.170 76.800 171.430 ;
        RECT 75.620 170.830 75.880 171.090 ;
        RECT 64.580 170.490 64.840 170.750 ;
        RECT 71.020 170.490 71.280 170.750 ;
        RECT 73.320 170.490 73.580 170.750 ;
        RECT 74.700 170.490 74.960 170.750 ;
        RECT 76.540 170.490 76.800 170.750 ;
        RECT 105.060 171.170 105.320 171.430 ;
        RECT 108.740 171.170 109.000 171.430 ;
        RECT 114.260 171.510 114.520 171.770 ;
        RECT 116.560 171.510 116.820 171.770 ;
        RECT 117.940 171.850 118.200 172.110 ;
        RECT 119.780 171.510 120.040 171.770 ;
        RECT 124.380 171.510 124.640 171.770 ;
        RECT 123.000 171.170 123.260 171.430 ;
        RECT 99.540 170.490 99.800 170.750 ;
        RECT 102.760 170.490 103.020 170.750 ;
        RECT 114.720 170.490 114.980 170.750 ;
        RECT 27.770 169.980 28.030 170.240 ;
        RECT 28.090 169.980 28.350 170.240 ;
        RECT 28.410 169.980 28.670 170.240 ;
        RECT 28.730 169.980 28.990 170.240 ;
        RECT 29.050 169.980 29.310 170.240 ;
        RECT 62.615 169.980 62.875 170.240 ;
        RECT 62.935 169.980 63.195 170.240 ;
        RECT 63.255 169.980 63.515 170.240 ;
        RECT 63.575 169.980 63.835 170.240 ;
        RECT 63.895 169.980 64.155 170.240 ;
        RECT 97.460 169.980 97.720 170.240 ;
        RECT 97.780 169.980 98.040 170.240 ;
        RECT 98.100 169.980 98.360 170.240 ;
        RECT 98.420 169.980 98.680 170.240 ;
        RECT 98.740 169.980 99.000 170.240 ;
        RECT 132.305 169.980 132.565 170.240 ;
        RECT 132.625 169.980 132.885 170.240 ;
        RECT 132.945 169.980 133.205 170.240 ;
        RECT 133.265 169.980 133.525 170.240 ;
        RECT 133.585 169.980 133.845 170.240 ;
        RECT 16.740 169.470 17.000 169.730 ;
        RECT 18.120 169.470 18.380 169.730 ;
        RECT 26.860 169.470 27.120 169.730 ;
        RECT 30.540 169.470 30.800 169.730 ;
        RECT 36.980 169.470 37.240 169.730 ;
        RECT 15.820 169.130 16.080 169.390 ;
        RECT 26.400 168.790 26.660 169.050 ;
        RECT 22.720 168.110 22.980 168.370 ;
        RECT 27.320 168.450 27.580 168.710 ;
        RECT 19.040 167.770 19.300 168.030 ;
        RECT 28.240 168.450 28.500 168.710 ;
        RECT 35.600 168.450 35.860 168.710 ;
        RECT 40.660 169.470 40.920 169.730 ;
        RECT 42.960 169.470 43.220 169.730 ;
        RECT 48.940 169.470 49.200 169.730 ;
        RECT 49.400 169.470 49.660 169.730 ;
        RECT 45.260 169.130 45.520 169.390 ;
        RECT 93.100 169.470 93.360 169.730 ;
        RECT 108.740 169.470 109.000 169.730 ;
        RECT 114.720 169.470 114.980 169.730 ;
        RECT 118.860 169.470 119.120 169.730 ;
        RECT 124.380 169.470 124.640 169.730 ;
        RECT 39.280 168.790 39.540 169.050 ;
        RECT 48.480 168.790 48.740 169.050 ;
        RECT 42.500 168.450 42.760 168.710 ;
        RECT 32.840 168.110 33.100 168.370 ;
        RECT 33.760 168.110 34.020 168.370 ;
        RECT 56.300 169.130 56.560 169.390 ;
        RECT 58.140 169.130 58.400 169.390 ;
        RECT 58.600 169.130 58.860 169.390 ;
        RECT 74.240 169.130 74.500 169.390 ;
        RECT 77.000 169.130 77.260 169.390 ;
        RECT 95.400 169.130 95.660 169.390 ;
        RECT 111.960 169.130 112.220 169.390 ;
        RECT 64.580 168.790 64.840 169.050 ;
        RECT 57.220 168.450 57.480 168.710 ;
        RECT 58.140 168.450 58.400 168.710 ;
        RECT 72.400 168.790 72.660 169.050 ;
        RECT 76.080 168.790 76.340 169.050 ;
        RECT 85.280 168.450 85.540 168.710 ;
        RECT 95.400 168.450 95.660 168.710 ;
        RECT 96.780 168.450 97.040 168.710 ;
        RECT 98.160 168.450 98.420 168.710 ;
        RECT 98.620 168.450 98.880 168.710 ;
        RECT 99.540 168.450 99.800 168.710 ;
        RECT 100.000 168.450 100.260 168.710 ;
        RECT 100.920 168.790 101.180 169.050 ;
        RECT 109.200 168.790 109.460 169.050 ;
        RECT 68.260 168.110 68.520 168.370 ;
        RECT 83.440 168.110 83.700 168.370 ;
        RECT 113.340 168.450 113.600 168.710 ;
        RECT 116.100 168.450 116.360 168.710 ;
        RECT 118.860 168.450 119.120 168.710 ;
        RECT 119.780 168.450 120.040 168.710 ;
        RECT 121.160 168.450 121.420 168.710 ;
        RECT 122.540 168.450 122.800 168.710 ;
        RECT 38.820 167.770 39.080 168.030 ;
        RECT 41.580 167.770 41.840 168.030 ;
        RECT 50.320 167.770 50.580 168.030 ;
        RECT 51.700 167.770 51.960 168.030 ;
        RECT 53.540 167.770 53.800 168.030 ;
        RECT 63.200 167.770 63.460 168.030 ;
        RECT 75.160 167.770 75.420 168.030 ;
        RECT 78.380 167.770 78.640 168.030 ;
        RECT 91.260 167.770 91.520 168.030 ;
        RECT 117.940 168.110 118.200 168.370 ;
        RECT 110.580 167.770 110.840 168.030 ;
        RECT 114.260 167.770 114.520 168.030 ;
        RECT 116.560 167.770 116.820 168.030 ;
        RECT 45.190 167.260 45.450 167.520 ;
        RECT 45.510 167.260 45.770 167.520 ;
        RECT 45.830 167.260 46.090 167.520 ;
        RECT 46.150 167.260 46.410 167.520 ;
        RECT 46.470 167.260 46.730 167.520 ;
        RECT 80.035 167.260 80.295 167.520 ;
        RECT 80.355 167.260 80.615 167.520 ;
        RECT 80.675 167.260 80.935 167.520 ;
        RECT 80.995 167.260 81.255 167.520 ;
        RECT 81.315 167.260 81.575 167.520 ;
        RECT 114.880 167.260 115.140 167.520 ;
        RECT 115.200 167.260 115.460 167.520 ;
        RECT 115.520 167.260 115.780 167.520 ;
        RECT 115.840 167.260 116.100 167.520 ;
        RECT 116.160 167.260 116.420 167.520 ;
        RECT 149.725 167.260 149.985 167.520 ;
        RECT 150.045 167.260 150.305 167.520 ;
        RECT 150.365 167.260 150.625 167.520 ;
        RECT 150.685 167.260 150.945 167.520 ;
        RECT 151.005 167.260 151.265 167.520 ;
        RECT 28.240 166.750 28.500 167.010 ;
        RECT 31.000 166.750 31.260 167.010 ;
        RECT 32.840 166.750 33.100 167.010 ;
        RECT 35.600 166.750 35.860 167.010 ;
        RECT 52.160 166.750 52.420 167.010 ;
        RECT 67.340 166.750 67.600 167.010 ;
        RECT 68.260 166.750 68.520 167.010 ;
        RECT 73.320 166.750 73.580 167.010 ;
        RECT 26.400 166.070 26.660 166.330 ;
        RECT 53.540 166.410 53.800 166.670 ;
        RECT 74.240 166.410 74.500 166.670 ;
        RECT 75.160 166.410 75.420 166.670 ;
        RECT 42.040 166.070 42.300 166.330 ;
        RECT 51.700 166.070 51.960 166.330 ;
        RECT 43.880 165.730 44.140 165.990 ;
        RECT 56.300 166.070 56.560 166.330 ;
        RECT 63.200 166.070 63.460 166.330 ;
        RECT 69.180 166.070 69.440 166.330 ;
        RECT 73.320 166.070 73.580 166.330 ;
        RECT 79.300 166.750 79.560 167.010 ;
        RECT 74.700 165.730 74.960 165.990 ;
        RECT 75.160 165.730 75.420 165.990 ;
        RECT 82.520 166.070 82.780 166.330 ;
        RECT 31.920 165.390 32.180 165.650 ;
        RECT 52.620 165.390 52.880 165.650 ;
        RECT 53.080 165.390 53.340 165.650 ;
        RECT 76.080 165.390 76.340 165.650 ;
        RECT 98.160 166.750 98.420 167.010 ;
        RECT 98.620 166.750 98.880 167.010 ;
        RECT 102.760 166.750 103.020 167.010 ;
        RECT 95.400 166.410 95.660 166.670 ;
        RECT 100.000 166.410 100.260 166.670 ;
        RECT 116.560 166.750 116.820 167.010 ;
        RECT 112.420 166.410 112.680 166.670 ;
        RECT 92.640 166.070 92.900 166.330 ;
        RECT 95.860 166.070 96.120 166.330 ;
        RECT 96.320 166.070 96.580 166.330 ;
        RECT 104.600 166.070 104.860 166.330 ;
        RECT 111.040 166.070 111.300 166.330 ;
        RECT 124.840 166.410 125.100 166.670 ;
        RECT 110.580 165.730 110.840 165.990 ;
        RECT 111.960 165.730 112.220 165.990 ;
        RECT 127.140 166.070 127.400 166.330 ;
        RECT 117.940 165.730 118.200 165.990 ;
        RECT 111.040 165.390 111.300 165.650 ;
        RECT 32.840 165.050 33.100 165.310 ;
        RECT 35.600 165.050 35.860 165.310 ;
        RECT 43.420 165.050 43.680 165.310 ;
        RECT 52.160 165.050 52.420 165.310 ;
        RECT 71.480 165.050 71.740 165.310 ;
        RECT 77.460 165.050 77.720 165.310 ;
        RECT 95.400 165.050 95.660 165.310 ;
        RECT 107.820 165.050 108.080 165.310 ;
        RECT 119.320 165.050 119.580 165.310 ;
        RECT 121.160 165.050 121.420 165.310 ;
        RECT 27.770 164.540 28.030 164.800 ;
        RECT 28.090 164.540 28.350 164.800 ;
        RECT 28.410 164.540 28.670 164.800 ;
        RECT 28.730 164.540 28.990 164.800 ;
        RECT 29.050 164.540 29.310 164.800 ;
        RECT 62.615 164.540 62.875 164.800 ;
        RECT 62.935 164.540 63.195 164.800 ;
        RECT 63.255 164.540 63.515 164.800 ;
        RECT 63.575 164.540 63.835 164.800 ;
        RECT 63.895 164.540 64.155 164.800 ;
        RECT 97.460 164.540 97.720 164.800 ;
        RECT 97.780 164.540 98.040 164.800 ;
        RECT 98.100 164.540 98.360 164.800 ;
        RECT 98.420 164.540 98.680 164.800 ;
        RECT 98.740 164.540 99.000 164.800 ;
        RECT 132.305 164.540 132.565 164.800 ;
        RECT 132.625 164.540 132.885 164.800 ;
        RECT 132.945 164.540 133.205 164.800 ;
        RECT 133.265 164.540 133.525 164.800 ;
        RECT 133.585 164.540 133.845 164.800 ;
        RECT 26.400 164.030 26.660 164.290 ;
        RECT 16.280 163.010 16.540 163.270 ;
        RECT 19.040 163.010 19.300 163.270 ;
        RECT 37.900 164.030 38.160 164.290 ;
        RECT 51.700 164.030 51.960 164.290 ;
        RECT 30.540 163.350 30.800 163.610 ;
        RECT 31.460 163.350 31.720 163.610 ;
        RECT 33.760 163.010 34.020 163.270 ;
        RECT 39.740 163.010 40.000 163.270 ;
        RECT 41.120 163.010 41.380 163.270 ;
        RECT 43.420 163.010 43.680 163.270 ;
        RECT 37.440 162.670 37.700 162.930 ;
        RECT 50.320 163.350 50.580 163.610 ;
        RECT 53.540 164.030 53.800 164.290 ;
        RECT 65.960 164.030 66.220 164.290 ;
        RECT 69.180 164.030 69.440 164.290 ;
        RECT 74.240 164.030 74.500 164.290 ;
        RECT 75.160 164.030 75.420 164.290 ;
        RECT 77.920 164.030 78.180 164.290 ;
        RECT 96.320 164.030 96.580 164.290 ;
        RECT 107.820 164.030 108.080 164.290 ;
        RECT 95.860 163.690 96.120 163.950 ;
        RECT 52.620 163.010 52.880 163.270 ;
        RECT 78.380 163.350 78.640 163.610 ;
        RECT 92.180 163.350 92.440 163.610 ;
        RECT 56.300 163.010 56.560 163.270 ;
        RECT 56.760 163.010 57.020 163.270 ;
        RECT 70.560 163.010 70.820 163.270 ;
        RECT 38.360 162.330 38.620 162.590 ;
        RECT 43.420 162.330 43.680 162.590 ;
        RECT 50.780 162.330 51.040 162.590 ;
        RECT 53.080 162.330 53.340 162.590 ;
        RECT 71.480 162.670 71.740 162.930 ;
        RECT 71.940 162.670 72.200 162.930 ;
        RECT 72.860 162.670 73.120 162.930 ;
        RECT 77.000 163.010 77.260 163.270 ;
        RECT 93.560 163.010 93.820 163.270 ;
        RECT 57.680 162.330 57.940 162.590 ;
        RECT 90.800 162.670 91.060 162.930 ;
        RECT 99.080 163.010 99.340 163.270 ;
        RECT 100.000 162.670 100.260 162.930 ;
        RECT 82.520 162.330 82.780 162.590 ;
        RECT 85.280 162.330 85.540 162.590 ;
        RECT 106.440 162.330 106.700 162.590 ;
        RECT 45.190 161.820 45.450 162.080 ;
        RECT 45.510 161.820 45.770 162.080 ;
        RECT 45.830 161.820 46.090 162.080 ;
        RECT 46.150 161.820 46.410 162.080 ;
        RECT 46.470 161.820 46.730 162.080 ;
        RECT 80.035 161.820 80.295 162.080 ;
        RECT 80.355 161.820 80.615 162.080 ;
        RECT 80.675 161.820 80.935 162.080 ;
        RECT 80.995 161.820 81.255 162.080 ;
        RECT 81.315 161.820 81.575 162.080 ;
        RECT 114.880 161.820 115.140 162.080 ;
        RECT 115.200 161.820 115.460 162.080 ;
        RECT 115.520 161.820 115.780 162.080 ;
        RECT 115.840 161.820 116.100 162.080 ;
        RECT 116.160 161.820 116.420 162.080 ;
        RECT 149.725 161.820 149.985 162.080 ;
        RECT 150.045 161.820 150.305 162.080 ;
        RECT 150.365 161.820 150.625 162.080 ;
        RECT 150.685 161.820 150.945 162.080 ;
        RECT 151.005 161.820 151.265 162.080 ;
        RECT 43.420 161.310 43.680 161.570 ;
        RECT 56.760 161.310 57.020 161.570 ;
        RECT 75.160 161.310 75.420 161.570 ;
        RECT 77.000 161.310 77.260 161.570 ;
        RECT 74.700 160.970 74.960 161.230 ;
        RECT 26.860 160.630 27.120 160.890 ;
        RECT 37.440 160.630 37.700 160.890 ;
        RECT 38.820 160.630 39.080 160.890 ;
        RECT 41.120 160.630 41.380 160.890 ;
        RECT 44.800 160.630 45.060 160.890 ;
        RECT 49.860 160.630 50.120 160.890 ;
        RECT 50.780 160.630 51.040 160.890 ;
        RECT 58.600 160.630 58.860 160.890 ;
        RECT 16.280 160.290 16.540 160.550 ;
        RECT 64.580 160.290 64.840 160.550 ;
        RECT 52.620 159.950 52.880 160.210 ;
        RECT 56.300 159.950 56.560 160.210 ;
        RECT 71.480 160.630 71.740 160.890 ;
        RECT 75.160 160.630 75.420 160.890 ;
        RECT 77.000 160.630 77.260 160.890 ;
        RECT 70.560 160.290 70.820 160.550 ;
        RECT 74.240 160.290 74.500 160.550 ;
        RECT 31.460 159.610 31.720 159.870 ;
        RECT 39.740 159.610 40.000 159.870 ;
        RECT 52.160 159.610 52.420 159.870 ;
        RECT 65.960 159.610 66.220 159.870 ;
        RECT 71.940 159.610 72.200 159.870 ;
        RECT 76.080 160.290 76.340 160.550 ;
        RECT 76.540 160.290 76.800 160.550 ;
        RECT 81.140 160.290 81.400 160.550 ;
        RECT 81.600 160.290 81.860 160.550 ;
        RECT 82.520 160.630 82.780 160.890 ;
        RECT 83.440 160.630 83.700 160.890 ;
        RECT 83.900 160.630 84.160 160.890 ;
        RECT 101.840 161.310 102.100 161.570 ;
        RECT 106.440 161.310 106.700 161.570 ;
        RECT 111.960 161.310 112.220 161.570 ;
        RECT 92.180 160.630 92.440 160.890 ;
        RECT 96.780 160.630 97.040 160.890 ;
        RECT 86.660 160.290 86.920 160.550 ;
        RECT 90.800 160.290 91.060 160.550 ;
        RECT 93.560 160.290 93.820 160.550 ;
        RECT 78.380 159.610 78.640 159.870 ;
        RECT 80.680 159.950 80.940 160.210 ;
        RECT 81.140 159.610 81.400 159.870 ;
        RECT 81.600 159.610 81.860 159.870 ;
        RECT 93.100 159.610 93.360 159.870 ;
        RECT 27.770 159.100 28.030 159.360 ;
        RECT 28.090 159.100 28.350 159.360 ;
        RECT 28.410 159.100 28.670 159.360 ;
        RECT 28.730 159.100 28.990 159.360 ;
        RECT 29.050 159.100 29.310 159.360 ;
        RECT 62.615 159.100 62.875 159.360 ;
        RECT 62.935 159.100 63.195 159.360 ;
        RECT 63.255 159.100 63.515 159.360 ;
        RECT 63.575 159.100 63.835 159.360 ;
        RECT 63.895 159.100 64.155 159.360 ;
        RECT 97.460 159.100 97.720 159.360 ;
        RECT 97.780 159.100 98.040 159.360 ;
        RECT 98.100 159.100 98.360 159.360 ;
        RECT 98.420 159.100 98.680 159.360 ;
        RECT 98.740 159.100 99.000 159.360 ;
        RECT 132.305 159.100 132.565 159.360 ;
        RECT 132.625 159.100 132.885 159.360 ;
        RECT 132.945 159.100 133.205 159.360 ;
        RECT 133.265 159.100 133.525 159.360 ;
        RECT 133.585 159.100 133.845 159.360 ;
        RECT 26.860 158.590 27.120 158.850 ;
        RECT 53.080 158.590 53.340 158.850 ;
        RECT 57.680 158.590 57.940 158.850 ;
        RECT 58.600 158.590 58.860 158.850 ;
        RECT 70.560 158.590 70.820 158.850 ;
        RECT 72.860 158.590 73.120 158.850 ;
        RECT 75.620 158.590 75.880 158.850 ;
        RECT 78.380 158.590 78.640 158.850 ;
        RECT 84.820 158.590 85.080 158.850 ;
        RECT 93.560 158.590 93.820 158.850 ;
        RECT 75.160 157.910 75.420 158.170 ;
        RECT 25.020 157.570 25.280 157.830 ;
        RECT 25.480 157.570 25.740 157.830 ;
        RECT 71.940 157.570 72.200 157.830 ;
        RECT 42.040 157.230 42.300 157.490 ;
        RECT 60.440 157.230 60.700 157.490 ;
        RECT 41.120 156.890 41.380 157.150 ;
        RECT 51.240 156.890 51.500 157.150 ;
        RECT 51.700 156.890 51.960 157.150 ;
        RECT 53.080 156.890 53.340 157.150 ;
        RECT 57.220 156.890 57.480 157.150 ;
        RECT 71.020 156.890 71.280 157.150 ;
        RECT 74.240 156.890 74.500 157.150 ;
        RECT 76.540 156.890 76.800 157.150 ;
        RECT 78.380 156.890 78.640 157.150 ;
        RECT 84.360 157.570 84.620 157.830 ;
        RECT 85.740 157.570 86.000 157.830 ;
        RECT 91.720 157.910 91.980 158.170 ;
        RECT 88.040 157.570 88.300 157.830 ;
        RECT 83.440 156.890 83.700 157.150 ;
        RECT 87.580 157.230 87.840 157.490 ;
        RECT 89.420 157.230 89.680 157.490 ;
        RECT 90.340 157.230 90.600 157.490 ;
        RECT 92.640 157.910 92.900 158.170 ;
        RECT 105.060 158.250 105.320 158.510 ;
        RECT 124.840 158.250 125.100 158.510 ;
        RECT 95.400 157.570 95.660 157.830 ;
        RECT 99.080 157.910 99.340 158.170 ;
        RECT 101.840 157.910 102.100 158.170 ;
        RECT 103.220 157.910 103.480 158.170 ;
        RECT 98.160 157.570 98.420 157.830 ;
        RECT 95.860 156.890 96.120 157.150 ;
        RECT 101.380 157.570 101.640 157.830 ;
        RECT 110.120 157.570 110.380 157.830 ;
        RECT 101.380 156.890 101.640 157.150 ;
        RECT 109.200 156.890 109.460 157.150 ;
        RECT 45.190 156.380 45.450 156.640 ;
        RECT 45.510 156.380 45.770 156.640 ;
        RECT 45.830 156.380 46.090 156.640 ;
        RECT 46.150 156.380 46.410 156.640 ;
        RECT 46.470 156.380 46.730 156.640 ;
        RECT 80.035 156.380 80.295 156.640 ;
        RECT 80.355 156.380 80.615 156.640 ;
        RECT 80.675 156.380 80.935 156.640 ;
        RECT 80.995 156.380 81.255 156.640 ;
        RECT 81.315 156.380 81.575 156.640 ;
        RECT 114.880 156.380 115.140 156.640 ;
        RECT 115.200 156.380 115.460 156.640 ;
        RECT 115.520 156.380 115.780 156.640 ;
        RECT 115.840 156.380 116.100 156.640 ;
        RECT 116.160 156.380 116.420 156.640 ;
        RECT 149.725 156.380 149.985 156.640 ;
        RECT 150.045 156.380 150.305 156.640 ;
        RECT 150.365 156.380 150.625 156.640 ;
        RECT 150.685 156.380 150.945 156.640 ;
        RECT 151.005 156.380 151.265 156.640 ;
        RECT 25.480 155.870 25.740 156.130 ;
        RECT 32.380 155.870 32.640 156.130 ;
        RECT 31.460 155.530 31.720 155.790 ;
        RECT 19.040 155.190 19.300 155.450 ;
        RECT 31.000 155.190 31.260 155.450 ;
        RECT 31.920 155.190 32.180 155.450 ;
        RECT 34.220 155.190 34.480 155.450 ;
        RECT 39.740 155.530 40.000 155.790 ;
        RECT 42.500 155.870 42.760 156.130 ;
        RECT 44.800 155.530 45.060 155.790 ;
        RECT 35.140 154.850 35.400 155.110 ;
        RECT 39.280 155.190 39.540 155.450 ;
        RECT 38.360 154.850 38.620 155.110 ;
        RECT 41.120 154.850 41.380 155.110 ;
        RECT 42.040 155.190 42.300 155.450 ;
        RECT 42.960 155.190 43.220 155.450 ;
        RECT 45.260 155.190 45.520 155.450 ;
        RECT 49.860 155.870 50.120 156.130 ;
        RECT 48.480 155.530 48.740 155.790 ;
        RECT 53.080 155.190 53.340 155.450 ;
        RECT 57.220 155.870 57.480 156.130 ;
        RECT 59.980 155.870 60.240 156.130 ;
        RECT 65.960 155.870 66.220 156.130 ;
        RECT 71.020 155.870 71.280 156.130 ;
        RECT 73.780 155.870 74.040 156.130 ;
        RECT 56.760 155.530 57.020 155.790 ;
        RECT 56.300 155.190 56.560 155.450 ;
        RECT 64.580 155.190 64.840 155.450 ;
        RECT 82.980 155.530 83.240 155.790 ;
        RECT 83.440 155.530 83.700 155.790 ;
        RECT 85.740 155.870 86.000 156.130 ;
        RECT 95.860 155.870 96.120 156.130 ;
        RECT 98.160 155.870 98.420 156.130 ;
        RECT 101.840 155.870 102.100 156.130 ;
        RECT 84.360 155.530 84.620 155.790 ;
        RECT 86.200 155.530 86.460 155.790 ;
        RECT 89.420 155.530 89.680 155.790 ;
        RECT 91.260 155.530 91.520 155.790 ;
        RECT 87.580 155.190 87.840 155.450 ;
        RECT 88.040 155.190 88.300 155.450 ;
        RECT 90.340 155.190 90.600 155.450 ;
        RECT 38.820 154.510 39.080 154.770 ;
        RECT 40.200 154.510 40.460 154.770 ;
        RECT 75.620 154.850 75.880 155.110 ;
        RECT 84.820 154.850 85.080 155.110 ;
        RECT 43.880 154.510 44.140 154.770 ;
        RECT 51.700 154.510 51.960 154.770 ;
        RECT 17.200 154.170 17.460 154.430 ;
        RECT 31.920 154.170 32.180 154.430 ;
        RECT 61.820 154.170 62.080 154.430 ;
        RECT 73.320 154.170 73.580 154.430 ;
        RECT 73.780 154.170 74.040 154.430 ;
        RECT 75.160 154.170 75.420 154.430 ;
        RECT 91.260 154.510 91.520 154.770 ;
        RECT 94.480 154.850 94.740 155.110 ;
        RECT 95.860 154.850 96.120 155.110 ;
        RECT 101.840 155.190 102.100 155.450 ;
        RECT 107.820 155.190 108.080 155.450 ;
        RECT 109.200 155.190 109.460 155.450 ;
        RECT 94.940 154.510 95.200 154.770 ;
        RECT 88.040 154.170 88.300 154.430 ;
        RECT 96.320 154.170 96.580 154.430 ;
        RECT 105.520 154.850 105.780 155.110 ;
        RECT 101.380 154.170 101.640 154.430 ;
        RECT 108.740 154.170 109.000 154.430 ;
        RECT 27.770 153.660 28.030 153.920 ;
        RECT 28.090 153.660 28.350 153.920 ;
        RECT 28.410 153.660 28.670 153.920 ;
        RECT 28.730 153.660 28.990 153.920 ;
        RECT 29.050 153.660 29.310 153.920 ;
        RECT 62.615 153.660 62.875 153.920 ;
        RECT 62.935 153.660 63.195 153.920 ;
        RECT 63.255 153.660 63.515 153.920 ;
        RECT 63.575 153.660 63.835 153.920 ;
        RECT 63.895 153.660 64.155 153.920 ;
        RECT 97.460 153.660 97.720 153.920 ;
        RECT 97.780 153.660 98.040 153.920 ;
        RECT 98.100 153.660 98.360 153.920 ;
        RECT 98.420 153.660 98.680 153.920 ;
        RECT 98.740 153.660 99.000 153.920 ;
        RECT 132.305 153.660 132.565 153.920 ;
        RECT 132.625 153.660 132.885 153.920 ;
        RECT 132.945 153.660 133.205 153.920 ;
        RECT 133.265 153.660 133.525 153.920 ;
        RECT 133.585 153.660 133.845 153.920 ;
        RECT 31.000 153.150 31.260 153.410 ;
        RECT 42.040 153.150 42.300 153.410 ;
        RECT 42.500 153.150 42.760 153.410 ;
        RECT 42.960 153.150 43.220 153.410 ;
        RECT 45.260 153.150 45.520 153.410 ;
        RECT 56.300 153.150 56.560 153.410 ;
        RECT 84.820 153.150 85.080 153.410 ;
        RECT 30.540 152.810 30.800 153.070 ;
        RECT 24.560 152.470 24.820 152.730 ;
        RECT 16.280 152.130 16.540 152.390 ;
        RECT 17.200 152.130 17.460 152.390 ;
        RECT 27.320 152.130 27.580 152.390 ;
        RECT 29.620 151.450 29.880 151.710 ;
        RECT 32.380 152.130 32.640 152.390 ;
        RECT 35.140 152.130 35.400 152.390 ;
        RECT 40.200 152.130 40.460 152.390 ;
        RECT 51.700 152.810 51.960 153.070 ;
        RECT 31.460 151.790 31.720 152.050 ;
        RECT 36.980 151.790 37.240 152.050 ;
        RECT 38.820 151.790 39.080 152.050 ;
        RECT 41.120 151.790 41.380 152.050 ;
        RECT 43.880 151.790 44.140 152.050 ;
        RECT 51.240 152.130 51.500 152.390 ;
        RECT 52.160 151.790 52.420 152.050 ;
        RECT 53.080 152.130 53.340 152.390 ;
        RECT 67.800 152.470 68.060 152.730 ;
        RECT 82.520 152.470 82.780 152.730 ;
        RECT 61.820 152.130 62.080 152.390 ;
        RECT 64.580 152.130 64.840 152.390 ;
        RECT 66.420 152.130 66.680 152.390 ;
        RECT 73.320 152.130 73.580 152.390 ;
        RECT 74.240 152.130 74.500 152.390 ;
        RECT 74.700 152.130 74.960 152.390 ;
        RECT 78.380 152.130 78.640 152.390 ;
        RECT 76.080 151.790 76.340 152.050 ;
        RECT 86.200 152.130 86.460 152.390 ;
        RECT 87.120 152.810 87.380 153.070 ;
        RECT 95.400 153.150 95.660 153.410 ;
        RECT 98.160 153.150 98.420 153.410 ;
        RECT 102.300 153.150 102.560 153.410 ;
        RECT 111.040 152.810 111.300 153.070 ;
        RECT 91.260 152.130 91.520 152.390 ;
        RECT 93.560 152.130 93.820 152.390 ;
        RECT 94.020 152.130 94.280 152.390 ;
        RECT 31.920 151.450 32.180 151.710 ;
        RECT 44.800 151.450 45.060 151.710 ;
        RECT 57.680 151.450 57.940 151.710 ;
        RECT 65.500 151.450 65.760 151.710 ;
        RECT 72.400 151.450 72.660 151.710 ;
        RECT 73.780 151.450 74.040 151.710 ;
        RECT 76.540 151.450 76.800 151.710 ;
        RECT 83.440 151.450 83.700 151.710 ;
        RECT 95.860 152.130 96.120 152.390 ;
        RECT 96.320 151.450 96.580 151.710 ;
        RECT 118.860 152.470 119.120 152.730 ;
        RECT 123.000 152.470 123.260 152.730 ;
        RECT 97.700 152.130 97.960 152.390 ;
        RECT 100.920 152.130 101.180 152.390 ;
        RECT 109.200 151.790 109.460 152.050 ;
        RECT 97.240 151.450 97.500 151.710 ;
        RECT 45.190 150.940 45.450 151.200 ;
        RECT 45.510 150.940 45.770 151.200 ;
        RECT 45.830 150.940 46.090 151.200 ;
        RECT 46.150 150.940 46.410 151.200 ;
        RECT 46.470 150.940 46.730 151.200 ;
        RECT 80.035 150.940 80.295 151.200 ;
        RECT 80.355 150.940 80.615 151.200 ;
        RECT 80.675 150.940 80.935 151.200 ;
        RECT 80.995 150.940 81.255 151.200 ;
        RECT 81.315 150.940 81.575 151.200 ;
        RECT 114.880 150.940 115.140 151.200 ;
        RECT 115.200 150.940 115.460 151.200 ;
        RECT 115.520 150.940 115.780 151.200 ;
        RECT 115.840 150.940 116.100 151.200 ;
        RECT 116.160 150.940 116.420 151.200 ;
        RECT 149.725 150.940 149.985 151.200 ;
        RECT 150.045 150.940 150.305 151.200 ;
        RECT 150.365 150.940 150.625 151.200 ;
        RECT 150.685 150.940 150.945 151.200 ;
        RECT 151.005 150.940 151.265 151.200 ;
        RECT 19.040 150.430 19.300 150.690 ;
        RECT 29.620 150.430 29.880 150.690 ;
        RECT 40.660 150.430 40.920 150.690 ;
        RECT 74.240 150.430 74.500 150.690 ;
        RECT 76.540 150.430 76.800 150.690 ;
        RECT 94.940 150.430 95.200 150.690 ;
        RECT 98.160 150.430 98.420 150.690 ;
        RECT 108.740 150.430 109.000 150.690 ;
        RECT 109.200 150.430 109.460 150.690 ;
        RECT 111.040 150.430 111.300 150.690 ;
        RECT 31.000 149.750 31.260 150.010 ;
        RECT 35.600 149.750 35.860 150.010 ;
        RECT 38.820 149.750 39.080 150.010 ;
        RECT 20.420 149.410 20.680 149.670 ;
        RECT 34.220 149.410 34.480 149.670 ;
        RECT 40.200 149.750 40.460 150.010 ;
        RECT 45.720 149.750 45.980 150.010 ;
        RECT 75.620 149.750 75.880 150.010 ;
        RECT 51.240 149.410 51.500 149.670 ;
        RECT 51.700 149.410 51.960 149.670 ;
        RECT 79.300 149.410 79.560 149.670 ;
        RECT 27.320 149.070 27.580 149.330 ;
        RECT 56.760 149.070 57.020 149.330 ;
        RECT 61.820 149.070 62.080 149.330 ;
        RECT 93.560 149.750 93.820 150.010 ;
        RECT 94.480 149.750 94.740 150.010 ;
        RECT 99.080 149.410 99.340 149.670 ;
        RECT 101.840 149.410 102.100 149.670 ;
        RECT 103.680 149.750 103.940 150.010 ;
        RECT 105.060 149.750 105.320 150.010 ;
        RECT 107.820 149.750 108.080 150.010 ;
        RECT 108.280 149.750 108.540 150.010 ;
        RECT 111.500 149.750 111.760 150.010 ;
        RECT 113.340 150.090 113.600 150.350 ;
        RECT 120.700 150.090 120.960 150.350 ;
        RECT 114.720 149.750 114.980 150.010 ;
        RECT 123.000 149.750 123.260 150.010 ;
        RECT 25.020 148.730 25.280 148.990 ;
        RECT 37.440 148.730 37.700 148.990 ;
        RECT 68.260 148.730 68.520 148.990 ;
        RECT 94.940 148.730 95.200 148.990 ;
        RECT 103.680 148.730 103.940 148.990 ;
        RECT 109.660 148.730 109.920 148.990 ;
        RECT 110.120 148.730 110.380 148.990 ;
        RECT 116.560 148.730 116.820 148.990 ;
        RECT 27.770 148.220 28.030 148.480 ;
        RECT 28.090 148.220 28.350 148.480 ;
        RECT 28.410 148.220 28.670 148.480 ;
        RECT 28.730 148.220 28.990 148.480 ;
        RECT 29.050 148.220 29.310 148.480 ;
        RECT 62.615 148.220 62.875 148.480 ;
        RECT 62.935 148.220 63.195 148.480 ;
        RECT 63.255 148.220 63.515 148.480 ;
        RECT 63.575 148.220 63.835 148.480 ;
        RECT 63.895 148.220 64.155 148.480 ;
        RECT 97.460 148.220 97.720 148.480 ;
        RECT 97.780 148.220 98.040 148.480 ;
        RECT 98.100 148.220 98.360 148.480 ;
        RECT 98.420 148.220 98.680 148.480 ;
        RECT 98.740 148.220 99.000 148.480 ;
        RECT 132.305 148.220 132.565 148.480 ;
        RECT 132.625 148.220 132.885 148.480 ;
        RECT 132.945 148.220 133.205 148.480 ;
        RECT 133.265 148.220 133.525 148.480 ;
        RECT 133.585 148.220 133.845 148.480 ;
        RECT 30.540 147.710 30.800 147.970 ;
        RECT 45.720 147.710 45.980 147.970 ;
        RECT 51.240 147.710 51.500 147.970 ;
        RECT 24.100 147.370 24.360 147.630 ;
        RECT 23.640 146.690 23.900 146.950 ;
        RECT 26.860 146.690 27.120 146.950 ;
        RECT 27.780 146.690 28.040 146.950 ;
        RECT 31.000 146.690 31.260 146.950 ;
        RECT 34.220 146.690 34.480 146.950 ;
        RECT 37.900 146.690 38.160 146.950 ;
        RECT 53.080 147.030 53.340 147.290 ;
        RECT 57.220 147.030 57.480 147.290 ;
        RECT 39.740 146.350 40.000 146.610 ;
        RECT 40.200 146.350 40.460 146.610 ;
        RECT 56.300 146.690 56.560 146.950 ;
        RECT 58.140 146.690 58.400 146.950 ;
        RECT 61.820 147.370 62.080 147.630 ;
        RECT 65.040 147.030 65.300 147.290 ;
        RECT 68.720 147.710 68.980 147.970 ;
        RECT 108.280 147.710 108.540 147.970 ;
        RECT 114.720 147.710 114.980 147.970 ;
        RECT 77.920 147.370 78.180 147.630 ;
        RECT 67.340 147.030 67.600 147.290 ;
        RECT 25.480 146.010 25.740 146.270 ;
        RECT 38.820 146.010 39.080 146.270 ;
        RECT 47.100 146.010 47.360 146.270 ;
        RECT 52.160 146.010 52.420 146.270 ;
        RECT 53.080 146.010 53.340 146.270 ;
        RECT 56.760 146.010 57.020 146.270 ;
        RECT 59.980 146.010 60.240 146.270 ;
        RECT 61.360 146.010 61.620 146.270 ;
        RECT 61.820 146.010 62.080 146.270 ;
        RECT 65.960 146.010 66.220 146.270 ;
        RECT 66.880 146.690 67.140 146.950 ;
        RECT 68.260 146.690 68.520 146.950 ;
        RECT 70.100 146.690 70.360 146.950 ;
        RECT 77.460 146.350 77.720 146.610 ;
        RECT 78.840 146.690 79.100 146.950 ;
        RECT 82.520 146.690 82.780 146.950 ;
        RECT 83.440 146.690 83.700 146.950 ;
        RECT 86.660 146.690 86.920 146.950 ;
        RECT 94.480 147.370 94.740 147.630 ;
        RECT 102.300 147.370 102.560 147.630 ;
        RECT 100.000 147.030 100.260 147.290 ;
        RECT 88.960 146.350 89.220 146.610 ;
        RECT 93.560 146.350 93.820 146.610 ;
        RECT 109.660 147.370 109.920 147.630 ;
        RECT 111.500 147.030 111.760 147.290 ;
        RECT 110.580 146.690 110.840 146.950 ;
        RECT 113.340 146.690 113.600 146.950 ;
        RECT 111.500 146.350 111.760 146.610 ;
        RECT 66.880 146.010 67.140 146.270 ;
        RECT 77.920 146.010 78.180 146.270 ;
        RECT 78.380 146.010 78.640 146.270 ;
        RECT 79.300 146.010 79.560 146.270 ;
        RECT 100.000 146.010 100.260 146.270 ;
        RECT 117.940 146.690 118.200 146.950 ;
        RECT 119.320 146.690 119.580 146.950 ;
        RECT 116.560 146.350 116.820 146.610 ;
        RECT 45.190 145.500 45.450 145.760 ;
        RECT 45.510 145.500 45.770 145.760 ;
        RECT 45.830 145.500 46.090 145.760 ;
        RECT 46.150 145.500 46.410 145.760 ;
        RECT 46.470 145.500 46.730 145.760 ;
        RECT 80.035 145.500 80.295 145.760 ;
        RECT 80.355 145.500 80.615 145.760 ;
        RECT 80.675 145.500 80.935 145.760 ;
        RECT 80.995 145.500 81.255 145.760 ;
        RECT 81.315 145.500 81.575 145.760 ;
        RECT 114.880 145.500 115.140 145.760 ;
        RECT 115.200 145.500 115.460 145.760 ;
        RECT 115.520 145.500 115.780 145.760 ;
        RECT 115.840 145.500 116.100 145.760 ;
        RECT 116.160 145.500 116.420 145.760 ;
        RECT 149.725 145.500 149.985 145.760 ;
        RECT 150.045 145.500 150.305 145.760 ;
        RECT 150.365 145.500 150.625 145.760 ;
        RECT 150.685 145.500 150.945 145.760 ;
        RECT 151.005 145.500 151.265 145.760 ;
        RECT 24.100 144.990 24.360 145.250 ;
        RECT 25.480 144.990 25.740 145.250 ;
        RECT 39.740 144.990 40.000 145.250 ;
        RECT 57.680 144.990 57.940 145.250 ;
        RECT 61.360 144.990 61.620 145.250 ;
        RECT 65.040 144.990 65.300 145.250 ;
        RECT 70.100 144.990 70.360 145.250 ;
        RECT 77.460 144.990 77.720 145.250 ;
        RECT 78.380 144.990 78.640 145.250 ;
        RECT 86.200 144.990 86.460 145.250 ;
        RECT 88.960 144.990 89.220 145.250 ;
        RECT 94.940 144.990 95.200 145.250 ;
        RECT 35.600 144.650 35.860 144.910 ;
        RECT 24.560 143.970 24.820 144.230 ;
        RECT 27.320 144.310 27.580 144.570 ;
        RECT 38.360 144.310 38.620 144.570 ;
        RECT 47.100 144.310 47.360 144.570 ;
        RECT 51.700 144.310 51.960 144.570 ;
        RECT 61.820 144.650 62.080 144.910 ;
        RECT 66.880 144.650 67.140 144.910 ;
        RECT 72.400 144.650 72.660 144.910 ;
        RECT 65.040 144.310 65.300 144.570 ;
        RECT 78.840 144.310 79.100 144.570 ;
        RECT 82.060 144.310 82.320 144.570 ;
        RECT 31.460 143.970 31.720 144.230 ;
        RECT 37.440 143.970 37.700 144.230 ;
        RECT 48.940 143.970 49.200 144.230 ;
        RECT 53.080 143.970 53.340 144.230 ;
        RECT 58.140 143.970 58.400 144.230 ;
        RECT 56.760 143.630 57.020 143.890 ;
        RECT 59.060 143.630 59.320 143.890 ;
        RECT 60.900 143.290 61.160 143.550 ;
        RECT 61.820 143.290 62.080 143.550 ;
        RECT 64.580 143.290 64.840 143.550 ;
        RECT 78.380 143.970 78.640 144.230 ;
        RECT 93.100 144.310 93.360 144.570 ;
        RECT 103.220 144.650 103.480 144.910 ;
        RECT 103.680 144.310 103.940 144.570 ;
        RECT 116.560 144.310 116.820 144.570 ;
        RECT 82.980 143.630 83.240 143.890 ;
        RECT 102.300 143.630 102.560 143.890 ;
        RECT 83.440 143.290 83.700 143.550 ;
        RECT 87.580 143.290 87.840 143.550 ;
        RECT 105.060 143.290 105.320 143.550 ;
        RECT 119.780 143.290 120.040 143.550 ;
        RECT 27.770 142.780 28.030 143.040 ;
        RECT 28.090 142.780 28.350 143.040 ;
        RECT 28.410 142.780 28.670 143.040 ;
        RECT 28.730 142.780 28.990 143.040 ;
        RECT 29.050 142.780 29.310 143.040 ;
        RECT 62.615 142.780 62.875 143.040 ;
        RECT 62.935 142.780 63.195 143.040 ;
        RECT 63.255 142.780 63.515 143.040 ;
        RECT 63.575 142.780 63.835 143.040 ;
        RECT 63.895 142.780 64.155 143.040 ;
        RECT 97.460 142.780 97.720 143.040 ;
        RECT 97.780 142.780 98.040 143.040 ;
        RECT 98.100 142.780 98.360 143.040 ;
        RECT 98.420 142.780 98.680 143.040 ;
        RECT 98.740 142.780 99.000 143.040 ;
        RECT 132.305 142.780 132.565 143.040 ;
        RECT 132.625 142.780 132.885 143.040 ;
        RECT 132.945 142.780 133.205 143.040 ;
        RECT 133.265 142.780 133.525 143.040 ;
        RECT 133.585 142.780 133.845 143.040 ;
        RECT 38.360 142.270 38.620 142.530 ;
        RECT 47.100 142.270 47.360 142.530 ;
        RECT 53.080 142.270 53.340 142.530 ;
        RECT 65.040 142.270 65.300 142.530 ;
        RECT 105.060 142.270 105.320 142.530 ;
        RECT 18.580 141.250 18.840 141.510 ;
        RECT 24.560 140.910 24.820 141.170 ;
        RECT 28.700 141.250 28.960 141.510 ;
        RECT 31.000 141.250 31.260 141.510 ;
        RECT 32.380 141.250 32.640 141.510 ;
        RECT 36.980 141.250 37.240 141.510 ;
        RECT 60.900 141.930 61.160 142.190 ;
        RECT 33.760 140.910 34.020 141.170 ;
        RECT 36.520 140.910 36.780 141.170 ;
        RECT 17.200 140.570 17.460 140.830 ;
        RECT 29.160 140.570 29.420 140.830 ;
        RECT 31.000 140.570 31.260 140.830 ;
        RECT 31.920 140.570 32.180 140.830 ;
        RECT 44.340 140.910 44.600 141.170 ;
        RECT 65.500 141.590 65.760 141.850 ;
        RECT 94.480 141.590 94.740 141.850 ;
        RECT 103.220 141.590 103.480 141.850 ;
        RECT 57.680 141.250 57.940 141.510 ;
        RECT 61.820 141.250 62.080 141.510 ;
        RECT 76.540 141.250 76.800 141.510 ;
        RECT 77.460 141.250 77.720 141.510 ;
        RECT 100.000 141.250 100.260 141.510 ;
        RECT 103.680 141.250 103.940 141.510 ;
        RECT 105.520 141.250 105.780 141.510 ;
        RECT 105.980 141.250 106.240 141.510 ;
        RECT 107.820 141.250 108.080 141.510 ;
        RECT 110.120 141.250 110.380 141.510 ;
        RECT 111.500 141.250 111.760 141.510 ;
        RECT 44.800 140.570 45.060 140.830 ;
        RECT 47.100 140.570 47.360 140.830 ;
        RECT 75.620 140.570 75.880 140.830 ;
        RECT 77.000 140.570 77.260 140.830 ;
        RECT 102.760 140.570 103.020 140.830 ;
        RECT 105.520 140.570 105.780 140.830 ;
        RECT 108.280 140.570 108.540 140.830 ;
        RECT 109.660 140.570 109.920 140.830 ;
        RECT 118.400 140.910 118.660 141.170 ;
        RECT 119.780 140.910 120.040 141.170 ;
        RECT 113.800 140.570 114.060 140.830 ;
        RECT 45.190 140.060 45.450 140.320 ;
        RECT 45.510 140.060 45.770 140.320 ;
        RECT 45.830 140.060 46.090 140.320 ;
        RECT 46.150 140.060 46.410 140.320 ;
        RECT 46.470 140.060 46.730 140.320 ;
        RECT 80.035 140.060 80.295 140.320 ;
        RECT 80.355 140.060 80.615 140.320 ;
        RECT 80.675 140.060 80.935 140.320 ;
        RECT 80.995 140.060 81.255 140.320 ;
        RECT 81.315 140.060 81.575 140.320 ;
        RECT 114.880 140.060 115.140 140.320 ;
        RECT 115.200 140.060 115.460 140.320 ;
        RECT 115.520 140.060 115.780 140.320 ;
        RECT 115.840 140.060 116.100 140.320 ;
        RECT 116.160 140.060 116.420 140.320 ;
        RECT 149.725 140.060 149.985 140.320 ;
        RECT 150.045 140.060 150.305 140.320 ;
        RECT 150.365 140.060 150.625 140.320 ;
        RECT 150.685 140.060 150.945 140.320 ;
        RECT 151.005 140.060 151.265 140.320 ;
        RECT 16.280 139.210 16.540 139.470 ;
        RECT 37.900 139.550 38.160 139.810 ;
        RECT 23.640 139.210 23.900 139.470 ;
        RECT 17.200 138.870 17.460 139.130 ;
        RECT 28.700 139.210 28.960 139.470 ;
        RECT 29.160 139.210 29.420 139.470 ;
        RECT 33.760 139.210 34.020 139.470 ;
        RECT 24.560 138.530 24.820 138.790 ;
        RECT 31.000 138.870 31.260 139.130 ;
        RECT 31.920 138.870 32.180 139.130 ;
        RECT 32.840 138.870 33.100 139.130 ;
        RECT 47.100 139.550 47.360 139.810 ;
        RECT 59.980 139.550 60.240 139.810 ;
        RECT 60.440 139.550 60.700 139.810 ;
        RECT 49.400 139.210 49.660 139.470 ;
        RECT 64.580 139.210 64.840 139.470 ;
        RECT 65.500 139.210 65.760 139.470 ;
        RECT 79.300 139.550 79.560 139.810 ;
        RECT 76.540 139.210 76.800 139.470 ;
        RECT 77.460 139.210 77.720 139.470 ;
        RECT 82.060 139.210 82.320 139.470 ;
        RECT 57.680 138.870 57.940 139.130 ;
        RECT 59.060 138.870 59.320 139.130 ;
        RECT 31.460 138.530 31.720 138.790 ;
        RECT 53.540 138.530 53.800 138.790 ;
        RECT 55.380 138.530 55.640 138.790 ;
        RECT 59.980 138.530 60.240 138.790 ;
        RECT 25.940 138.190 26.200 138.450 ;
        RECT 27.320 138.190 27.580 138.450 ;
        RECT 78.380 138.530 78.640 138.790 ;
        RECT 77.920 138.190 78.180 138.450 ;
        RECT 79.300 138.870 79.560 139.130 ;
        RECT 80.220 138.870 80.480 139.130 ;
        RECT 89.880 139.550 90.140 139.810 ;
        RECT 25.480 137.850 25.740 138.110 ;
        RECT 56.760 137.850 57.020 138.110 ;
        RECT 60.440 137.850 60.700 138.110 ;
        RECT 66.880 137.850 67.140 138.110 ;
        RECT 72.860 137.850 73.120 138.110 ;
        RECT 73.320 137.850 73.580 138.110 ;
        RECT 76.080 137.850 76.340 138.110 ;
        RECT 84.360 138.870 84.620 139.130 ;
        RECT 86.200 139.210 86.460 139.470 ;
        RECT 87.580 138.870 87.840 139.130 ;
        RECT 89.420 138.870 89.680 139.130 ;
        RECT 89.880 138.870 90.140 139.130 ;
        RECT 96.780 139.210 97.040 139.470 ;
        RECT 105.060 139.550 105.320 139.810 ;
        RECT 105.980 139.550 106.240 139.810 ;
        RECT 107.820 139.550 108.080 139.810 ;
        RECT 113.800 139.550 114.060 139.810 ;
        RECT 116.560 139.550 116.820 139.810 ;
        RECT 102.300 139.210 102.560 139.470 ;
        RECT 105.520 138.870 105.780 139.130 ;
        RECT 81.140 138.190 81.400 138.450 ;
        RECT 82.520 137.850 82.780 138.110 ;
        RECT 83.440 137.850 83.700 138.110 ;
        RECT 86.200 137.850 86.460 138.110 ;
        RECT 88.960 137.850 89.220 138.110 ;
        RECT 98.620 138.530 98.880 138.790 ;
        RECT 101.380 138.530 101.640 138.790 ;
        RECT 92.180 138.190 92.440 138.450 ;
        RECT 93.560 137.850 93.820 138.110 ;
        RECT 102.760 138.530 103.020 138.790 ;
        RECT 103.220 138.190 103.480 138.450 ;
        RECT 110.120 138.530 110.380 138.790 ;
        RECT 117.940 138.530 118.200 138.790 ;
        RECT 106.440 137.850 106.700 138.110 ;
        RECT 27.770 137.340 28.030 137.600 ;
        RECT 28.090 137.340 28.350 137.600 ;
        RECT 28.410 137.340 28.670 137.600 ;
        RECT 28.730 137.340 28.990 137.600 ;
        RECT 29.050 137.340 29.310 137.600 ;
        RECT 62.615 137.340 62.875 137.600 ;
        RECT 62.935 137.340 63.195 137.600 ;
        RECT 63.255 137.340 63.515 137.600 ;
        RECT 63.575 137.340 63.835 137.600 ;
        RECT 63.895 137.340 64.155 137.600 ;
        RECT 97.460 137.340 97.720 137.600 ;
        RECT 97.780 137.340 98.040 137.600 ;
        RECT 98.100 137.340 98.360 137.600 ;
        RECT 98.420 137.340 98.680 137.600 ;
        RECT 98.740 137.340 99.000 137.600 ;
        RECT 132.305 137.340 132.565 137.600 ;
        RECT 132.625 137.340 132.885 137.600 ;
        RECT 132.945 137.340 133.205 137.600 ;
        RECT 133.265 137.340 133.525 137.600 ;
        RECT 133.585 137.340 133.845 137.600 ;
        RECT 18.580 136.830 18.840 137.090 ;
        RECT 25.480 136.830 25.740 137.090 ;
        RECT 25.940 136.830 26.200 137.090 ;
        RECT 31.920 136.830 32.180 137.090 ;
        RECT 36.520 136.830 36.780 137.090 ;
        RECT 47.100 136.830 47.360 137.090 ;
        RECT 53.540 136.830 53.800 137.090 ;
        RECT 57.220 136.830 57.480 137.090 ;
        RECT 60.900 136.830 61.160 137.090 ;
        RECT 60.440 136.490 60.700 136.750 ;
        RECT 67.800 136.830 68.060 137.090 ;
        RECT 20.420 135.810 20.680 136.070 ;
        RECT 27.320 135.810 27.580 136.070 ;
        RECT 38.820 135.810 39.080 136.070 ;
        RECT 44.340 136.150 44.600 136.410 ;
        RECT 44.800 135.810 45.060 136.070 ;
        RECT 52.160 136.150 52.420 136.410 ;
        RECT 51.700 135.810 51.960 136.070 ;
        RECT 53.080 135.810 53.340 136.070 ;
        RECT 57.220 135.810 57.480 136.070 ;
        RECT 59.060 136.150 59.320 136.410 ;
        RECT 62.280 136.150 62.540 136.410 ;
        RECT 64.580 136.150 64.840 136.410 ;
        RECT 59.520 135.810 59.780 136.070 ;
        RECT 43.880 135.130 44.140 135.390 ;
        RECT 57.680 135.470 57.940 135.730 ;
        RECT 59.980 135.470 60.240 135.730 ;
        RECT 67.800 135.470 68.060 135.730 ;
        RECT 73.320 136.830 73.580 137.090 ;
        RECT 76.080 136.830 76.340 137.090 ;
        RECT 82.060 136.490 82.320 136.750 ;
        RECT 72.860 136.150 73.120 136.410 ;
        RECT 84.360 136.150 84.620 136.410 ;
        RECT 88.960 136.150 89.220 136.410 ;
        RECT 75.620 135.470 75.880 135.730 ;
        RECT 77.000 135.470 77.260 135.730 ;
        RECT 80.220 135.810 80.480 136.070 ;
        RECT 83.440 135.810 83.700 136.070 ;
        RECT 84.820 135.810 85.080 136.070 ;
        RECT 78.380 135.470 78.640 135.730 ;
        RECT 82.520 135.470 82.780 135.730 ;
        RECT 89.880 135.810 90.140 136.070 ;
        RECT 93.560 135.810 93.820 136.070 ;
        RECT 96.780 136.830 97.040 137.090 ;
        RECT 94.480 136.150 94.740 136.410 ;
        RECT 96.320 136.490 96.580 136.750 ;
        RECT 108.280 136.490 108.540 136.750 ;
        RECT 59.520 135.130 59.780 135.390 ;
        RECT 61.360 135.130 61.620 135.390 ;
        RECT 62.280 135.130 62.540 135.390 ;
        RECT 72.400 135.130 72.660 135.390 ;
        RECT 73.780 135.130 74.040 135.390 ;
        RECT 76.080 135.130 76.340 135.390 ;
        RECT 83.900 135.130 84.160 135.390 ;
        RECT 84.360 135.130 84.620 135.390 ;
        RECT 106.900 135.470 107.160 135.730 ;
        RECT 111.500 135.470 111.760 135.730 ;
        RECT 92.180 135.130 92.440 135.390 ;
        RECT 94.480 135.130 94.740 135.390 ;
        RECT 110.120 135.130 110.380 135.390 ;
        RECT 45.190 134.620 45.450 134.880 ;
        RECT 45.510 134.620 45.770 134.880 ;
        RECT 45.830 134.620 46.090 134.880 ;
        RECT 46.150 134.620 46.410 134.880 ;
        RECT 46.470 134.620 46.730 134.880 ;
        RECT 80.035 134.620 80.295 134.880 ;
        RECT 80.355 134.620 80.615 134.880 ;
        RECT 80.675 134.620 80.935 134.880 ;
        RECT 80.995 134.620 81.255 134.880 ;
        RECT 81.315 134.620 81.575 134.880 ;
        RECT 114.880 134.620 115.140 134.880 ;
        RECT 115.200 134.620 115.460 134.880 ;
        RECT 115.520 134.620 115.780 134.880 ;
        RECT 115.840 134.620 116.100 134.880 ;
        RECT 116.160 134.620 116.420 134.880 ;
        RECT 149.725 134.620 149.985 134.880 ;
        RECT 150.045 134.620 150.305 134.880 ;
        RECT 150.365 134.620 150.625 134.880 ;
        RECT 150.685 134.620 150.945 134.880 ;
        RECT 151.005 134.620 151.265 134.880 ;
        RECT 31.460 134.110 31.720 134.370 ;
        RECT 30.080 133.770 30.340 134.030 ;
        RECT 35.600 133.430 35.860 133.690 ;
        RECT 36.980 133.430 37.240 133.690 ;
        RECT 39.280 133.430 39.540 133.690 ;
        RECT 43.880 133.770 44.140 134.030 ;
        RECT 46.640 133.770 46.900 134.030 ;
        RECT 44.340 133.090 44.600 133.350 ;
        RECT 51.700 133.770 51.960 134.030 ;
        RECT 57.220 134.110 57.480 134.370 ;
        RECT 68.260 134.110 68.520 134.370 ;
        RECT 69.180 134.110 69.440 134.370 ;
        RECT 73.780 134.110 74.040 134.370 ;
        RECT 37.440 132.410 37.700 132.670 ;
        RECT 42.500 132.410 42.760 132.670 ;
        RECT 46.640 132.750 46.900 133.010 ;
        RECT 60.900 133.430 61.160 133.690 ;
        RECT 57.680 132.750 57.940 133.010 ;
        RECT 75.160 133.770 75.420 134.030 ;
        RECT 88.960 133.770 89.220 134.030 ;
        RECT 72.400 133.430 72.660 133.690 ;
        RECT 101.380 133.430 101.640 133.690 ;
        RECT 104.140 133.430 104.400 133.690 ;
        RECT 104.600 133.430 104.860 133.690 ;
        RECT 106.900 133.430 107.160 133.690 ;
        RECT 67.800 133.090 68.060 133.350 ;
        RECT 76.080 133.090 76.340 133.350 ;
        RECT 108.280 133.430 108.540 133.690 ;
        RECT 110.120 133.430 110.380 133.690 ;
        RECT 73.780 132.750 74.040 133.010 ;
        RECT 74.700 132.750 74.960 133.010 ;
        RECT 106.440 132.750 106.700 133.010 ;
        RECT 48.480 132.410 48.740 132.670 ;
        RECT 53.080 132.410 53.340 132.670 ;
        RECT 56.300 132.410 56.560 132.670 ;
        RECT 65.960 132.410 66.220 132.670 ;
        RECT 69.180 132.410 69.440 132.670 ;
        RECT 77.000 132.410 77.260 132.670 ;
        RECT 82.980 132.410 83.240 132.670 ;
        RECT 90.340 132.410 90.600 132.670 ;
        RECT 112.880 132.410 113.140 132.670 ;
        RECT 27.770 131.900 28.030 132.160 ;
        RECT 28.090 131.900 28.350 132.160 ;
        RECT 28.410 131.900 28.670 132.160 ;
        RECT 28.730 131.900 28.990 132.160 ;
        RECT 29.050 131.900 29.310 132.160 ;
        RECT 62.615 131.900 62.875 132.160 ;
        RECT 62.935 131.900 63.195 132.160 ;
        RECT 63.255 131.900 63.515 132.160 ;
        RECT 63.575 131.900 63.835 132.160 ;
        RECT 63.895 131.900 64.155 132.160 ;
        RECT 97.460 131.900 97.720 132.160 ;
        RECT 97.780 131.900 98.040 132.160 ;
        RECT 98.100 131.900 98.360 132.160 ;
        RECT 98.420 131.900 98.680 132.160 ;
        RECT 98.740 131.900 99.000 132.160 ;
        RECT 132.305 131.900 132.565 132.160 ;
        RECT 132.625 131.900 132.885 132.160 ;
        RECT 132.945 131.900 133.205 132.160 ;
        RECT 133.265 131.900 133.525 132.160 ;
        RECT 133.585 131.900 133.845 132.160 ;
        RECT 27.320 131.390 27.580 131.650 ;
        RECT 37.440 131.390 37.700 131.650 ;
        RECT 42.500 131.390 42.760 131.650 ;
        RECT 37.900 130.370 38.160 130.630 ;
        RECT 41.580 130.370 41.840 130.630 ;
        RECT 48.480 131.390 48.740 131.650 ;
        RECT 54.920 131.390 55.180 131.650 ;
        RECT 56.760 131.390 57.020 131.650 ;
        RECT 61.360 131.390 61.620 131.650 ;
        RECT 65.960 131.390 66.220 131.650 ;
        RECT 56.300 131.050 56.560 131.310 ;
        RECT 44.340 130.030 44.600 130.290 ;
        RECT 48.940 130.370 49.200 130.630 ;
        RECT 55.380 130.710 55.640 130.970 ;
        RECT 57.680 131.050 57.940 131.310 ;
        RECT 57.680 130.370 57.940 130.630 ;
        RECT 57.220 130.030 57.480 130.290 ;
        RECT 75.620 130.710 75.880 130.970 ;
        RECT 42.040 129.690 42.300 129.950 ;
        RECT 43.420 129.690 43.680 129.950 ;
        RECT 54.460 129.690 54.720 129.950 ;
        RECT 59.060 129.690 59.320 129.950 ;
        RECT 60.440 129.690 60.700 129.950 ;
        RECT 66.420 129.690 66.680 129.950 ;
        RECT 73.780 130.030 74.040 130.290 ;
        RECT 75.160 130.370 75.420 130.630 ;
        RECT 82.980 131.390 83.240 131.650 ;
        RECT 78.840 131.050 79.100 131.310 ;
        RECT 82.060 130.370 82.320 130.630 ;
        RECT 84.360 131.050 84.620 131.310 ;
        RECT 99.080 131.390 99.340 131.650 ;
        RECT 85.280 130.370 85.540 130.630 ;
        RECT 104.600 131.050 104.860 131.310 ;
        RECT 104.140 130.710 104.400 130.970 ;
        RECT 118.400 131.390 118.660 131.650 ;
        RECT 102.300 130.370 102.560 130.630 ;
        RECT 112.880 130.370 113.140 130.630 ;
        RECT 79.300 130.030 79.560 130.290 ;
        RECT 84.820 130.030 85.080 130.290 ;
        RECT 74.700 129.690 74.960 129.950 ;
        RECT 76.080 129.690 76.340 129.950 ;
        RECT 85.280 129.690 85.540 129.950 ;
        RECT 86.200 129.690 86.460 129.950 ;
        RECT 89.420 129.690 89.680 129.950 ;
        RECT 45.190 129.180 45.450 129.440 ;
        RECT 45.510 129.180 45.770 129.440 ;
        RECT 45.830 129.180 46.090 129.440 ;
        RECT 46.150 129.180 46.410 129.440 ;
        RECT 46.470 129.180 46.730 129.440 ;
        RECT 80.035 129.180 80.295 129.440 ;
        RECT 80.355 129.180 80.615 129.440 ;
        RECT 80.675 129.180 80.935 129.440 ;
        RECT 80.995 129.180 81.255 129.440 ;
        RECT 81.315 129.180 81.575 129.440 ;
        RECT 114.880 129.180 115.140 129.440 ;
        RECT 115.200 129.180 115.460 129.440 ;
        RECT 115.520 129.180 115.780 129.440 ;
        RECT 115.840 129.180 116.100 129.440 ;
        RECT 116.160 129.180 116.420 129.440 ;
        RECT 149.725 129.180 149.985 129.440 ;
        RECT 150.045 129.180 150.305 129.440 ;
        RECT 150.365 129.180 150.625 129.440 ;
        RECT 150.685 129.180 150.945 129.440 ;
        RECT 151.005 129.180 151.265 129.440 ;
        RECT 39.280 128.670 39.540 128.930 ;
        RECT 53.080 128.670 53.340 128.930 ;
        RECT 54.460 128.670 54.720 128.930 ;
        RECT 42.040 127.990 42.300 128.250 ;
        RECT 45.260 126.970 45.520 127.230 ;
        RECT 49.400 127.650 49.660 127.910 ;
        RECT 52.160 127.990 52.420 128.250 ;
        RECT 54.000 128.330 54.260 128.590 ;
        RECT 59.060 128.330 59.320 128.590 ;
        RECT 66.880 128.670 67.140 128.930 ;
        RECT 75.160 128.670 75.420 128.930 ;
        RECT 79.300 128.670 79.560 128.930 ;
        RECT 54.920 127.650 55.180 127.910 ;
        RECT 54.460 127.310 54.720 127.570 ;
        RECT 60.440 127.990 60.700 128.250 ;
        RECT 67.340 127.990 67.600 128.250 ;
        RECT 64.580 127.650 64.840 127.910 ;
        RECT 78.840 128.330 79.100 128.590 ;
        RECT 82.520 128.670 82.780 128.930 ;
        RECT 84.820 128.670 85.080 128.930 ;
        RECT 86.200 128.670 86.460 128.930 ;
        RECT 89.420 128.670 89.680 128.930 ;
        RECT 85.280 128.330 85.540 128.590 ;
        RECT 82.520 127.990 82.780 128.250 ;
        RECT 83.440 127.990 83.700 128.250 ;
        RECT 90.340 128.330 90.600 128.590 ;
        RECT 60.900 127.310 61.160 127.570 ;
        RECT 65.040 127.310 65.300 127.570 ;
        RECT 82.520 127.310 82.780 127.570 ;
        RECT 92.640 127.650 92.900 127.910 ;
        RECT 59.060 126.970 59.320 127.230 ;
        RECT 99.080 127.990 99.340 128.250 ;
        RECT 88.960 126.970 89.220 127.230 ;
        RECT 91.260 126.970 91.520 127.230 ;
        RECT 27.770 126.460 28.030 126.720 ;
        RECT 28.090 126.460 28.350 126.720 ;
        RECT 28.410 126.460 28.670 126.720 ;
        RECT 28.730 126.460 28.990 126.720 ;
        RECT 29.050 126.460 29.310 126.720 ;
        RECT 62.615 126.460 62.875 126.720 ;
        RECT 62.935 126.460 63.195 126.720 ;
        RECT 63.255 126.460 63.515 126.720 ;
        RECT 63.575 126.460 63.835 126.720 ;
        RECT 63.895 126.460 64.155 126.720 ;
        RECT 97.460 126.460 97.720 126.720 ;
        RECT 97.780 126.460 98.040 126.720 ;
        RECT 98.100 126.460 98.360 126.720 ;
        RECT 98.420 126.460 98.680 126.720 ;
        RECT 98.740 126.460 99.000 126.720 ;
        RECT 132.305 126.460 132.565 126.720 ;
        RECT 132.625 126.460 132.885 126.720 ;
        RECT 132.945 126.460 133.205 126.720 ;
        RECT 133.265 126.460 133.525 126.720 ;
        RECT 133.585 126.460 133.845 126.720 ;
        RECT 43.420 125.950 43.680 126.210 ;
        RECT 65.040 125.950 65.300 126.210 ;
        RECT 67.340 125.950 67.600 126.210 ;
        RECT 92.640 125.950 92.900 126.210 ;
        RECT 66.420 125.270 66.680 125.530 ;
        RECT 91.260 125.270 91.520 125.530 ;
        RECT 41.580 124.930 41.840 125.190 ;
        RECT 45.260 124.590 45.520 124.850 ;
        RECT 64.580 124.930 64.840 125.190 ;
        RECT 96.320 124.930 96.580 125.190 ;
        RECT 59.060 124.590 59.320 124.850 ;
        RECT 47.560 124.250 47.820 124.510 ;
        RECT 45.190 123.740 45.450 124.000 ;
        RECT 45.510 123.740 45.770 124.000 ;
        RECT 45.830 123.740 46.090 124.000 ;
        RECT 46.150 123.740 46.410 124.000 ;
        RECT 46.470 123.740 46.730 124.000 ;
        RECT 80.035 123.740 80.295 124.000 ;
        RECT 80.355 123.740 80.615 124.000 ;
        RECT 80.675 123.740 80.935 124.000 ;
        RECT 80.995 123.740 81.255 124.000 ;
        RECT 81.315 123.740 81.575 124.000 ;
        RECT 114.880 123.740 115.140 124.000 ;
        RECT 115.200 123.740 115.460 124.000 ;
        RECT 115.520 123.740 115.780 124.000 ;
        RECT 115.840 123.740 116.100 124.000 ;
        RECT 116.160 123.740 116.420 124.000 ;
        RECT 149.725 123.740 149.985 124.000 ;
        RECT 150.045 123.740 150.305 124.000 ;
        RECT 150.365 123.740 150.625 124.000 ;
        RECT 150.685 123.740 150.945 124.000 ;
        RECT 151.005 123.740 151.265 124.000 ;
        RECT 54.460 123.230 54.720 123.490 ;
        RECT 49.400 122.890 49.660 123.150 ;
        RECT 47.560 122.550 47.820 122.810 ;
        RECT 27.770 121.020 28.030 121.280 ;
        RECT 28.090 121.020 28.350 121.280 ;
        RECT 28.410 121.020 28.670 121.280 ;
        RECT 28.730 121.020 28.990 121.280 ;
        RECT 29.050 121.020 29.310 121.280 ;
        RECT 62.615 121.020 62.875 121.280 ;
        RECT 62.935 121.020 63.195 121.280 ;
        RECT 63.255 121.020 63.515 121.280 ;
        RECT 63.575 121.020 63.835 121.280 ;
        RECT 63.895 121.020 64.155 121.280 ;
        RECT 97.460 121.020 97.720 121.280 ;
        RECT 97.780 121.020 98.040 121.280 ;
        RECT 98.100 121.020 98.360 121.280 ;
        RECT 98.420 121.020 98.680 121.280 ;
        RECT 98.740 121.020 99.000 121.280 ;
        RECT 132.305 121.020 132.565 121.280 ;
        RECT 132.625 121.020 132.885 121.280 ;
        RECT 132.945 121.020 133.205 121.280 ;
        RECT 133.265 121.020 133.525 121.280 ;
        RECT 133.585 121.020 133.845 121.280 ;
        RECT 45.190 118.300 45.450 118.560 ;
        RECT 45.510 118.300 45.770 118.560 ;
        RECT 45.830 118.300 46.090 118.560 ;
        RECT 46.150 118.300 46.410 118.560 ;
        RECT 46.470 118.300 46.730 118.560 ;
        RECT 80.035 118.300 80.295 118.560 ;
        RECT 80.355 118.300 80.615 118.560 ;
        RECT 80.675 118.300 80.935 118.560 ;
        RECT 80.995 118.300 81.255 118.560 ;
        RECT 81.315 118.300 81.575 118.560 ;
        RECT 114.880 118.300 115.140 118.560 ;
        RECT 115.200 118.300 115.460 118.560 ;
        RECT 115.520 118.300 115.780 118.560 ;
        RECT 115.840 118.300 116.100 118.560 ;
        RECT 116.160 118.300 116.420 118.560 ;
        RECT 149.725 118.300 149.985 118.560 ;
        RECT 150.045 118.300 150.305 118.560 ;
        RECT 150.365 118.300 150.625 118.560 ;
        RECT 150.685 118.300 150.945 118.560 ;
        RECT 151.005 118.300 151.265 118.560 ;
        RECT 27.770 115.580 28.030 115.840 ;
        RECT 28.090 115.580 28.350 115.840 ;
        RECT 28.410 115.580 28.670 115.840 ;
        RECT 28.730 115.580 28.990 115.840 ;
        RECT 29.050 115.580 29.310 115.840 ;
        RECT 62.615 115.580 62.875 115.840 ;
        RECT 62.935 115.580 63.195 115.840 ;
        RECT 63.255 115.580 63.515 115.840 ;
        RECT 63.575 115.580 63.835 115.840 ;
        RECT 63.895 115.580 64.155 115.840 ;
        RECT 97.460 115.580 97.720 115.840 ;
        RECT 97.780 115.580 98.040 115.840 ;
        RECT 98.100 115.580 98.360 115.840 ;
        RECT 98.420 115.580 98.680 115.840 ;
        RECT 98.740 115.580 99.000 115.840 ;
        RECT 132.305 115.580 132.565 115.840 ;
        RECT 132.625 115.580 132.885 115.840 ;
        RECT 132.945 115.580 133.205 115.840 ;
        RECT 133.265 115.580 133.525 115.840 ;
        RECT 133.585 115.580 133.845 115.840 ;
        RECT 45.190 112.860 45.450 113.120 ;
        RECT 45.510 112.860 45.770 113.120 ;
        RECT 45.830 112.860 46.090 113.120 ;
        RECT 46.150 112.860 46.410 113.120 ;
        RECT 46.470 112.860 46.730 113.120 ;
        RECT 80.035 112.860 80.295 113.120 ;
        RECT 80.355 112.860 80.615 113.120 ;
        RECT 80.675 112.860 80.935 113.120 ;
        RECT 80.995 112.860 81.255 113.120 ;
        RECT 81.315 112.860 81.575 113.120 ;
        RECT 114.880 112.860 115.140 113.120 ;
        RECT 115.200 112.860 115.460 113.120 ;
        RECT 115.520 112.860 115.780 113.120 ;
        RECT 115.840 112.860 116.100 113.120 ;
        RECT 116.160 112.860 116.420 113.120 ;
        RECT 149.725 112.860 149.985 113.120 ;
        RECT 150.045 112.860 150.305 113.120 ;
        RECT 150.365 112.860 150.625 113.120 ;
        RECT 150.685 112.860 150.945 113.120 ;
        RECT 151.005 112.860 151.265 113.120 ;
        RECT 27.770 110.140 28.030 110.400 ;
        RECT 28.090 110.140 28.350 110.400 ;
        RECT 28.410 110.140 28.670 110.400 ;
        RECT 28.730 110.140 28.990 110.400 ;
        RECT 29.050 110.140 29.310 110.400 ;
        RECT 62.615 110.140 62.875 110.400 ;
        RECT 62.935 110.140 63.195 110.400 ;
        RECT 63.255 110.140 63.515 110.400 ;
        RECT 63.575 110.140 63.835 110.400 ;
        RECT 63.895 110.140 64.155 110.400 ;
        RECT 97.460 110.140 97.720 110.400 ;
        RECT 97.780 110.140 98.040 110.400 ;
        RECT 98.100 110.140 98.360 110.400 ;
        RECT 98.420 110.140 98.680 110.400 ;
        RECT 98.740 110.140 99.000 110.400 ;
        RECT 132.305 110.140 132.565 110.400 ;
        RECT 132.625 110.140 132.885 110.400 ;
        RECT 132.945 110.140 133.205 110.400 ;
        RECT 133.265 110.140 133.525 110.400 ;
        RECT 133.585 110.140 133.845 110.400 ;
        RECT 45.190 107.420 45.450 107.680 ;
        RECT 45.510 107.420 45.770 107.680 ;
        RECT 45.830 107.420 46.090 107.680 ;
        RECT 46.150 107.420 46.410 107.680 ;
        RECT 46.470 107.420 46.730 107.680 ;
        RECT 80.035 107.420 80.295 107.680 ;
        RECT 80.355 107.420 80.615 107.680 ;
        RECT 80.675 107.420 80.935 107.680 ;
        RECT 80.995 107.420 81.255 107.680 ;
        RECT 81.315 107.420 81.575 107.680 ;
        RECT 114.880 107.420 115.140 107.680 ;
        RECT 115.200 107.420 115.460 107.680 ;
        RECT 115.520 107.420 115.780 107.680 ;
        RECT 115.840 107.420 116.100 107.680 ;
        RECT 116.160 107.420 116.420 107.680 ;
        RECT 149.725 107.420 149.985 107.680 ;
        RECT 150.045 107.420 150.305 107.680 ;
        RECT 150.365 107.420 150.625 107.680 ;
        RECT 150.685 107.420 150.945 107.680 ;
        RECT 151.005 107.420 151.265 107.680 ;
        RECT 27.770 104.700 28.030 104.960 ;
        RECT 28.090 104.700 28.350 104.960 ;
        RECT 28.410 104.700 28.670 104.960 ;
        RECT 28.730 104.700 28.990 104.960 ;
        RECT 29.050 104.700 29.310 104.960 ;
        RECT 62.615 104.700 62.875 104.960 ;
        RECT 62.935 104.700 63.195 104.960 ;
        RECT 63.255 104.700 63.515 104.960 ;
        RECT 63.575 104.700 63.835 104.960 ;
        RECT 63.895 104.700 64.155 104.960 ;
        RECT 97.460 104.700 97.720 104.960 ;
        RECT 97.780 104.700 98.040 104.960 ;
        RECT 98.100 104.700 98.360 104.960 ;
        RECT 98.420 104.700 98.680 104.960 ;
        RECT 98.740 104.700 99.000 104.960 ;
        RECT 132.305 104.700 132.565 104.960 ;
        RECT 132.625 104.700 132.885 104.960 ;
        RECT 132.945 104.700 133.205 104.960 ;
        RECT 133.265 104.700 133.525 104.960 ;
        RECT 133.585 104.700 133.845 104.960 ;
        RECT 45.190 101.980 45.450 102.240 ;
        RECT 45.510 101.980 45.770 102.240 ;
        RECT 45.830 101.980 46.090 102.240 ;
        RECT 46.150 101.980 46.410 102.240 ;
        RECT 46.470 101.980 46.730 102.240 ;
        RECT 80.035 101.980 80.295 102.240 ;
        RECT 80.355 101.980 80.615 102.240 ;
        RECT 80.675 101.980 80.935 102.240 ;
        RECT 80.995 101.980 81.255 102.240 ;
        RECT 81.315 101.980 81.575 102.240 ;
        RECT 114.880 101.980 115.140 102.240 ;
        RECT 115.200 101.980 115.460 102.240 ;
        RECT 115.520 101.980 115.780 102.240 ;
        RECT 115.840 101.980 116.100 102.240 ;
        RECT 116.160 101.980 116.420 102.240 ;
        RECT 149.725 101.980 149.985 102.240 ;
        RECT 150.045 101.980 150.305 102.240 ;
        RECT 150.365 101.980 150.625 102.240 ;
        RECT 150.685 101.980 150.945 102.240 ;
        RECT 151.005 101.980 151.265 102.240 ;
        RECT 27.770 99.260 28.030 99.520 ;
        RECT 28.090 99.260 28.350 99.520 ;
        RECT 28.410 99.260 28.670 99.520 ;
        RECT 28.730 99.260 28.990 99.520 ;
        RECT 29.050 99.260 29.310 99.520 ;
        RECT 62.615 99.260 62.875 99.520 ;
        RECT 62.935 99.260 63.195 99.520 ;
        RECT 63.255 99.260 63.515 99.520 ;
        RECT 63.575 99.260 63.835 99.520 ;
        RECT 63.895 99.260 64.155 99.520 ;
        RECT 97.460 99.260 97.720 99.520 ;
        RECT 97.780 99.260 98.040 99.520 ;
        RECT 98.100 99.260 98.360 99.520 ;
        RECT 98.420 99.260 98.680 99.520 ;
        RECT 98.740 99.260 99.000 99.520 ;
        RECT 132.305 99.260 132.565 99.520 ;
        RECT 132.625 99.260 132.885 99.520 ;
        RECT 132.945 99.260 133.205 99.520 ;
        RECT 133.265 99.260 133.525 99.520 ;
        RECT 133.585 99.260 133.845 99.520 ;
        RECT 45.190 96.540 45.450 96.800 ;
        RECT 45.510 96.540 45.770 96.800 ;
        RECT 45.830 96.540 46.090 96.800 ;
        RECT 46.150 96.540 46.410 96.800 ;
        RECT 46.470 96.540 46.730 96.800 ;
        RECT 80.035 96.540 80.295 96.800 ;
        RECT 80.355 96.540 80.615 96.800 ;
        RECT 80.675 96.540 80.935 96.800 ;
        RECT 80.995 96.540 81.255 96.800 ;
        RECT 81.315 96.540 81.575 96.800 ;
        RECT 114.880 96.540 115.140 96.800 ;
        RECT 115.200 96.540 115.460 96.800 ;
        RECT 115.520 96.540 115.780 96.800 ;
        RECT 115.840 96.540 116.100 96.800 ;
        RECT 116.160 96.540 116.420 96.800 ;
        RECT 149.725 96.540 149.985 96.800 ;
        RECT 150.045 96.540 150.305 96.800 ;
        RECT 150.365 96.540 150.625 96.800 ;
        RECT 150.685 96.540 150.945 96.800 ;
        RECT 151.005 96.540 151.265 96.800 ;
        RECT 27.770 93.820 28.030 94.080 ;
        RECT 28.090 93.820 28.350 94.080 ;
        RECT 28.410 93.820 28.670 94.080 ;
        RECT 28.730 93.820 28.990 94.080 ;
        RECT 29.050 93.820 29.310 94.080 ;
        RECT 62.615 93.820 62.875 94.080 ;
        RECT 62.935 93.820 63.195 94.080 ;
        RECT 63.255 93.820 63.515 94.080 ;
        RECT 63.575 93.820 63.835 94.080 ;
        RECT 63.895 93.820 64.155 94.080 ;
        RECT 97.460 93.820 97.720 94.080 ;
        RECT 97.780 93.820 98.040 94.080 ;
        RECT 98.100 93.820 98.360 94.080 ;
        RECT 98.420 93.820 98.680 94.080 ;
        RECT 98.740 93.820 99.000 94.080 ;
        RECT 132.305 93.820 132.565 94.080 ;
        RECT 132.625 93.820 132.885 94.080 ;
        RECT 132.945 93.820 133.205 94.080 ;
        RECT 133.265 93.820 133.525 94.080 ;
        RECT 133.585 93.820 133.845 94.080 ;
        RECT 45.190 91.100 45.450 91.360 ;
        RECT 45.510 91.100 45.770 91.360 ;
        RECT 45.830 91.100 46.090 91.360 ;
        RECT 46.150 91.100 46.410 91.360 ;
        RECT 46.470 91.100 46.730 91.360 ;
        RECT 80.035 91.100 80.295 91.360 ;
        RECT 80.355 91.100 80.615 91.360 ;
        RECT 80.675 91.100 80.935 91.360 ;
        RECT 80.995 91.100 81.255 91.360 ;
        RECT 81.315 91.100 81.575 91.360 ;
        RECT 114.880 91.100 115.140 91.360 ;
        RECT 115.200 91.100 115.460 91.360 ;
        RECT 115.520 91.100 115.780 91.360 ;
        RECT 115.840 91.100 116.100 91.360 ;
        RECT 116.160 91.100 116.420 91.360 ;
        RECT 149.725 91.100 149.985 91.360 ;
        RECT 150.045 91.100 150.305 91.360 ;
        RECT 150.365 91.100 150.625 91.360 ;
        RECT 150.685 91.100 150.945 91.360 ;
        RECT 151.005 91.100 151.265 91.360 ;
        RECT 27.770 88.380 28.030 88.640 ;
        RECT 28.090 88.380 28.350 88.640 ;
        RECT 28.410 88.380 28.670 88.640 ;
        RECT 28.730 88.380 28.990 88.640 ;
        RECT 29.050 88.380 29.310 88.640 ;
        RECT 62.615 88.380 62.875 88.640 ;
        RECT 62.935 88.380 63.195 88.640 ;
        RECT 63.255 88.380 63.515 88.640 ;
        RECT 63.575 88.380 63.835 88.640 ;
        RECT 63.895 88.380 64.155 88.640 ;
        RECT 97.460 88.380 97.720 88.640 ;
        RECT 97.780 88.380 98.040 88.640 ;
        RECT 98.100 88.380 98.360 88.640 ;
        RECT 98.420 88.380 98.680 88.640 ;
        RECT 98.740 88.380 99.000 88.640 ;
        RECT 132.305 88.380 132.565 88.640 ;
        RECT 132.625 88.380 132.885 88.640 ;
        RECT 132.945 88.380 133.205 88.640 ;
        RECT 133.265 88.380 133.525 88.640 ;
        RECT 133.585 88.380 133.845 88.640 ;
        RECT 45.190 85.660 45.450 85.920 ;
        RECT 45.510 85.660 45.770 85.920 ;
        RECT 45.830 85.660 46.090 85.920 ;
        RECT 46.150 85.660 46.410 85.920 ;
        RECT 46.470 85.660 46.730 85.920 ;
        RECT 80.035 85.660 80.295 85.920 ;
        RECT 80.355 85.660 80.615 85.920 ;
        RECT 80.675 85.660 80.935 85.920 ;
        RECT 80.995 85.660 81.255 85.920 ;
        RECT 81.315 85.660 81.575 85.920 ;
        RECT 114.880 85.660 115.140 85.920 ;
        RECT 115.200 85.660 115.460 85.920 ;
        RECT 115.520 85.660 115.780 85.920 ;
        RECT 115.840 85.660 116.100 85.920 ;
        RECT 116.160 85.660 116.420 85.920 ;
        RECT 149.725 85.660 149.985 85.920 ;
        RECT 150.045 85.660 150.305 85.920 ;
        RECT 150.365 85.660 150.625 85.920 ;
        RECT 150.685 85.660 150.945 85.920 ;
        RECT 151.005 85.660 151.265 85.920 ;
        RECT 27.770 82.940 28.030 83.200 ;
        RECT 28.090 82.940 28.350 83.200 ;
        RECT 28.410 82.940 28.670 83.200 ;
        RECT 28.730 82.940 28.990 83.200 ;
        RECT 29.050 82.940 29.310 83.200 ;
        RECT 62.615 82.940 62.875 83.200 ;
        RECT 62.935 82.940 63.195 83.200 ;
        RECT 63.255 82.940 63.515 83.200 ;
        RECT 63.575 82.940 63.835 83.200 ;
        RECT 63.895 82.940 64.155 83.200 ;
        RECT 97.460 82.940 97.720 83.200 ;
        RECT 97.780 82.940 98.040 83.200 ;
        RECT 98.100 82.940 98.360 83.200 ;
        RECT 98.420 82.940 98.680 83.200 ;
        RECT 98.740 82.940 99.000 83.200 ;
        RECT 132.305 82.940 132.565 83.200 ;
        RECT 132.625 82.940 132.885 83.200 ;
        RECT 132.945 82.940 133.205 83.200 ;
        RECT 133.265 82.940 133.525 83.200 ;
        RECT 133.585 82.940 133.845 83.200 ;
        RECT 45.190 80.220 45.450 80.480 ;
        RECT 45.510 80.220 45.770 80.480 ;
        RECT 45.830 80.220 46.090 80.480 ;
        RECT 46.150 80.220 46.410 80.480 ;
        RECT 46.470 80.220 46.730 80.480 ;
        RECT 80.035 80.220 80.295 80.480 ;
        RECT 80.355 80.220 80.615 80.480 ;
        RECT 80.675 80.220 80.935 80.480 ;
        RECT 80.995 80.220 81.255 80.480 ;
        RECT 81.315 80.220 81.575 80.480 ;
        RECT 114.880 80.220 115.140 80.480 ;
        RECT 115.200 80.220 115.460 80.480 ;
        RECT 115.520 80.220 115.780 80.480 ;
        RECT 115.840 80.220 116.100 80.480 ;
        RECT 116.160 80.220 116.420 80.480 ;
        RECT 149.725 80.220 149.985 80.480 ;
        RECT 150.045 80.220 150.305 80.480 ;
        RECT 150.365 80.220 150.625 80.480 ;
        RECT 150.685 80.220 150.945 80.480 ;
        RECT 151.005 80.220 151.265 80.480 ;
        RECT 27.770 77.500 28.030 77.760 ;
        RECT 28.090 77.500 28.350 77.760 ;
        RECT 28.410 77.500 28.670 77.760 ;
        RECT 28.730 77.500 28.990 77.760 ;
        RECT 29.050 77.500 29.310 77.760 ;
        RECT 62.615 77.500 62.875 77.760 ;
        RECT 62.935 77.500 63.195 77.760 ;
        RECT 63.255 77.500 63.515 77.760 ;
        RECT 63.575 77.500 63.835 77.760 ;
        RECT 63.895 77.500 64.155 77.760 ;
        RECT 97.460 77.500 97.720 77.760 ;
        RECT 97.780 77.500 98.040 77.760 ;
        RECT 98.100 77.500 98.360 77.760 ;
        RECT 98.420 77.500 98.680 77.760 ;
        RECT 98.740 77.500 99.000 77.760 ;
        RECT 132.305 77.500 132.565 77.760 ;
        RECT 132.625 77.500 132.885 77.760 ;
        RECT 132.945 77.500 133.205 77.760 ;
        RECT 133.265 77.500 133.525 77.760 ;
        RECT 133.585 77.500 133.845 77.760 ;
        RECT 45.190 74.780 45.450 75.040 ;
        RECT 45.510 74.780 45.770 75.040 ;
        RECT 45.830 74.780 46.090 75.040 ;
        RECT 46.150 74.780 46.410 75.040 ;
        RECT 46.470 74.780 46.730 75.040 ;
        RECT 80.035 74.780 80.295 75.040 ;
        RECT 80.355 74.780 80.615 75.040 ;
        RECT 80.675 74.780 80.935 75.040 ;
        RECT 80.995 74.780 81.255 75.040 ;
        RECT 81.315 74.780 81.575 75.040 ;
        RECT 114.880 74.780 115.140 75.040 ;
        RECT 115.200 74.780 115.460 75.040 ;
        RECT 115.520 74.780 115.780 75.040 ;
        RECT 115.840 74.780 116.100 75.040 ;
        RECT 116.160 74.780 116.420 75.040 ;
        RECT 149.725 74.780 149.985 75.040 ;
        RECT 150.045 74.780 150.305 75.040 ;
        RECT 150.365 74.780 150.625 75.040 ;
        RECT 150.685 74.780 150.945 75.040 ;
        RECT 151.005 74.780 151.265 75.040 ;
        RECT 55.340 55.020 76.610 59.300 ;
        RECT 95.400 55.090 105.220 59.770 ;
        RECT 62.000 49.290 62.940 49.650 ;
        RECT 64.680 49.300 65.590 49.700 ;
        RECT 78.760 49.160 79.750 49.640 ;
        RECT 78.760 48.380 79.750 48.860 ;
        RECT 78.750 47.580 79.740 48.060 ;
        RECT 64.630 46.910 65.640 47.280 ;
        RECT 77.540 46.870 78.230 47.310 ;
        RECT 78.750 46.800 79.740 47.280 ;
        RECT 81.010 47.560 82.950 51.910 ;
        RECT 117.310 54.830 134.530 58.370 ;
        RECT 62.000 44.650 62.940 45.010 ;
        RECT 64.680 44.630 65.590 45.030 ;
        RECT 78.740 46.010 79.730 46.490 ;
        RECT 78.750 45.210 79.740 45.690 ;
        RECT 78.770 44.420 79.760 44.900 ;
        RECT 64.630 42.350 65.640 42.720 ;
        RECT 78.760 43.640 79.750 44.120 ;
        RECT 78.770 42.840 79.760 43.320 ;
        RECT 62.010 40.080 62.950 40.440 ;
        RECT 64.670 40.060 65.580 40.460 ;
        RECT 73.610 42.040 74.520 42.400 ;
        RECT 78.760 42.060 79.750 42.540 ;
        RECT 78.770 41.260 79.760 41.740 ;
        RECT 106.985 41.740 108.715 43.470 ;
        RECT 73.590 39.820 74.540 40.100 ;
        RECT 64.630 37.770 65.640 38.140 ;
        RECT 78.760 40.480 79.750 40.960 ;
        RECT 78.750 39.680 79.740 40.160 ;
        RECT 73.600 37.490 74.510 37.850 ;
        RECT 78.760 38.900 79.750 39.380 ;
        RECT 78.760 38.100 79.750 38.580 ;
        RECT 62.030 35.540 62.940 35.840 ;
        RECT 64.690 35.490 65.590 35.840 ;
        RECT 78.760 37.310 79.750 37.790 ;
        RECT 95.110 38.110 96.110 39.110 ;
        RECT 97.400 38.090 98.400 39.090 ;
        RECT 99.690 38.070 100.690 39.070 ;
        RECT 101.950 38.090 102.950 39.090 ;
        RECT 104.240 38.090 105.240 39.090 ;
        RECT 64.760 34.690 65.790 35.110 ;
        RECT 61.960 31.020 62.410 33.080 ;
        RECT 63.890 31.040 64.310 33.030 ;
        RECT 73.580 35.110 74.540 35.620 ;
        RECT 78.770 36.520 79.760 37.000 ;
        RECT 78.760 35.730 79.750 36.210 ;
        RECT 124.230 48.890 125.170 49.250 ;
        RECT 126.910 48.900 127.820 49.300 ;
        RECT 140.990 48.760 141.980 49.240 ;
        RECT 140.990 47.980 141.980 48.460 ;
        RECT 140.980 47.180 141.970 47.660 ;
        RECT 126.860 46.510 127.870 46.880 ;
        RECT 139.770 46.470 140.460 46.910 ;
        RECT 140.980 46.400 141.970 46.880 ;
        RECT 143.240 47.160 145.180 51.510 ;
        RECT 124.230 44.250 125.170 44.610 ;
        RECT 126.910 44.230 127.820 44.630 ;
        RECT 140.970 45.610 141.960 46.090 ;
        RECT 140.980 44.810 141.970 45.290 ;
        RECT 141.000 44.020 141.990 44.500 ;
        RECT 126.860 41.950 127.870 42.320 ;
        RECT 140.990 43.240 141.980 43.720 ;
        RECT 141.000 42.440 141.990 42.920 ;
        RECT 124.240 39.680 125.180 40.040 ;
        RECT 126.900 39.660 127.810 40.060 ;
        RECT 135.840 41.640 136.750 42.000 ;
        RECT 140.990 41.660 141.980 42.140 ;
        RECT 141.000 40.860 141.990 41.340 ;
        RECT 135.820 39.420 136.770 39.700 ;
        RECT 95.580 36.400 104.840 36.500 ;
        RECT 78.770 34.950 79.760 35.430 ;
        RECT 95.500 35.670 104.860 36.400 ;
        RECT 126.860 37.370 127.870 37.740 ;
        RECT 140.990 40.080 141.980 40.560 ;
        RECT 140.980 39.280 141.970 39.760 ;
        RECT 135.830 37.090 136.740 37.450 ;
        RECT 140.990 38.500 141.980 38.980 ;
        RECT 140.990 37.700 141.980 38.180 ;
        RECT 78.760 34.140 79.750 34.620 ;
        RECT 78.760 33.320 79.720 33.760 ;
        RECT 54.960 28.560 55.960 30.370 ;
        RECT 66.615 29.635 67.210 30.230 ;
        RECT 64.290 28.820 64.810 29.340 ;
        RECT 73.570 32.950 74.550 33.210 ;
        RECT 73.580 30.620 74.540 30.940 ;
        RECT 73.570 28.360 74.540 28.630 ;
        RECT 55.540 25.470 55.800 26.470 ;
        RECT 57.840 25.470 58.120 26.470 ;
        RECT 60.120 25.470 60.400 26.470 ;
        RECT 62.410 25.470 62.690 26.470 ;
        RECT 64.710 25.470 64.990 26.470 ;
        RECT 73.590 26.100 74.540 26.360 ;
        RECT 55.560 23.840 64.950 24.420 ;
        RECT 55.390 11.400 64.190 18.240 ;
        RECT 74.330 11.280 83.680 18.120 ;
        RECT 124.260 35.140 125.170 35.440 ;
        RECT 126.920 35.090 127.820 35.440 ;
        RECT 140.990 36.910 141.980 37.390 ;
        RECT 126.990 34.290 128.020 34.710 ;
        RECT 124.190 30.620 124.640 32.680 ;
        RECT 126.120 30.640 126.540 32.630 ;
        RECT 135.810 34.710 136.770 35.220 ;
        RECT 141.000 36.120 141.990 36.600 ;
        RECT 140.990 35.330 141.980 35.810 ;
        RECT 141.000 34.550 141.990 35.030 ;
        RECT 140.990 33.740 141.980 34.220 ;
        RECT 140.990 32.920 141.950 33.360 ;
        RECT 117.190 28.160 118.190 29.970 ;
        RECT 128.845 29.235 129.440 29.830 ;
        RECT 126.520 28.420 127.040 28.940 ;
        RECT 135.800 32.550 136.780 32.810 ;
        RECT 135.810 30.220 136.770 30.540 ;
        RECT 135.800 27.960 136.770 28.230 ;
        RECT 117.770 25.070 118.030 26.070 ;
        RECT 120.070 25.070 120.350 26.070 ;
        RECT 122.350 25.070 122.630 26.070 ;
        RECT 124.640 25.070 124.920 26.070 ;
        RECT 126.940 25.070 127.220 26.070 ;
        RECT 135.820 25.700 136.770 25.960 ;
        RECT 117.790 23.440 127.180 24.020 ;
        RECT 94.640 11.670 105.730 18.200 ;
        RECT 117.320 13.120 127.600 18.610 ;
        RECT 135.980 13.520 146.160 18.400 ;
      LAYER met2 ;
        RECT 126.905 223.880 127.295 223.890 ;
        RECT 57.745 223.710 58.135 223.720 ;
        RECT 14.890 223.430 58.135 223.710 ;
        RECT 14.890 215.190 15.170 223.430 ;
        RECT 57.745 223.420 58.135 223.430 ;
        RECT 95.850 223.600 127.295 223.880 ;
        RECT 73.880 220.870 74.180 220.925 ;
        RECT 45.250 220.590 74.180 220.870 ;
        RECT 25.010 216.495 25.290 217.190 ;
        RECT 35.130 216.915 35.410 217.190 ;
        RECT 35.120 216.525 35.420 216.915 ;
        RECT 25.000 216.105 25.300 216.495 ;
        RECT 25.010 215.190 25.290 216.105 ;
        RECT 35.130 215.190 35.410 216.525 ;
        RECT 45.250 216.095 45.530 220.590 ;
        RECT 73.880 220.535 74.180 220.590 ;
        RECT 85.675 218.450 86.065 218.750 ;
        RECT 79.535 218.030 79.925 218.040 ;
        RECT 75.610 217.750 79.925 218.030 ;
        RECT 55.315 217.100 55.705 217.400 ;
        RECT 69.115 217.190 69.505 217.200 ;
        RECT 45.240 215.705 45.540 216.095 ;
        RECT 45.250 215.190 45.530 215.705 ;
        RECT 55.370 215.190 55.650 217.100 ;
        RECT 65.490 216.910 69.505 217.190 ;
        RECT 65.490 215.190 65.770 216.910 ;
        RECT 69.115 216.900 69.505 216.910 ;
        RECT 75.610 215.190 75.890 217.750 ;
        RECT 79.535 217.740 79.925 217.750 ;
        RECT 85.730 215.190 86.010 218.450 ;
        RECT 95.850 215.190 96.130 223.600 ;
        RECT 126.905 223.590 127.295 223.600 ;
        RECT 143.810 221.410 144.110 221.465 ;
        RECT 116.090 221.130 144.110 221.410 ;
        RECT 105.960 217.795 106.260 218.185 ;
        RECT 105.970 215.190 106.250 217.795 ;
        RECT 116.090 215.190 116.370 221.130 ;
        RECT 143.810 221.075 144.110 221.130 ;
        RECT 151.190 220.015 151.490 220.405 ;
        RECT 151.200 219.270 151.480 220.015 ;
        RECT 136.330 218.990 151.480 219.270 ;
        RECT 126.200 218.165 126.500 218.555 ;
        RECT 126.210 215.190 126.490 218.165 ;
        RECT 136.330 215.190 136.610 218.990 ;
        RECT 146.395 217.400 146.785 217.700 ;
        RECT 146.450 215.190 146.730 217.400 ;
        RECT 14.960 210.220 15.100 215.190 ;
        RECT 25.080 210.220 25.220 215.190 ;
        RECT 27.770 213.445 29.310 213.815 ;
        RECT 35.200 210.220 35.340 215.190 ;
        RECT 45.320 212.000 45.460 215.190 ;
        RECT 44.860 211.860 45.460 212.000 ;
        RECT 14.900 209.900 15.160 210.220 ;
        RECT 25.020 209.900 25.280 210.220 ;
        RECT 35.140 209.900 35.400 210.220 ;
        RECT 19.500 209.560 19.760 209.880 ;
        RECT 21.340 209.560 21.600 209.880 ;
        RECT 32.840 209.560 33.100 209.880 ;
        RECT 36.060 209.560 36.320 209.880 ;
        RECT 37.900 209.560 38.160 209.880 ;
        RECT 43.420 209.560 43.680 209.880 ;
        RECT 15.360 201.060 15.620 201.380 ;
        RECT 14.900 193.240 15.160 193.560 ;
        RECT 13.980 192.220 14.240 192.540 ;
        RECT 14.040 190.160 14.180 192.220 ;
        RECT 13.980 189.840 14.240 190.160 ;
        RECT 14.440 189.500 14.700 189.820 ;
        RECT 14.500 182.660 14.640 189.500 ;
        RECT 14.960 188.800 15.100 193.240 ;
        RECT 15.420 193.220 15.560 201.060 ;
        RECT 19.040 193.240 19.300 193.560 ;
        RECT 15.360 192.900 15.620 193.220 ;
        RECT 15.420 190.500 15.560 192.900 ;
        RECT 19.100 191.520 19.240 193.240 ;
        RECT 19.040 191.200 19.300 191.520 ;
        RECT 15.360 190.180 15.620 190.500 ;
        RECT 14.900 188.480 15.160 188.800 ;
        RECT 17.200 188.140 17.460 188.460 ;
        RECT 19.040 188.140 19.300 188.460 ;
        RECT 16.740 186.780 17.000 187.100 ;
        RECT 14.040 182.520 14.640 182.660 ;
        RECT 14.040 179.620 14.180 182.520 ;
        RECT 15.820 182.360 16.080 182.680 ;
        RECT 13.980 179.300 14.240 179.620 ;
        RECT 14.040 171.800 14.180 179.300 ;
        RECT 15.880 176.220 16.020 182.360 ;
        RECT 16.800 177.240 16.940 186.780 ;
        RECT 17.260 186.080 17.400 188.140 ;
        RECT 19.100 186.080 19.240 188.140 ;
        RECT 19.560 187.635 19.700 209.560 ;
        RECT 19.960 209.220 20.220 209.540 ;
        RECT 20.020 201.380 20.160 209.220 ;
        RECT 21.400 207.840 21.540 209.560 ;
        RECT 30.080 209.220 30.340 209.540 ;
        RECT 26.860 208.540 27.120 208.860 ;
        RECT 21.340 207.520 21.600 207.840 ;
        RECT 26.920 207.500 27.060 208.540 ;
        RECT 27.770 208.005 29.310 208.375 ;
        RECT 26.860 207.240 27.120 207.500 ;
        RECT 26.860 207.180 27.520 207.240 ;
        RECT 26.920 207.100 27.520 207.180 ;
        RECT 26.860 206.500 27.120 206.820 ;
        RECT 19.960 201.060 20.220 201.380 ;
        RECT 20.420 200.720 20.680 201.040 ;
        RECT 20.480 199.680 20.620 200.720 ;
        RECT 24.100 200.380 24.360 200.700 ;
        RECT 24.160 199.680 24.300 200.380 ;
        RECT 26.920 199.680 27.060 206.500 ;
        RECT 20.420 199.360 20.680 199.680 ;
        RECT 24.100 199.590 24.360 199.680 ;
        RECT 24.100 199.450 25.220 199.590 ;
        RECT 24.100 199.360 24.360 199.450 ;
        RECT 25.080 199.000 25.220 199.450 ;
        RECT 26.860 199.360 27.120 199.680 ;
        RECT 25.020 198.680 25.280 199.000 ;
        RECT 27.380 198.660 27.520 207.100 ;
        RECT 30.140 206.140 30.280 209.220 ;
        RECT 30.540 208.540 30.800 208.860 ;
        RECT 29.620 205.820 29.880 206.140 ;
        RECT 30.080 205.820 30.340 206.140 ;
        RECT 27.770 202.565 29.310 202.935 ;
        RECT 27.320 198.340 27.580 198.660 ;
        RECT 27.380 196.620 27.520 198.340 ;
        RECT 29.680 197.890 29.820 205.820 ;
        RECT 30.140 199.680 30.280 205.820 ;
        RECT 30.600 203.420 30.740 208.540 ;
        RECT 31.000 207.520 31.260 207.840 ;
        RECT 31.060 204.100 31.200 207.520 ;
        RECT 32.900 207.500 33.040 209.560 ;
        RECT 33.300 208.540 33.560 208.860 ;
        RECT 32.840 207.180 33.100 207.500 ;
        RECT 33.360 205.120 33.500 208.540 ;
        RECT 33.300 204.800 33.560 205.120 ;
        RECT 31.000 203.780 31.260 204.100 ;
        RECT 30.540 203.100 30.800 203.420 ;
        RECT 30.080 199.360 30.340 199.680 ;
        RECT 30.080 197.890 30.340 197.980 ;
        RECT 29.680 197.750 30.340 197.890 ;
        RECT 30.080 197.660 30.340 197.750 ;
        RECT 27.770 197.125 29.310 197.495 ;
        RECT 27.320 196.300 27.580 196.620 ;
        RECT 25.940 193.240 26.200 193.560 ;
        RECT 26.860 193.240 27.120 193.560 ;
        RECT 22.720 190.180 22.980 190.500 ;
        RECT 20.420 189.500 20.680 189.820 ;
        RECT 20.480 187.780 20.620 189.500 ;
        RECT 19.490 187.265 19.770 187.635 ;
        RECT 20.420 187.460 20.680 187.780 ;
        RECT 17.200 185.760 17.460 186.080 ;
        RECT 19.040 185.760 19.300 186.080 ;
        RECT 20.480 185.060 20.620 187.460 ;
        RECT 22.780 187.440 22.920 190.180 ;
        RECT 26.000 188.800 26.140 193.240 ;
        RECT 26.920 191.520 27.060 193.240 ;
        RECT 29.620 192.220 29.880 192.540 ;
        RECT 27.770 191.685 29.310 192.055 ;
        RECT 29.680 191.520 29.820 192.220 ;
        RECT 26.860 191.200 27.120 191.520 ;
        RECT 29.620 191.200 29.880 191.520 ;
        RECT 29.620 190.410 29.880 190.500 ;
        RECT 30.140 190.410 30.280 197.660 ;
        RECT 29.620 190.270 30.280 190.410 ;
        RECT 29.620 190.180 29.880 190.270 ;
        RECT 26.860 189.840 27.120 190.160 ;
        RECT 26.400 189.500 26.660 189.820 ;
        RECT 25.940 188.480 26.200 188.800 ;
        RECT 24.560 188.140 24.820 188.460 ;
        RECT 22.720 187.120 22.980 187.440 ;
        RECT 24.620 186.080 24.760 188.140 ;
        RECT 24.560 185.760 24.820 186.080 ;
        RECT 20.420 184.740 20.680 185.060 ;
        RECT 25.480 184.740 25.740 185.060 ;
        RECT 25.540 184.380 25.680 184.740 ;
        RECT 26.460 184.720 26.600 189.500 ;
        RECT 26.920 186.080 27.060 189.840 ;
        RECT 31.060 188.460 31.200 203.780 ;
        RECT 31.920 200.720 32.180 201.040 ;
        RECT 31.980 199.680 32.120 200.720 ;
        RECT 31.920 199.360 32.180 199.680 ;
        RECT 32.840 198.680 33.100 199.000 ;
        RECT 35.600 198.680 35.860 199.000 ;
        RECT 32.900 191.520 33.040 198.680 ;
        RECT 35.660 197.980 35.800 198.680 ;
        RECT 35.140 197.660 35.400 197.980 ;
        RECT 35.600 197.660 35.860 197.980 ;
        RECT 35.200 194.240 35.340 197.660 ;
        RECT 35.140 193.920 35.400 194.240 ;
        RECT 35.140 192.900 35.400 193.220 ;
        RECT 35.200 192.540 35.340 192.900 ;
        RECT 34.680 192.220 34.940 192.540 ;
        RECT 35.140 192.220 35.400 192.540 ;
        RECT 32.840 191.200 33.100 191.520 ;
        RECT 34.740 190.500 34.880 192.220 ;
        RECT 34.680 190.180 34.940 190.500 ;
        RECT 31.000 188.140 31.260 188.460 ;
        RECT 30.540 187.800 30.800 188.120 ;
        RECT 31.460 187.800 31.720 188.120 ;
        RECT 27.320 186.780 27.580 187.100 ;
        RECT 27.380 186.080 27.520 186.780 ;
        RECT 27.770 186.245 29.310 186.615 ;
        RECT 26.860 185.760 27.120 186.080 ;
        RECT 27.320 185.760 27.580 186.080 ;
        RECT 26.400 184.400 26.660 184.720 ;
        RECT 30.070 184.545 30.350 184.915 ;
        RECT 30.080 184.400 30.340 184.545 ;
        RECT 25.480 184.060 25.740 184.380 ;
        RECT 17.660 182.360 17.920 182.680 ;
        RECT 17.200 181.340 17.460 181.660 ;
        RECT 17.260 179.620 17.400 181.340 ;
        RECT 17.200 179.300 17.460 179.620 ;
        RECT 17.720 177.920 17.860 182.360 ;
        RECT 25.540 182.340 25.680 184.060 ;
        RECT 25.480 182.020 25.740 182.340 ;
        RECT 18.580 181.340 18.840 181.660 ;
        RECT 20.420 181.340 20.680 181.660 ;
        RECT 17.660 177.600 17.920 177.920 ;
        RECT 18.640 177.240 18.780 181.340 ;
        RECT 20.480 180.640 20.620 181.340 ;
        RECT 27.770 180.805 29.310 181.175 ;
        RECT 20.420 180.320 20.680 180.640 ;
        RECT 23.640 178.960 23.900 179.280 ;
        RECT 22.720 178.620 22.980 178.940 ;
        RECT 22.780 177.240 22.920 178.620 ;
        RECT 23.700 177.920 23.840 178.960 ;
        RECT 25.020 178.620 25.280 178.940 ;
        RECT 23.640 177.600 23.900 177.920 ;
        RECT 16.740 176.920 17.000 177.240 ;
        RECT 18.580 176.920 18.840 177.240 ;
        RECT 22.720 176.920 22.980 177.240 ;
        RECT 15.820 175.900 16.080 176.220 ;
        RECT 13.980 171.480 14.240 171.800 ;
        RECT 15.880 170.780 16.020 175.900 ;
        RECT 16.280 173.180 16.540 173.500 ;
        RECT 16.340 172.140 16.480 173.180 ;
        RECT 16.280 171.820 16.540 172.140 ;
        RECT 15.820 170.460 16.080 170.780 ;
        RECT 15.880 169.420 16.020 170.460 ;
        RECT 16.800 169.760 16.940 176.920 ;
        RECT 25.080 176.560 25.220 178.620 ;
        RECT 25.020 176.240 25.280 176.560 ;
        RECT 26.860 175.900 27.120 176.220 ;
        RECT 18.120 173.860 18.380 174.180 ;
        RECT 18.180 169.760 18.320 173.860 ;
        RECT 26.400 171.820 26.660 172.140 ;
        RECT 22.720 170.460 22.980 170.780 ;
        RECT 16.740 169.440 17.000 169.760 ;
        RECT 18.120 169.440 18.380 169.760 ;
        RECT 15.820 169.100 16.080 169.420 ;
        RECT 22.780 168.400 22.920 170.460 ;
        RECT 26.460 169.275 26.600 171.820 ;
        RECT 26.920 169.760 27.060 175.900 ;
        RECT 27.770 175.365 29.310 175.735 ;
        RECT 27.320 170.800 27.580 171.120 ;
        RECT 26.860 169.440 27.120 169.760 ;
        RECT 26.390 168.905 26.670 169.275 ;
        RECT 26.400 168.760 26.660 168.905 ;
        RECT 22.720 168.080 22.980 168.400 ;
        RECT 19.040 167.740 19.300 168.060 ;
        RECT 19.100 163.300 19.240 167.740 ;
        RECT 26.460 166.360 26.600 168.760 ;
        RECT 27.380 168.740 27.520 170.800 ;
        RECT 27.770 169.925 29.310 170.295 ;
        RECT 27.320 168.420 27.580 168.740 ;
        RECT 28.240 168.420 28.500 168.740 ;
        RECT 28.300 167.040 28.440 168.420 ;
        RECT 28.240 166.720 28.500 167.040 ;
        RECT 26.400 166.040 26.660 166.360 ;
        RECT 26.460 164.320 26.600 166.040 ;
        RECT 27.770 164.485 29.310 164.855 ;
        RECT 26.400 164.000 26.660 164.320 ;
        RECT 16.280 162.980 16.540 163.300 ;
        RECT 19.040 162.980 19.300 163.300 ;
        RECT 16.340 160.580 16.480 162.980 ;
        RECT 26.860 160.600 27.120 160.920 ;
        RECT 16.280 160.260 16.540 160.580 ;
        RECT 16.340 152.420 16.480 160.260 ;
        RECT 26.920 158.880 27.060 160.600 ;
        RECT 27.770 159.045 29.310 159.415 ;
        RECT 26.860 158.560 27.120 158.880 ;
        RECT 25.020 157.540 25.280 157.860 ;
        RECT 25.480 157.540 25.740 157.860 ;
        RECT 19.040 155.160 19.300 155.480 ;
        RECT 17.200 154.140 17.460 154.460 ;
        RECT 17.260 152.420 17.400 154.140 ;
        RECT 16.280 152.100 16.540 152.420 ;
        RECT 17.200 152.100 17.460 152.420 ;
        RECT 16.340 139.500 16.480 152.100 ;
        RECT 19.100 150.720 19.240 155.160 ;
        RECT 24.560 152.440 24.820 152.760 ;
        RECT 19.040 150.400 19.300 150.720 ;
        RECT 20.420 149.380 20.680 149.700 ;
        RECT 18.580 141.220 18.840 141.540 ;
        RECT 17.200 140.540 17.460 140.860 ;
        RECT 16.280 139.180 16.540 139.500 ;
        RECT 17.260 139.160 17.400 140.540 ;
        RECT 17.200 138.840 17.460 139.160 ;
        RECT 18.640 137.120 18.780 141.220 ;
        RECT 18.580 136.800 18.840 137.120 ;
        RECT 20.480 136.100 20.620 149.380 ;
        RECT 24.100 147.340 24.360 147.660 ;
        RECT 23.640 146.660 23.900 146.980 ;
        RECT 23.700 139.500 23.840 146.660 ;
        RECT 24.160 145.280 24.300 147.340 ;
        RECT 24.100 144.960 24.360 145.280 ;
        RECT 24.620 144.260 24.760 152.440 ;
        RECT 25.080 149.020 25.220 157.540 ;
        RECT 25.540 156.160 25.680 157.540 ;
        RECT 25.480 155.840 25.740 156.160 ;
        RECT 27.770 153.605 29.310 153.975 ;
        RECT 27.320 152.100 27.580 152.420 ;
        RECT 27.380 149.360 27.520 152.100 ;
        RECT 29.620 151.420 29.880 151.740 ;
        RECT 29.680 150.720 29.820 151.420 ;
        RECT 29.620 150.400 29.880 150.720 ;
        RECT 27.320 149.040 27.580 149.360 ;
        RECT 25.020 148.700 25.280 149.020 ;
        RECT 27.380 147.400 27.520 149.040 ;
        RECT 27.770 148.165 29.310 148.535 ;
        RECT 27.380 147.260 27.980 147.400 ;
        RECT 27.840 146.980 27.980 147.260 ;
        RECT 26.860 146.660 27.120 146.980 ;
        RECT 27.780 146.660 28.040 146.980 ;
        RECT 25.480 145.980 25.740 146.300 ;
        RECT 25.540 145.280 25.680 145.980 ;
        RECT 25.480 144.960 25.740 145.280 ;
        RECT 26.920 144.680 27.060 146.660 ;
        RECT 26.920 144.600 27.520 144.680 ;
        RECT 26.920 144.540 27.580 144.600 ;
        RECT 27.320 144.280 27.580 144.540 ;
        RECT 24.560 143.940 24.820 144.260 ;
        RECT 24.560 140.880 24.820 141.200 ;
        RECT 23.640 139.180 23.900 139.500 ;
        RECT 24.620 138.820 24.760 140.880 ;
        RECT 24.560 138.500 24.820 138.820 ;
        RECT 27.380 138.480 27.520 144.280 ;
        RECT 27.770 142.725 29.310 143.095 ;
        RECT 28.700 141.220 28.960 141.540 ;
        RECT 28.760 139.500 28.900 141.220 ;
        RECT 29.160 140.540 29.420 140.860 ;
        RECT 29.220 139.500 29.360 140.540 ;
        RECT 28.700 139.180 28.960 139.500 ;
        RECT 29.160 139.180 29.420 139.500 ;
        RECT 25.940 138.160 26.200 138.480 ;
        RECT 27.320 138.160 27.580 138.480 ;
        RECT 25.480 137.820 25.740 138.140 ;
        RECT 25.540 137.120 25.680 137.820 ;
        RECT 26.000 137.120 26.140 138.160 ;
        RECT 27.770 137.285 29.310 137.655 ;
        RECT 25.480 136.800 25.740 137.120 ;
        RECT 25.940 136.800 26.200 137.120 ;
        RECT 20.420 135.780 20.680 136.100 ;
        RECT 27.320 135.780 27.580 136.100 ;
        RECT 27.380 134.360 27.520 135.780 ;
        RECT 30.140 134.360 30.280 184.400 ;
        RECT 30.600 183.020 30.740 187.800 ;
        RECT 31.000 186.780 31.260 187.100 ;
        RECT 31.060 186.080 31.200 186.780 ;
        RECT 31.000 185.760 31.260 186.080 ;
        RECT 31.520 184.380 31.660 187.800 ;
        RECT 32.840 184.740 33.100 185.060 ;
        RECT 31.460 184.060 31.720 184.380 ;
        RECT 32.900 183.360 33.040 184.740 ;
        RECT 32.840 183.040 33.100 183.360 ;
        RECT 30.540 182.700 30.800 183.020 ;
        RECT 34.220 179.980 34.480 180.300 ;
        RECT 32.380 178.620 32.640 178.940 ;
        RECT 32.440 177.240 32.580 178.620 ;
        RECT 32.380 176.920 32.640 177.240 ;
        RECT 33.300 176.920 33.560 177.240 ;
        RECT 32.440 171.800 32.580 176.920 ;
        RECT 33.360 173.500 33.500 176.920 ;
        RECT 33.760 176.580 34.020 176.900 ;
        RECT 33.300 173.180 33.560 173.500 ;
        RECT 32.380 171.480 32.640 171.800 ;
        RECT 30.540 170.460 30.800 170.780 ;
        RECT 31.000 170.460 31.260 170.780 ;
        RECT 30.600 169.760 30.740 170.460 ;
        RECT 30.540 169.440 30.800 169.760 ;
        RECT 31.060 167.040 31.200 170.460 ;
        RECT 31.000 166.720 31.260 167.040 ;
        RECT 31.920 165.360 32.180 165.680 ;
        RECT 30.540 163.320 30.800 163.640 ;
        RECT 31.460 163.320 31.720 163.640 ;
        RECT 30.600 153.100 30.740 163.320 ;
        RECT 31.520 159.900 31.660 163.320 ;
        RECT 31.460 159.580 31.720 159.900 ;
        RECT 31.520 155.820 31.660 159.580 ;
        RECT 31.460 155.500 31.720 155.820 ;
        RECT 31.980 155.480 32.120 165.360 ;
        RECT 32.440 156.160 32.580 171.480 ;
        RECT 33.360 171.460 33.500 173.180 ;
        RECT 33.820 171.460 33.960 176.580 ;
        RECT 33.300 171.140 33.560 171.460 ;
        RECT 33.760 171.140 34.020 171.460 ;
        RECT 33.820 168.400 33.960 171.140 ;
        RECT 32.840 168.080 33.100 168.400 ;
        RECT 33.760 168.080 34.020 168.400 ;
        RECT 32.900 167.040 33.040 168.080 ;
        RECT 32.840 166.720 33.100 167.040 ;
        RECT 32.840 165.020 33.100 165.340 ;
        RECT 32.380 155.840 32.640 156.160 ;
        RECT 31.000 155.160 31.260 155.480 ;
        RECT 31.920 155.160 32.180 155.480 ;
        RECT 31.060 153.440 31.200 155.160 ;
        RECT 31.980 154.880 32.120 155.160 ;
        RECT 31.980 154.740 32.580 154.880 ;
        RECT 31.920 154.140 32.180 154.460 ;
        RECT 31.000 153.120 31.260 153.440 ;
        RECT 30.540 152.780 30.800 153.100 ;
        RECT 30.600 148.000 30.740 152.780 ;
        RECT 31.460 151.760 31.720 152.080 ;
        RECT 31.000 149.720 31.260 150.040 ;
        RECT 30.540 147.680 30.800 148.000 ;
        RECT 31.060 146.980 31.200 149.720 ;
        RECT 31.000 146.660 31.260 146.980 ;
        RECT 31.060 141.540 31.200 146.660 ;
        RECT 31.520 144.260 31.660 151.760 ;
        RECT 31.980 151.740 32.120 154.140 ;
        RECT 32.440 152.420 32.580 154.740 ;
        RECT 32.380 152.100 32.640 152.420 ;
        RECT 31.920 151.420 32.180 151.740 ;
        RECT 31.460 143.940 31.720 144.260 ;
        RECT 31.000 141.220 31.260 141.540 ;
        RECT 31.980 140.860 32.120 151.420 ;
        RECT 32.440 141.540 32.580 152.100 ;
        RECT 32.380 141.220 32.640 141.540 ;
        RECT 31.000 140.540 31.260 140.860 ;
        RECT 31.920 140.540 32.180 140.860 ;
        RECT 31.060 139.160 31.200 140.540 ;
        RECT 32.900 139.160 33.040 165.020 ;
        RECT 33.820 163.300 33.960 168.080 ;
        RECT 33.760 162.980 34.020 163.300 ;
        RECT 34.280 156.070 34.420 179.980 ;
        RECT 34.740 177.920 34.880 190.180 ;
        RECT 35.200 188.120 35.340 192.220 ;
        RECT 35.140 187.800 35.400 188.120 ;
        RECT 35.140 184.915 35.400 185.060 ;
        RECT 35.130 184.545 35.410 184.915 ;
        RECT 35.140 182.700 35.400 183.020 ;
        RECT 35.200 180.300 35.340 182.700 ;
        RECT 36.120 182.660 36.260 209.560 ;
        RECT 37.960 204.100 38.100 209.560 ;
        RECT 38.820 209.220 39.080 209.540 ;
        RECT 38.360 208.540 38.620 208.860 ;
        RECT 38.420 206.820 38.560 208.540 ;
        RECT 38.360 206.500 38.620 206.820 ;
        RECT 38.880 205.120 39.020 209.220 ;
        RECT 42.960 208.880 43.220 209.200 ;
        RECT 39.740 206.500 40.000 206.820 ;
        RECT 38.820 204.800 39.080 205.120 ;
        RECT 37.900 203.780 38.160 204.100 ;
        RECT 38.360 202.080 38.620 202.400 ;
        RECT 38.420 200.700 38.560 202.080 ;
        RECT 39.800 201.380 39.940 206.500 ;
        RECT 42.500 204.120 42.760 204.440 ;
        RECT 41.120 203.780 41.380 204.100 ;
        RECT 40.200 203.440 40.460 203.760 ;
        RECT 39.740 201.060 40.000 201.380 ;
        RECT 38.360 200.380 38.620 200.700 ;
        RECT 37.900 195.280 38.160 195.600 ;
        RECT 37.960 193.220 38.100 195.280 ;
        RECT 37.900 192.900 38.160 193.220 ;
        RECT 38.420 192.960 38.560 200.380 ;
        RECT 38.420 192.880 39.480 192.960 ;
        RECT 38.420 192.820 39.540 192.880 ;
        RECT 38.420 192.540 38.560 192.820 ;
        RECT 39.280 192.560 39.540 192.820 ;
        RECT 37.440 192.220 37.700 192.540 ;
        RECT 38.360 192.220 38.620 192.540 ;
        RECT 38.820 192.220 39.080 192.540 ;
        RECT 37.500 191.520 37.640 192.220 ;
        RECT 38.880 191.520 39.020 192.220 ;
        RECT 37.440 191.200 37.700 191.520 ;
        RECT 38.820 191.200 39.080 191.520 ;
        RECT 39.340 186.080 39.480 192.560 ;
        RECT 38.360 185.760 38.620 186.080 ;
        RECT 39.280 185.760 39.540 186.080 ;
        RECT 38.420 184.380 38.560 185.760 ;
        RECT 37.440 184.060 37.700 184.380 ;
        RECT 38.360 184.290 38.620 184.380 ;
        RECT 37.960 184.150 38.620 184.290 ;
        RECT 37.500 183.360 37.640 184.060 ;
        RECT 37.440 183.040 37.700 183.360 ;
        RECT 36.120 182.520 37.180 182.660 ;
        RECT 35.140 179.980 35.400 180.300 ;
        RECT 36.060 179.640 36.320 179.960 ;
        RECT 35.140 179.300 35.400 179.620 ;
        RECT 34.680 177.600 34.940 177.920 ;
        RECT 35.200 173.840 35.340 179.300 ;
        RECT 36.120 177.920 36.260 179.640 ;
        RECT 36.060 177.600 36.320 177.920 ;
        RECT 35.600 176.920 35.860 177.240 ;
        RECT 35.140 173.520 35.400 173.840 ;
        RECT 35.660 168.740 35.800 176.920 ;
        RECT 36.060 176.580 36.320 176.900 ;
        RECT 36.120 170.780 36.260 176.580 ;
        RECT 36.520 175.900 36.780 176.220 ;
        RECT 36.580 174.180 36.720 175.900 ;
        RECT 37.040 174.715 37.180 182.520 ;
        RECT 37.440 178.960 37.700 179.280 ;
        RECT 37.500 175.200 37.640 178.960 ;
        RECT 37.440 174.880 37.700 175.200 ;
        RECT 36.970 174.345 37.250 174.715 ;
        RECT 36.520 173.860 36.780 174.180 ;
        RECT 36.980 173.520 37.240 173.840 ;
        RECT 37.040 171.460 37.180 173.520 ;
        RECT 36.980 171.140 37.240 171.460 ;
        RECT 36.060 170.460 36.320 170.780 ;
        RECT 37.040 169.760 37.180 171.140 ;
        RECT 36.980 169.440 37.240 169.760 ;
        RECT 35.600 168.420 35.860 168.740 ;
        RECT 35.600 166.720 35.860 167.040 ;
        RECT 35.660 165.340 35.800 166.720 ;
        RECT 35.600 165.020 35.860 165.340 ;
        RECT 37.960 164.320 38.100 184.150 ;
        RECT 38.360 184.060 38.620 184.150 ;
        RECT 39.800 177.240 39.940 201.060 ;
        RECT 40.260 200.700 40.400 203.440 ;
        RECT 41.180 202.400 41.320 203.780 ;
        RECT 41.120 202.080 41.380 202.400 ;
        RECT 42.040 201.740 42.300 202.060 ;
        RECT 40.200 200.380 40.460 200.700 ;
        RECT 41.580 198.340 41.840 198.660 ;
        RECT 41.640 196.960 41.780 198.340 ;
        RECT 41.580 196.640 41.840 196.960 ;
        RECT 40.200 193.240 40.460 193.560 ;
        RECT 40.260 185.400 40.400 193.240 ;
        RECT 40.660 192.220 40.920 192.540 ;
        RECT 40.720 190.500 40.860 192.220 ;
        RECT 40.660 190.180 40.920 190.500 ;
        RECT 41.580 187.800 41.840 188.120 ;
        RECT 41.120 185.420 41.380 185.740 ;
        RECT 40.200 185.080 40.460 185.400 ;
        RECT 40.660 185.080 40.920 185.400 ;
        RECT 40.720 183.360 40.860 185.080 ;
        RECT 40.660 183.040 40.920 183.360 ;
        RECT 40.660 181.680 40.920 182.000 ;
        RECT 39.740 176.920 40.000 177.240 ;
        RECT 38.820 176.240 39.080 176.560 ;
        RECT 38.360 175.900 38.620 176.220 ;
        RECT 38.420 174.180 38.560 175.900 ;
        RECT 38.880 174.520 39.020 176.240 ;
        RECT 38.820 174.200 39.080 174.520 ;
        RECT 38.360 173.860 38.620 174.180 ;
        RECT 38.820 173.180 39.080 173.500 ;
        RECT 38.880 168.060 39.020 173.180 ;
        RECT 39.280 171.480 39.540 171.800 ;
        RECT 39.340 169.275 39.480 171.480 ;
        RECT 40.720 170.780 40.860 181.680 ;
        RECT 40.660 170.460 40.920 170.780 ;
        RECT 40.720 169.760 40.860 170.460 ;
        RECT 40.660 169.440 40.920 169.760 ;
        RECT 39.270 168.905 39.550 169.275 ;
        RECT 39.280 168.760 39.540 168.905 ;
        RECT 38.820 167.740 39.080 168.060 ;
        RECT 37.900 164.000 38.160 164.320 ;
        RECT 41.180 163.300 41.320 185.420 ;
        RECT 41.640 184.630 41.780 187.800 ;
        RECT 42.100 187.780 42.240 201.740 ;
        RECT 42.560 201.040 42.700 204.120 ;
        RECT 42.500 200.720 42.760 201.040 ;
        RECT 42.040 187.460 42.300 187.780 ;
        RECT 43.020 186.080 43.160 208.880 ;
        RECT 43.480 202.060 43.620 209.560 ;
        RECT 44.860 209.200 45.000 211.860 ;
        RECT 45.190 210.725 46.730 211.095 ;
        RECT 48.020 209.560 48.280 209.880 ;
        RECT 53.080 209.560 53.340 209.880 ;
        RECT 47.560 209.220 47.820 209.540 ;
        RECT 44.800 208.880 45.060 209.200 ;
        RECT 45.720 208.540 45.980 208.860 ;
        RECT 44.800 206.160 45.060 206.480 ;
        RECT 44.860 205.120 45.000 206.160 ;
        RECT 45.780 206.140 45.920 208.540 ;
        RECT 47.620 207.840 47.760 209.220 ;
        RECT 47.560 207.520 47.820 207.840 ;
        RECT 47.100 207.180 47.360 207.500 ;
        RECT 45.720 205.820 45.980 206.140 ;
        RECT 45.190 205.285 46.730 205.655 ;
        RECT 47.160 205.120 47.300 207.180 ;
        RECT 44.800 204.800 45.060 205.120 ;
        RECT 46.180 204.800 46.440 205.120 ;
        RECT 47.100 204.800 47.360 205.120 ;
        RECT 46.240 204.440 46.380 204.800 ;
        RECT 46.180 204.120 46.440 204.440 ;
        RECT 47.560 204.350 47.820 204.440 ;
        RECT 48.080 204.350 48.220 209.560 ;
        RECT 52.160 206.730 52.420 206.820 ;
        RECT 47.560 204.210 48.220 204.350 ;
        RECT 47.560 204.120 47.820 204.210 ;
        RECT 48.080 202.400 48.220 204.210 ;
        RECT 51.300 206.590 52.420 206.730 ;
        RECT 48.020 202.080 48.280 202.400 ;
        RECT 43.420 201.740 43.680 202.060 ;
        RECT 43.480 196.960 43.620 201.740 ;
        RECT 48.020 201.060 48.280 201.380 ;
        RECT 47.100 200.720 47.360 201.040 ;
        RECT 45.190 199.845 46.730 200.215 ;
        RECT 43.420 196.640 43.680 196.960 ;
        RECT 44.800 194.940 45.060 195.260 ;
        RECT 44.860 192.880 45.000 194.940 ;
        RECT 45.190 194.405 46.730 194.775 ;
        RECT 47.160 194.240 47.300 200.720 ;
        RECT 48.080 199.680 48.220 201.060 ;
        RECT 48.020 199.360 48.280 199.680 ;
        RECT 49.860 198.680 50.120 199.000 ;
        RECT 47.100 193.920 47.360 194.240 ;
        RECT 47.100 193.470 47.360 193.560 ;
        RECT 47.100 193.330 47.760 193.470 ;
        RECT 47.100 193.240 47.360 193.330 ;
        RECT 44.800 192.560 45.060 192.880 ;
        RECT 44.860 191.520 45.000 192.560 ;
        RECT 47.100 192.220 47.360 192.540 ;
        RECT 44.800 191.200 45.060 191.520 ;
        RECT 45.190 188.965 46.730 189.335 ;
        RECT 42.960 185.760 43.220 186.080 ;
        RECT 47.160 184.720 47.300 192.220 ;
        RECT 47.620 190.160 47.760 193.330 ;
        RECT 47.560 189.840 47.820 190.160 ;
        RECT 47.620 188.120 47.760 189.840 ;
        RECT 47.560 187.800 47.820 188.120 ;
        RECT 49.920 187.780 50.060 198.680 ;
        RECT 49.860 187.460 50.120 187.780 ;
        RECT 48.480 184.740 48.740 185.060 ;
        RECT 42.040 184.630 42.300 184.720 ;
        RECT 41.640 184.490 42.300 184.630 ;
        RECT 41.640 181.660 41.780 184.490 ;
        RECT 42.040 184.400 42.300 184.490 ;
        RECT 47.100 184.400 47.360 184.720 ;
        RECT 45.190 183.525 46.730 183.895 ;
        RECT 42.040 182.360 42.300 182.680 ;
        RECT 41.580 181.340 41.840 181.660 ;
        RECT 41.640 170.780 41.780 181.340 ;
        RECT 42.100 178.940 42.240 182.360 ;
        RECT 47.090 181.825 47.370 182.195 ;
        RECT 42.960 180.320 43.220 180.640 ;
        RECT 42.040 178.620 42.300 178.940 ;
        RECT 42.100 174.860 42.240 178.620 ;
        RECT 42.500 174.880 42.760 175.200 ;
        RECT 42.040 174.540 42.300 174.860 ;
        RECT 42.040 173.520 42.300 173.840 ;
        RECT 42.100 171.800 42.240 173.520 ;
        RECT 42.040 171.480 42.300 171.800 ;
        RECT 41.580 170.460 41.840 170.780 ;
        RECT 41.640 168.060 41.780 170.460 ;
        RECT 41.580 167.740 41.840 168.060 ;
        RECT 42.100 166.360 42.240 171.480 ;
        RECT 42.560 168.740 42.700 174.880 ;
        RECT 43.020 174.180 43.160 180.320 ;
        RECT 47.160 179.620 47.300 181.825 ;
        RECT 48.540 179.960 48.680 184.740 ;
        RECT 49.860 184.400 50.120 184.720 ;
        RECT 49.920 181.660 50.060 184.400 ;
        RECT 50.780 182.360 51.040 182.680 ;
        RECT 49.860 181.340 50.120 181.660 ;
        RECT 49.920 180.640 50.060 181.340 ;
        RECT 49.860 180.320 50.120 180.640 ;
        RECT 48.480 179.640 48.740 179.960 ;
        RECT 43.420 179.300 43.680 179.620 ;
        RECT 43.880 179.300 44.140 179.620 ;
        RECT 47.100 179.300 47.360 179.620 ;
        RECT 50.320 179.300 50.580 179.620 ;
        RECT 42.960 173.860 43.220 174.180 ;
        RECT 43.480 173.500 43.620 179.300 ;
        RECT 43.940 174.180 44.080 179.300 ;
        RECT 45.190 178.085 46.730 178.455 ;
        RECT 49.400 176.920 49.660 177.240 ;
        RECT 44.340 174.200 44.600 174.520 ;
        RECT 44.800 174.200 45.060 174.520 ;
        RECT 43.880 173.860 44.140 174.180 ;
        RECT 43.420 173.180 43.680 173.500 ;
        RECT 43.940 172.560 44.080 173.860 ;
        RECT 44.400 173.500 44.540 174.200 ;
        RECT 44.340 173.180 44.600 173.500 ;
        RECT 43.480 172.480 44.080 172.560 ;
        RECT 43.420 172.420 44.080 172.480 ;
        RECT 43.420 172.160 43.680 172.420 ;
        RECT 42.960 171.480 43.220 171.800 ;
        RECT 43.020 169.760 43.160 171.480 ;
        RECT 44.860 171.460 45.000 174.200 ;
        RECT 45.190 172.645 46.730 173.015 ;
        RECT 45.260 171.820 45.520 172.140 ;
        RECT 44.800 171.140 45.060 171.460 ;
        RECT 42.960 169.440 43.220 169.760 ;
        RECT 45.320 169.420 45.460 171.820 ;
        RECT 48.940 171.480 49.200 171.800 ;
        RECT 48.480 170.460 48.740 170.780 ;
        RECT 45.260 169.100 45.520 169.420 ;
        RECT 48.540 169.080 48.680 170.460 ;
        RECT 49.000 169.760 49.140 171.480 ;
        RECT 49.460 169.760 49.600 176.920 ;
        RECT 50.380 174.520 50.520 179.300 ;
        RECT 50.840 174.520 50.980 182.360 ;
        RECT 50.320 174.200 50.580 174.520 ;
        RECT 50.780 174.200 51.040 174.520 ;
        RECT 51.300 172.140 51.440 206.590 ;
        RECT 52.160 206.500 52.420 206.590 ;
        RECT 51.700 201.060 51.960 201.380 ;
        RECT 51.760 199.680 51.900 201.060 ;
        RECT 52.160 200.380 52.420 200.700 ;
        RECT 52.220 199.680 52.360 200.380 ;
        RECT 53.140 199.680 53.280 209.560 ;
        RECT 55.440 207.840 55.580 215.190 ;
        RECT 62.615 213.445 64.155 213.815 ;
        RECT 65.560 213.280 65.700 215.190 ;
        RECT 65.500 212.960 65.760 213.280 ;
        RECT 64.120 211.940 64.380 212.260 ;
        RECT 55.840 209.560 56.100 209.880 ;
        RECT 58.140 209.560 58.400 209.880 ;
        RECT 55.380 207.520 55.640 207.840 ;
        RECT 51.700 199.360 51.960 199.680 ;
        RECT 52.160 199.360 52.420 199.680 ;
        RECT 53.080 199.360 53.340 199.680 ;
        RECT 51.700 198.340 51.960 198.660 ;
        RECT 51.760 194.240 51.900 198.340 ;
        RECT 55.900 195.940 56.040 209.560 ;
        RECT 56.300 197.660 56.560 197.980 ;
        RECT 56.360 195.940 56.500 197.660 ;
        RECT 57.680 196.640 57.940 196.960 ;
        RECT 55.840 195.620 56.100 195.940 ;
        RECT 56.300 195.620 56.560 195.940 ;
        RECT 51.700 193.920 51.960 194.240 ;
        RECT 54.460 193.920 54.720 194.240 ;
        RECT 53.540 192.220 53.800 192.540 ;
        RECT 53.600 191.520 53.740 192.220 ;
        RECT 53.540 191.200 53.800 191.520 ;
        RECT 54.000 191.200 54.260 191.520 ;
        RECT 54.060 190.920 54.200 191.200 ;
        RECT 54.520 191.180 54.660 193.920 ;
        RECT 52.680 190.780 54.200 190.920 ;
        RECT 54.460 190.860 54.720 191.180 ;
        RECT 52.680 189.820 52.820 190.780 ;
        RECT 54.520 190.500 54.660 190.860 ;
        RECT 53.540 190.180 53.800 190.500 ;
        RECT 54.460 190.180 54.720 190.500 ;
        RECT 55.380 190.180 55.640 190.500 ;
        RECT 52.620 189.500 52.880 189.820 ;
        RECT 53.080 189.500 53.340 189.820 ;
        RECT 52.160 188.140 52.420 188.460 ;
        RECT 51.700 187.800 51.960 188.120 ;
        RECT 51.760 182.660 51.900 187.800 ;
        RECT 52.220 185.990 52.360 188.140 ;
        RECT 53.140 187.100 53.280 189.500 ;
        RECT 53.600 188.460 53.740 190.180 ;
        RECT 53.540 188.140 53.800 188.460 ;
        RECT 53.080 186.780 53.340 187.100 ;
        RECT 53.080 185.990 53.340 186.080 ;
        RECT 52.220 185.850 53.340 185.990 ;
        RECT 53.080 185.760 53.340 185.850 ;
        RECT 52.160 185.080 52.420 185.400 ;
        RECT 52.220 184.380 52.360 185.080 ;
        RECT 52.160 184.060 52.420 184.380 ;
        RECT 53.080 184.060 53.340 184.380 ;
        RECT 53.140 183.360 53.280 184.060 ;
        RECT 53.080 183.040 53.340 183.360 ;
        RECT 54.520 182.660 54.660 190.180 ;
        RECT 55.440 188.800 55.580 190.180 ;
        RECT 55.380 188.480 55.640 188.800 ;
        RECT 55.900 188.120 56.040 195.620 ;
        RECT 56.360 192.880 56.500 195.620 ;
        RECT 56.300 192.560 56.560 192.880 ;
        RECT 57.220 192.220 57.480 192.540 ;
        RECT 57.280 190.840 57.420 192.220 ;
        RECT 57.220 190.520 57.480 190.840 ;
        RECT 56.760 189.500 57.020 189.820 ;
        RECT 56.820 188.460 56.960 189.500 ;
        RECT 56.760 188.140 57.020 188.460 ;
        RECT 55.840 187.800 56.100 188.120 ;
        RECT 51.760 182.520 52.360 182.660 ;
        RECT 51.700 181.340 51.960 181.660 ;
        RECT 51.760 179.620 51.900 181.340 ;
        RECT 51.700 179.300 51.960 179.620 ;
        RECT 51.240 171.820 51.500 172.140 ;
        RECT 48.940 169.440 49.200 169.760 ;
        RECT 49.400 169.440 49.660 169.760 ;
        RECT 48.480 168.760 48.740 169.080 ;
        RECT 42.500 168.420 42.760 168.740 ;
        RECT 45.190 167.205 46.730 167.575 ;
        RECT 42.040 166.040 42.300 166.360 ;
        RECT 43.880 165.700 44.140 166.020 ;
        RECT 43.420 165.020 43.680 165.340 ;
        RECT 43.480 163.300 43.620 165.020 ;
        RECT 39.740 162.980 40.000 163.300 ;
        RECT 41.120 162.980 41.380 163.300 ;
        RECT 43.420 163.210 43.680 163.300 ;
        RECT 43.020 163.070 43.680 163.210 ;
        RECT 37.440 162.640 37.700 162.960 ;
        RECT 37.500 160.920 37.640 162.640 ;
        RECT 38.360 162.300 38.620 162.620 ;
        RECT 37.440 160.600 37.700 160.920 ;
        RECT 33.820 155.930 34.420 156.070 ;
        RECT 33.820 141.200 33.960 155.930 ;
        RECT 34.220 155.160 34.480 155.480 ;
        RECT 34.280 149.700 34.420 155.160 ;
        RECT 38.420 155.140 38.560 162.300 ;
        RECT 38.820 160.600 39.080 160.920 ;
        RECT 35.140 154.820 35.400 155.140 ;
        RECT 38.360 154.820 38.620 155.140 ;
        RECT 35.200 152.420 35.340 154.820 ;
        RECT 38.880 154.800 39.020 160.600 ;
        RECT 39.800 159.900 39.940 162.980 ;
        RECT 41.180 160.920 41.320 162.980 ;
        RECT 41.120 160.600 41.380 160.920 ;
        RECT 39.740 159.580 40.000 159.900 ;
        RECT 42.040 157.200 42.300 157.520 ;
        RECT 41.120 156.860 41.380 157.180 ;
        RECT 39.740 155.730 40.000 155.820 ;
        RECT 39.740 155.590 40.860 155.730 ;
        RECT 39.740 155.500 40.000 155.590 ;
        RECT 39.280 155.160 39.540 155.480 ;
        RECT 39.340 154.880 39.480 155.160 ;
        RECT 39.340 154.800 40.400 154.880 ;
        RECT 38.820 154.480 39.080 154.800 ;
        RECT 39.340 154.740 40.460 154.800 ;
        RECT 40.200 154.480 40.460 154.740 ;
        RECT 35.140 152.100 35.400 152.420 ;
        RECT 40.200 152.100 40.460 152.420 ;
        RECT 36.980 151.760 37.240 152.080 ;
        RECT 38.820 151.760 39.080 152.080 ;
        RECT 35.600 149.720 35.860 150.040 ;
        RECT 34.220 149.380 34.480 149.700 ;
        RECT 34.280 146.980 34.420 149.380 ;
        RECT 34.220 146.660 34.480 146.980 ;
        RECT 35.660 144.940 35.800 149.720 ;
        RECT 35.600 144.620 35.860 144.940 ;
        RECT 37.040 141.540 37.180 151.760 ;
        RECT 38.880 150.040 39.020 151.760 ;
        RECT 40.260 150.040 40.400 152.100 ;
        RECT 40.720 150.720 40.860 155.590 ;
        RECT 41.180 155.140 41.320 156.860 ;
        RECT 42.100 155.480 42.240 157.200 ;
        RECT 42.500 155.840 42.760 156.160 ;
        RECT 42.040 155.160 42.300 155.480 ;
        RECT 41.120 154.820 41.380 155.140 ;
        RECT 41.180 152.080 41.320 154.820 ;
        RECT 42.100 153.440 42.240 155.160 ;
        RECT 42.560 153.440 42.700 155.840 ;
        RECT 43.020 155.480 43.160 163.070 ;
        RECT 43.420 162.980 43.680 163.070 ;
        RECT 43.420 162.300 43.680 162.620 ;
        RECT 43.480 161.600 43.620 162.300 ;
        RECT 43.420 161.280 43.680 161.600 ;
        RECT 42.960 155.160 43.220 155.480 ;
        RECT 43.020 153.440 43.160 155.160 ;
        RECT 43.940 154.800 44.080 165.700 ;
        RECT 45.190 161.765 46.730 162.135 ;
        RECT 44.800 160.600 45.060 160.920 ;
        RECT 44.860 155.820 45.000 160.600 ;
        RECT 45.190 156.325 46.730 156.695 ;
        RECT 48.540 155.820 48.680 168.760 ;
        RECT 44.800 155.500 45.060 155.820 ;
        RECT 48.480 155.500 48.740 155.820 ;
        RECT 45.260 155.160 45.520 155.480 ;
        RECT 43.880 154.480 44.140 154.800 ;
        RECT 42.040 153.120 42.300 153.440 ;
        RECT 42.500 153.120 42.760 153.440 ;
        RECT 42.960 153.120 43.220 153.440 ;
        RECT 43.940 152.080 44.080 154.480 ;
        RECT 45.320 153.440 45.460 155.160 ;
        RECT 45.260 153.120 45.520 153.440 ;
        RECT 41.120 151.760 41.380 152.080 ;
        RECT 43.880 151.760 44.140 152.080 ;
        RECT 44.800 151.420 45.060 151.740 ;
        RECT 40.660 150.400 40.920 150.720 ;
        RECT 44.860 150.120 45.000 151.420 ;
        RECT 45.190 150.885 46.730 151.255 ;
        RECT 44.860 150.040 45.920 150.120 ;
        RECT 38.820 149.720 39.080 150.040 ;
        RECT 40.200 149.720 40.460 150.040 ;
        RECT 44.860 149.980 45.980 150.040 ;
        RECT 45.720 149.720 45.980 149.980 ;
        RECT 37.440 148.700 37.700 149.020 ;
        RECT 37.500 144.260 37.640 148.700 ;
        RECT 37.900 146.660 38.160 146.980 ;
        RECT 37.440 143.940 37.700 144.260 ;
        RECT 36.980 141.220 37.240 141.540 ;
        RECT 33.760 140.880 34.020 141.200 ;
        RECT 36.520 140.880 36.780 141.200 ;
        RECT 33.820 139.500 33.960 140.880 ;
        RECT 33.760 139.180 34.020 139.500 ;
        RECT 31.000 138.840 31.260 139.160 ;
        RECT 31.920 138.840 32.180 139.160 ;
        RECT 32.840 138.840 33.100 139.160 ;
        RECT 31.460 138.500 31.720 138.820 ;
        RECT 31.520 134.400 31.660 138.500 ;
        RECT 31.980 137.120 32.120 138.840 ;
        RECT 36.580 137.120 36.720 140.880 ;
        RECT 37.960 139.840 38.100 146.660 ;
        RECT 40.260 146.640 40.400 149.720 ;
        RECT 45.780 148.000 45.920 149.720 ;
        RECT 45.720 147.680 45.980 148.000 ;
        RECT 39.740 146.320 40.000 146.640 ;
        RECT 40.200 146.320 40.460 146.640 ;
        RECT 38.820 145.980 39.080 146.300 ;
        RECT 38.360 144.280 38.620 144.600 ;
        RECT 38.420 142.560 38.560 144.280 ;
        RECT 38.360 142.240 38.620 142.560 ;
        RECT 37.900 139.520 38.160 139.840 ;
        RECT 31.920 136.800 32.180 137.120 ;
        RECT 36.520 136.800 36.780 137.120 ;
        RECT 27.380 134.220 30.280 134.360 ;
        RECT 27.380 131.680 27.520 134.220 ;
        RECT 30.140 134.060 30.280 134.220 ;
        RECT 31.460 134.080 31.720 134.400 ;
        RECT 30.080 133.740 30.340 134.060 ;
        RECT 35.600 133.630 35.860 133.720 ;
        RECT 36.980 133.630 37.240 133.720 ;
        RECT 35.600 133.490 37.240 133.630 ;
        RECT 35.600 133.400 35.860 133.490 ;
        RECT 36.980 133.400 37.240 133.490 ;
        RECT 37.440 132.380 37.700 132.700 ;
        RECT 27.770 131.845 29.310 132.215 ;
        RECT 37.500 131.680 37.640 132.380 ;
        RECT 27.320 131.360 27.580 131.680 ;
        RECT 37.440 131.360 37.700 131.680 ;
        RECT 37.960 130.660 38.100 139.520 ;
        RECT 38.880 136.100 39.020 145.980 ;
        RECT 39.800 145.280 39.940 146.320 ;
        RECT 47.100 145.980 47.360 146.300 ;
        RECT 45.190 145.445 46.730 145.815 ;
        RECT 39.740 144.960 40.000 145.280 ;
        RECT 47.160 144.600 47.300 145.980 ;
        RECT 47.100 144.280 47.360 144.600 ;
        RECT 47.160 142.560 47.300 144.280 ;
        RECT 48.940 143.940 49.200 144.260 ;
        RECT 47.100 142.240 47.360 142.560 ;
        RECT 44.340 140.880 44.600 141.200 ;
        RECT 44.400 136.440 44.540 140.880 ;
        RECT 44.800 140.540 45.060 140.860 ;
        RECT 47.100 140.540 47.360 140.860 ;
        RECT 44.340 136.120 44.600 136.440 ;
        RECT 44.860 136.100 45.000 140.540 ;
        RECT 45.190 140.005 46.730 140.375 ;
        RECT 47.160 139.840 47.300 140.540 ;
        RECT 47.100 139.520 47.360 139.840 ;
        RECT 47.100 136.800 47.360 137.120 ;
        RECT 38.820 135.780 39.080 136.100 ;
        RECT 44.800 135.780 45.060 136.100 ;
        RECT 43.880 135.100 44.140 135.420 ;
        RECT 43.940 134.060 44.080 135.100 ;
        RECT 45.190 134.565 46.730 134.935 ;
        RECT 47.160 134.360 47.300 136.800 ;
        RECT 46.700 134.220 47.300 134.360 ;
        RECT 46.700 134.060 46.840 134.220 ;
        RECT 43.880 133.740 44.140 134.060 ;
        RECT 46.640 133.740 46.900 134.060 ;
        RECT 39.280 133.400 39.540 133.720 ;
        RECT 37.900 130.340 38.160 130.660 ;
        RECT 39.340 128.960 39.480 133.400 ;
        RECT 44.340 133.060 44.600 133.380 ;
        RECT 42.500 132.380 42.760 132.700 ;
        RECT 42.560 131.680 42.700 132.380 ;
        RECT 42.500 131.360 42.760 131.680 ;
        RECT 41.580 130.340 41.840 130.660 ;
        RECT 39.280 128.640 39.540 128.960 ;
        RECT 27.770 126.405 29.310 126.775 ;
        RECT 41.640 125.220 41.780 130.340 ;
        RECT 44.400 130.320 44.540 133.060 ;
        RECT 46.700 133.040 46.840 133.740 ;
        RECT 46.640 132.720 46.900 133.040 ;
        RECT 48.480 132.380 48.740 132.700 ;
        RECT 48.540 131.680 48.680 132.380 ;
        RECT 48.480 131.360 48.740 131.680 ;
        RECT 49.000 130.660 49.140 143.940 ;
        RECT 49.460 139.500 49.600 169.440 ;
        RECT 50.320 167.740 50.580 168.060 ;
        RECT 51.700 167.740 51.960 168.060 ;
        RECT 50.380 163.640 50.520 167.740 ;
        RECT 51.760 166.360 51.900 167.740 ;
        RECT 52.220 167.040 52.360 182.520 ;
        RECT 53.140 182.520 54.660 182.660 ;
        RECT 52.160 166.720 52.420 167.040 ;
        RECT 53.140 166.440 53.280 182.520 ;
        RECT 53.540 181.340 53.800 181.660 ;
        RECT 54.920 181.340 55.180 181.660 ;
        RECT 53.600 179.620 53.740 181.340 ;
        RECT 54.980 180.640 55.120 181.340 ;
        RECT 54.920 180.320 55.180 180.640 ;
        RECT 54.980 179.960 55.120 180.320 ;
        RECT 54.920 179.640 55.180 179.960 ;
        RECT 53.540 179.300 53.800 179.620 ;
        RECT 53.600 172.480 53.740 179.300 ;
        RECT 55.900 177.920 56.040 187.800 ;
        RECT 57.740 186.080 57.880 196.640 ;
        RECT 57.680 185.760 57.940 186.080 ;
        RECT 56.760 184.740 57.020 185.060 ;
        RECT 56.820 183.020 56.960 184.740 ;
        RECT 56.760 182.700 57.020 183.020 ;
        RECT 56.300 182.360 56.560 182.680 ;
        RECT 56.360 180.640 56.500 182.360 ;
        RECT 56.300 180.320 56.560 180.640 ;
        RECT 56.300 178.620 56.560 178.940 ;
        RECT 55.840 177.600 56.100 177.920 ;
        RECT 56.360 174.520 56.500 178.620 ;
        RECT 56.820 177.580 56.960 182.700 ;
        RECT 58.200 182.000 58.340 209.560 ;
        RECT 64.180 209.200 64.320 211.940 ;
        RECT 64.580 209.560 64.840 209.880 ;
        RECT 74.700 209.560 74.960 209.880 ;
        RECT 64.120 208.880 64.380 209.200 ;
        RECT 61.820 208.540 62.080 208.860 ;
        RECT 61.880 207.840 62.020 208.540 ;
        RECT 62.615 208.005 64.155 208.375 ;
        RECT 61.820 207.520 62.080 207.840 ;
        RECT 64.120 206.840 64.380 207.160 ;
        RECT 64.180 205.120 64.320 206.840 ;
        RECT 64.120 204.800 64.380 205.120 ;
        RECT 58.600 204.120 58.860 204.440 ;
        RECT 58.660 187.100 58.800 204.120 ;
        RECT 62.615 202.565 64.155 202.935 ;
        RECT 62.615 197.125 64.155 197.495 ;
        RECT 63.660 195.620 63.920 195.940 ;
        RECT 61.360 195.280 61.620 195.600 ;
        RECT 62.280 195.280 62.540 195.600 ;
        RECT 60.440 194.940 60.700 195.260 ;
        RECT 60.500 194.240 60.640 194.940 ;
        RECT 61.420 194.240 61.560 195.280 ;
        RECT 62.340 194.240 62.480 195.280 ;
        RECT 63.200 194.940 63.460 195.260 ;
        RECT 60.440 193.920 60.700 194.240 ;
        RECT 61.360 193.920 61.620 194.240 ;
        RECT 62.280 193.920 62.540 194.240 ;
        RECT 63.260 193.220 63.400 194.940 ;
        RECT 63.720 193.220 63.860 195.620 ;
        RECT 64.120 193.920 64.380 194.240 ;
        RECT 64.180 193.220 64.320 193.920 ;
        RECT 63.200 192.900 63.460 193.220 ;
        RECT 63.660 192.900 63.920 193.220 ;
        RECT 64.120 192.900 64.380 193.220 ;
        RECT 61.820 192.220 62.080 192.540 ;
        RECT 61.880 188.800 62.020 192.220 ;
        RECT 62.615 191.685 64.155 192.055 ;
        RECT 61.820 188.480 62.080 188.800 ;
        RECT 58.600 186.780 58.860 187.100 ;
        RECT 61.820 186.780 62.080 187.100 ;
        RECT 60.440 185.760 60.700 186.080 ;
        RECT 58.140 181.680 58.400 182.000 ;
        RECT 57.680 181.340 57.940 181.660 ;
        RECT 57.740 179.960 57.880 181.340 ;
        RECT 57.680 179.640 57.940 179.960 ;
        RECT 58.600 179.300 58.860 179.620 ;
        RECT 57.220 177.600 57.480 177.920 ;
        RECT 56.760 177.260 57.020 177.580 ;
        RECT 56.300 174.200 56.560 174.520 ;
        RECT 54.920 173.860 55.180 174.180 ;
        RECT 54.980 172.480 55.120 173.860 ;
        RECT 53.540 172.160 53.800 172.480 ;
        RECT 54.920 172.160 55.180 172.480 ;
        RECT 56.360 169.420 56.500 174.200 ;
        RECT 57.280 171.800 57.420 177.600 ;
        RECT 58.660 176.900 58.800 179.300 ;
        RECT 59.520 178.960 59.780 179.280 ;
        RECT 59.580 177.240 59.720 178.960 ;
        RECT 59.980 178.620 60.240 178.940 ;
        RECT 60.040 177.920 60.180 178.620 ;
        RECT 59.980 177.600 60.240 177.920 ;
        RECT 59.520 176.920 59.780 177.240 ;
        RECT 57.680 176.755 57.940 176.900 ;
        RECT 57.670 176.385 57.950 176.755 ;
        RECT 58.140 176.580 58.400 176.900 ;
        RECT 58.600 176.580 58.860 176.900 ;
        RECT 58.200 175.200 58.340 176.580 ;
        RECT 58.140 175.110 58.400 175.200 ;
        RECT 58.140 174.970 58.800 175.110 ;
        RECT 58.140 174.880 58.400 174.970 ;
        RECT 57.220 171.480 57.480 171.800 ;
        RECT 58.140 171.480 58.400 171.800 ;
        RECT 58.200 169.420 58.340 171.480 ;
        RECT 58.660 169.420 58.800 174.970 ;
        RECT 59.580 170.780 59.720 176.920 ;
        RECT 59.520 170.460 59.780 170.780 ;
        RECT 59.980 170.460 60.240 170.780 ;
        RECT 56.300 169.100 56.560 169.420 ;
        RECT 58.140 169.100 58.400 169.420 ;
        RECT 58.600 169.100 58.860 169.420 ;
        RECT 57.220 168.420 57.480 168.740 ;
        RECT 58.140 168.420 58.400 168.740 ;
        RECT 53.540 167.740 53.800 168.060 ;
        RECT 53.600 166.700 53.740 167.740 ;
        RECT 51.700 166.040 51.960 166.360 ;
        RECT 52.680 166.300 53.280 166.440 ;
        RECT 53.540 166.380 53.800 166.700 ;
        RECT 51.760 164.320 51.900 166.040 ;
        RECT 52.680 165.680 52.820 166.300 ;
        RECT 52.620 165.360 52.880 165.680 ;
        RECT 53.080 165.360 53.340 165.680 ;
        RECT 52.160 165.020 52.420 165.340 ;
        RECT 51.700 164.000 51.960 164.320 ;
        RECT 50.320 163.320 50.580 163.640 ;
        RECT 50.780 162.300 51.040 162.620 ;
        RECT 50.840 160.920 50.980 162.300 ;
        RECT 49.860 160.600 50.120 160.920 ;
        RECT 50.780 160.600 51.040 160.920 ;
        RECT 49.920 156.160 50.060 160.600 ;
        RECT 51.760 158.960 51.900 164.000 ;
        RECT 52.220 159.900 52.360 165.020 ;
        RECT 52.620 162.980 52.880 163.300 ;
        RECT 52.680 160.240 52.820 162.980 ;
        RECT 53.140 162.620 53.280 165.360 ;
        RECT 53.600 164.320 53.740 166.380 ;
        RECT 56.300 166.040 56.560 166.360 ;
        RECT 53.540 164.000 53.800 164.320 ;
        RECT 56.360 163.300 56.500 166.040 ;
        RECT 56.300 162.980 56.560 163.300 ;
        RECT 56.760 162.980 57.020 163.300 ;
        RECT 53.080 162.300 53.340 162.620 ;
        RECT 52.620 159.920 52.880 160.240 ;
        RECT 52.160 159.580 52.420 159.900 ;
        RECT 51.760 158.820 52.360 158.960 ;
        RECT 53.140 158.880 53.280 162.300 ;
        RECT 56.360 160.240 56.500 162.980 ;
        RECT 56.820 161.600 56.960 162.980 ;
        RECT 56.760 161.280 57.020 161.600 ;
        RECT 56.300 159.920 56.560 160.240 ;
        RECT 51.240 156.860 51.500 157.180 ;
        RECT 51.700 156.860 51.960 157.180 ;
        RECT 49.860 155.840 50.120 156.160 ;
        RECT 51.300 152.420 51.440 156.860 ;
        RECT 51.760 154.800 51.900 156.860 ;
        RECT 51.700 154.480 51.960 154.800 ;
        RECT 51.760 153.100 51.900 154.480 ;
        RECT 51.700 152.780 51.960 153.100 ;
        RECT 51.240 152.100 51.500 152.420 ;
        RECT 51.760 149.700 51.900 152.780 ;
        RECT 52.220 152.080 52.360 158.820 ;
        RECT 53.080 158.560 53.340 158.880 ;
        RECT 57.280 157.600 57.420 168.420 ;
        RECT 57.680 162.300 57.940 162.620 ;
        RECT 57.740 158.880 57.880 162.300 ;
        RECT 57.680 158.560 57.940 158.880 ;
        RECT 56.820 157.460 57.420 157.600 ;
        RECT 53.080 156.860 53.340 157.180 ;
        RECT 53.140 155.480 53.280 156.860 ;
        RECT 56.820 155.820 56.960 157.460 ;
        RECT 57.220 156.860 57.480 157.180 ;
        RECT 57.280 156.160 57.420 156.860 ;
        RECT 57.220 155.840 57.480 156.160 ;
        RECT 56.760 155.500 57.020 155.820 ;
        RECT 53.080 155.160 53.340 155.480 ;
        RECT 56.300 155.160 56.560 155.480 ;
        RECT 53.140 152.420 53.280 155.160 ;
        RECT 56.360 153.440 56.500 155.160 ;
        RECT 56.300 153.120 56.560 153.440 ;
        RECT 53.080 152.100 53.340 152.420 ;
        RECT 52.160 151.760 52.420 152.080 ;
        RECT 51.240 149.380 51.500 149.700 ;
        RECT 51.700 149.380 51.960 149.700 ;
        RECT 51.300 148.000 51.440 149.380 ;
        RECT 51.240 147.680 51.500 148.000 ;
        RECT 51.760 144.600 51.900 149.380 ;
        RECT 52.220 146.300 52.360 151.760 ;
        RECT 53.140 147.320 53.280 152.100 ;
        RECT 56.820 149.360 56.960 155.500 ;
        RECT 57.680 151.420 57.940 151.740 ;
        RECT 56.760 149.040 57.020 149.360 ;
        RECT 53.080 147.000 53.340 147.320 ;
        RECT 56.820 147.230 56.960 149.040 ;
        RECT 57.220 147.230 57.480 147.320 ;
        RECT 56.820 147.090 57.480 147.230 ;
        RECT 57.220 147.000 57.480 147.090 ;
        RECT 56.300 146.720 56.560 146.980 ;
        RECT 56.300 146.660 57.420 146.720 ;
        RECT 56.360 146.580 57.420 146.660 ;
        RECT 52.160 145.980 52.420 146.300 ;
        RECT 53.080 145.980 53.340 146.300 ;
        RECT 56.760 145.980 57.020 146.300 ;
        RECT 51.700 144.280 51.960 144.600 ;
        RECT 49.400 139.180 49.660 139.500 ;
        RECT 52.220 136.440 52.360 145.980 ;
        RECT 53.140 144.260 53.280 145.980 ;
        RECT 53.080 143.940 53.340 144.260 ;
        RECT 53.140 142.560 53.280 143.940 ;
        RECT 56.820 143.920 56.960 145.980 ;
        RECT 56.760 143.600 57.020 143.920 ;
        RECT 53.080 142.240 53.340 142.560 ;
        RECT 52.160 136.120 52.420 136.440 ;
        RECT 51.700 135.780 51.960 136.100 ;
        RECT 51.760 134.060 51.900 135.780 ;
        RECT 51.700 133.740 51.960 134.060 ;
        RECT 48.940 130.340 49.200 130.660 ;
        RECT 44.340 130.000 44.600 130.320 ;
        RECT 42.040 129.660 42.300 129.980 ;
        RECT 43.420 129.660 43.680 129.980 ;
        RECT 42.100 128.280 42.240 129.660 ;
        RECT 42.040 127.960 42.300 128.280 ;
        RECT 43.480 126.240 43.620 129.660 ;
        RECT 45.190 129.125 46.730 129.495 ;
        RECT 52.220 128.280 52.360 136.120 ;
        RECT 53.140 136.100 53.280 142.240 ;
        RECT 53.540 138.500 53.800 138.820 ;
        RECT 55.380 138.500 55.640 138.820 ;
        RECT 53.600 137.120 53.740 138.500 ;
        RECT 53.540 136.800 53.800 137.120 ;
        RECT 53.080 135.780 53.340 136.100 ;
        RECT 53.140 132.700 53.280 135.780 ;
        RECT 53.080 132.380 53.340 132.700 ;
        RECT 54.920 131.360 55.180 131.680 ;
        RECT 54.460 129.660 54.720 129.980 ;
        RECT 54.520 128.960 54.660 129.660 ;
        RECT 53.080 128.640 53.340 128.960 ;
        RECT 54.460 128.640 54.720 128.960 ;
        RECT 53.140 128.360 53.280 128.640 ;
        RECT 54.000 128.360 54.260 128.620 ;
        RECT 53.140 128.300 54.260 128.360 ;
        RECT 52.160 127.960 52.420 128.280 ;
        RECT 53.140 128.220 54.200 128.300 ;
        RECT 54.980 127.940 55.120 131.360 ;
        RECT 55.440 131.000 55.580 138.500 ;
        RECT 56.760 137.820 57.020 138.140 ;
        RECT 56.300 132.380 56.560 132.700 ;
        RECT 56.360 131.340 56.500 132.380 ;
        RECT 56.820 131.680 56.960 137.820 ;
        RECT 57.280 137.120 57.420 146.580 ;
        RECT 57.740 145.280 57.880 151.420 ;
        RECT 58.200 146.980 58.340 168.420 ;
        RECT 58.600 160.600 58.860 160.920 ;
        RECT 58.660 158.880 58.800 160.600 ;
        RECT 58.600 158.560 58.860 158.880 ;
        RECT 60.040 156.160 60.180 170.460 ;
        RECT 60.500 157.520 60.640 185.760 ;
        RECT 61.880 185.060 62.020 186.780 ;
        RECT 62.615 186.245 64.155 186.615 ;
        RECT 61.820 184.740 62.080 185.060 ;
        RECT 61.360 182.760 61.620 183.020 ;
        RECT 61.360 182.700 63.860 182.760 ;
        RECT 61.420 182.680 63.860 182.700 ;
        RECT 60.900 182.360 61.160 182.680 ;
        RECT 61.420 182.620 63.920 182.680 ;
        RECT 64.640 182.660 64.780 209.560 ;
        RECT 74.760 207.840 74.900 209.560 ;
        RECT 75.680 208.860 75.820 215.190 ;
        RECT 80.035 210.725 81.575 211.095 ;
        RECT 85.800 210.220 85.940 215.190 ;
        RECT 95.920 212.260 96.060 215.190 ;
        RECT 97.460 213.445 99.000 213.815 ;
        RECT 106.040 213.280 106.180 215.190 ;
        RECT 105.980 212.960 106.240 213.280 ;
        RECT 116.160 212.260 116.300 215.190 ;
        RECT 126.280 212.260 126.420 215.190 ;
        RECT 132.305 213.445 133.845 213.815 ;
        RECT 136.400 212.260 136.540 215.190 ;
        RECT 86.660 211.940 86.920 212.260 ;
        RECT 95.860 211.940 96.120 212.260 ;
        RECT 104.600 211.940 104.860 212.260 ;
        RECT 116.100 211.940 116.360 212.260 ;
        RECT 126.220 211.940 126.480 212.260 ;
        RECT 136.340 211.940 136.600 212.260 ;
        RECT 86.720 210.560 86.860 211.940 ;
        RECT 89.420 211.260 89.680 211.580 ;
        RECT 99.080 211.260 99.340 211.580 ;
        RECT 86.660 210.240 86.920 210.560 ;
        RECT 83.440 209.900 83.700 210.220 ;
        RECT 85.740 209.900 86.000 210.220 ;
        RECT 79.300 208.880 79.560 209.200 ;
        RECT 75.620 208.540 75.880 208.860 ;
        RECT 74.700 207.520 74.960 207.840 ;
        RECT 70.560 206.500 70.820 206.820 ;
        RECT 72.400 206.500 72.660 206.820 ;
        RECT 65.500 205.820 65.760 206.140 ;
        RECT 68.260 205.820 68.520 206.140 ;
        RECT 65.040 201.740 65.300 202.060 ;
        RECT 65.100 188.800 65.240 201.740 ;
        RECT 65.040 188.480 65.300 188.800 ;
        RECT 65.040 187.460 65.300 187.780 ;
        RECT 63.660 182.360 63.920 182.620 ;
        RECT 64.180 182.520 64.780 182.660 ;
        RECT 65.100 182.660 65.240 187.460 ;
        RECT 65.560 186.080 65.700 205.820 ;
        RECT 68.320 205.120 68.460 205.820 ;
        RECT 68.260 204.800 68.520 205.120 ;
        RECT 69.640 204.120 69.900 204.440 ;
        RECT 70.100 204.120 70.360 204.440 ;
        RECT 66.420 203.440 66.680 203.760 ;
        RECT 67.340 203.440 67.600 203.760 ;
        RECT 66.480 199.340 66.620 203.440 ;
        RECT 66.420 199.020 66.680 199.340 ;
        RECT 66.480 193.560 66.620 199.020 ;
        RECT 66.880 196.300 67.140 196.620 ;
        RECT 66.940 195.260 67.080 196.300 ;
        RECT 66.880 194.940 67.140 195.260 ;
        RECT 66.420 193.240 66.680 193.560 ;
        RECT 65.960 191.200 66.220 191.520 ;
        RECT 65.500 185.760 65.760 186.080 ;
        RECT 66.020 182.660 66.160 191.200 ;
        RECT 66.480 189.820 66.620 193.240 ;
        RECT 66.940 192.880 67.080 194.940 ;
        RECT 67.400 193.560 67.540 203.440 ;
        RECT 69.700 201.380 69.840 204.120 ;
        RECT 69.640 201.060 69.900 201.380 ;
        RECT 67.800 200.380 68.060 200.700 ;
        RECT 67.860 196.960 68.000 200.380 ;
        RECT 69.700 199.680 69.840 201.060 ;
        RECT 69.640 199.360 69.900 199.680 ;
        RECT 67.800 196.640 68.060 196.960 ;
        RECT 70.160 196.280 70.300 204.120 ;
        RECT 70.100 195.960 70.360 196.280 ;
        RECT 67.340 193.240 67.600 193.560 ;
        RECT 68.720 192.900 68.980 193.220 ;
        RECT 66.880 192.560 67.140 192.880 ;
        RECT 67.340 192.220 67.600 192.540 ;
        RECT 66.420 189.500 66.680 189.820 ;
        RECT 67.400 188.120 67.540 192.220 ;
        RECT 67.800 188.480 68.060 188.800 ;
        RECT 67.340 187.800 67.600 188.120 ;
        RECT 66.880 187.460 67.140 187.780 ;
        RECT 66.420 186.780 66.680 187.100 ;
        RECT 66.480 185.740 66.620 186.780 ;
        RECT 66.420 185.420 66.680 185.740 ;
        RECT 66.940 184.720 67.080 187.460 ;
        RECT 67.400 186.080 67.540 187.800 ;
        RECT 67.860 186.080 68.000 188.480 ;
        RECT 67.340 185.760 67.600 186.080 ;
        RECT 67.800 185.760 68.060 186.080 ;
        RECT 66.880 184.400 67.140 184.720 ;
        RECT 65.100 182.520 65.700 182.660 ;
        RECT 66.020 182.520 66.620 182.660 ;
        RECT 60.960 179.620 61.100 182.360 ;
        RECT 64.180 182.000 64.320 182.520 ;
        RECT 64.120 181.680 64.380 182.000 ;
        RECT 65.560 181.660 65.700 182.520 ;
        RECT 65.500 181.340 65.760 181.660 ;
        RECT 62.615 180.805 64.155 181.175 ;
        RECT 60.900 179.300 61.160 179.620 ;
        RECT 64.580 176.240 64.840 176.560 ;
        RECT 62.615 175.365 64.155 175.735 ;
        RECT 63.660 174.880 63.920 175.200 ;
        RECT 63.720 174.715 63.860 174.880 ;
        RECT 63.650 174.345 63.930 174.715 ;
        RECT 64.640 174.180 64.780 176.240 ;
        RECT 64.580 173.860 64.840 174.180 ;
        RECT 65.560 173.840 65.700 181.340 ;
        RECT 66.480 180.040 66.620 182.520 ;
        RECT 66.020 179.900 66.620 180.040 ;
        RECT 66.020 177.580 66.160 179.900 ;
        RECT 66.410 179.105 66.690 179.475 ;
        RECT 65.960 177.260 66.220 177.580 ;
        RECT 65.500 173.520 65.760 173.840 ;
        RECT 65.040 173.180 65.300 173.500 ;
        RECT 65.100 172.480 65.240 173.180 ;
        RECT 65.040 172.160 65.300 172.480 ;
        RECT 64.580 170.460 64.840 170.780 ;
        RECT 62.615 169.925 64.155 170.295 ;
        RECT 64.640 169.080 64.780 170.460 ;
        RECT 64.580 168.760 64.840 169.080 ;
        RECT 63.200 167.740 63.460 168.060 ;
        RECT 63.260 166.360 63.400 167.740 ;
        RECT 63.200 166.040 63.460 166.360 ;
        RECT 62.615 164.485 64.155 164.855 ;
        RECT 66.020 164.320 66.160 177.260 ;
        RECT 65.960 164.000 66.220 164.320 ;
        RECT 64.580 160.260 64.840 160.580 ;
        RECT 62.615 159.045 64.155 159.415 ;
        RECT 60.440 157.200 60.700 157.520 ;
        RECT 59.980 155.840 60.240 156.160 ;
        RECT 64.640 155.480 64.780 160.260 ;
        RECT 65.960 159.580 66.220 159.900 ;
        RECT 66.020 156.160 66.160 159.580 ;
        RECT 65.960 155.840 66.220 156.160 ;
        RECT 64.580 155.160 64.840 155.480 ;
        RECT 61.820 154.140 62.080 154.460 ;
        RECT 61.880 152.420 62.020 154.140 ;
        RECT 62.615 153.605 64.155 153.975 ;
        RECT 64.640 152.420 64.780 155.160 ;
        RECT 66.480 152.420 66.620 179.105 ;
        RECT 66.940 176.900 67.080 184.400 ;
        RECT 68.260 181.680 68.520 182.000 ;
        RECT 67.800 179.980 68.060 180.300 ;
        RECT 67.860 179.475 68.000 179.980 ;
        RECT 67.790 179.105 68.070 179.475 ;
        RECT 67.340 178.620 67.600 178.940 ;
        RECT 66.880 176.580 67.140 176.900 ;
        RECT 67.400 167.040 67.540 178.620 ;
        RECT 68.320 177.580 68.460 181.680 ;
        RECT 68.780 179.960 68.920 192.900 ;
        RECT 69.640 189.500 69.900 189.820 ;
        RECT 69.700 188.120 69.840 189.500 ;
        RECT 69.180 187.800 69.440 188.120 ;
        RECT 69.640 187.800 69.900 188.120 ;
        RECT 70.100 187.800 70.360 188.120 ;
        RECT 69.240 186.080 69.380 187.800 ;
        RECT 69.180 185.760 69.440 186.080 ;
        RECT 69.700 183.020 69.840 187.800 ;
        RECT 70.160 186.955 70.300 187.800 ;
        RECT 70.090 186.585 70.370 186.955 ;
        RECT 69.640 182.700 69.900 183.020 ;
        RECT 70.620 182.340 70.760 206.500 ;
        RECT 71.480 205.820 71.740 206.140 ;
        RECT 71.540 204.440 71.680 205.820 ;
        RECT 72.460 205.120 72.600 206.500 ;
        RECT 77.920 205.820 78.180 206.140 ;
        RECT 72.400 204.800 72.660 205.120 ;
        RECT 77.980 204.780 78.120 205.820 ;
        RECT 79.360 205.120 79.500 208.880 ;
        RECT 82.520 208.540 82.780 208.860 ;
        RECT 82.060 206.500 82.320 206.820 ;
        RECT 80.035 205.285 81.575 205.655 ;
        RECT 82.120 205.120 82.260 206.500 ;
        RECT 79.300 204.800 79.560 205.120 ;
        RECT 82.060 204.800 82.320 205.120 ;
        RECT 77.920 204.460 78.180 204.780 ;
        RECT 71.020 204.120 71.280 204.440 ;
        RECT 71.480 204.120 71.740 204.440 ;
        RECT 71.080 202.400 71.220 204.120 ;
        RECT 73.780 203.440 74.040 203.760 ;
        RECT 73.840 202.400 73.980 203.440 ;
        RECT 71.020 202.080 71.280 202.400 ;
        RECT 73.780 202.080 74.040 202.400 ;
        RECT 77.980 202.060 78.120 204.460 ;
        RECT 78.380 203.100 78.640 203.420 ;
        RECT 77.920 201.740 78.180 202.060 ;
        RECT 78.440 201.380 78.580 203.100 ;
        RECT 78.380 201.060 78.640 201.380 ;
        RECT 71.480 200.720 71.740 201.040 ;
        RECT 71.940 200.720 72.200 201.040 ;
        RECT 71.020 198.340 71.280 198.660 ;
        RECT 71.080 196.960 71.220 198.340 ;
        RECT 71.020 196.640 71.280 196.960 ;
        RECT 71.540 195.940 71.680 200.720 ;
        RECT 72.000 197.980 72.140 200.720 ;
        RECT 79.360 199.590 79.500 204.800 ;
        RECT 82.060 203.780 82.320 204.100 ;
        RECT 80.035 199.845 81.575 200.215 ;
        RECT 80.220 199.590 80.480 199.680 ;
        RECT 79.360 199.450 80.480 199.590 ;
        RECT 76.990 198.825 77.270 199.195 ;
        RECT 78.380 199.020 78.640 199.340 ;
        RECT 77.000 198.680 77.260 198.825 ;
        RECT 71.940 197.660 72.200 197.980 ;
        RECT 73.780 197.660 74.040 197.980 ;
        RECT 72.000 195.940 72.140 197.660 ;
        RECT 71.480 195.620 71.740 195.940 ;
        RECT 71.940 195.620 72.200 195.940 ;
        RECT 72.000 191.520 72.140 195.620 ;
        RECT 73.320 193.920 73.580 194.240 ;
        RECT 72.400 192.900 72.660 193.220 ;
        RECT 71.940 191.200 72.200 191.520 ;
        RECT 71.020 189.500 71.280 189.820 ;
        RECT 71.080 188.120 71.220 189.500 ;
        RECT 71.020 187.800 71.280 188.120 ;
        RECT 71.480 187.120 71.740 187.440 ;
        RECT 71.540 186.080 71.680 187.120 ;
        RECT 71.480 185.760 71.740 186.080 ;
        RECT 72.000 185.400 72.140 191.200 ;
        RECT 72.460 190.160 72.600 192.900 ;
        RECT 73.380 190.840 73.520 193.920 ;
        RECT 73.840 193.560 73.980 197.660 ;
        RECT 78.440 195.940 78.580 199.020 ;
        RECT 78.840 197.660 79.100 197.980 ;
        RECT 77.920 195.620 78.180 195.940 ;
        RECT 78.380 195.620 78.640 195.940 ;
        RECT 77.980 194.240 78.120 195.620 ;
        RECT 78.440 194.240 78.580 195.620 ;
        RECT 78.900 195.600 79.040 197.660 ;
        RECT 79.360 196.960 79.500 199.450 ;
        RECT 80.220 199.360 80.480 199.450 ;
        RECT 81.140 198.340 81.400 198.660 ;
        RECT 79.300 196.640 79.560 196.960 ;
        RECT 81.200 195.600 81.340 198.340 ;
        RECT 82.120 196.960 82.260 203.780 ;
        RECT 82.580 201.720 82.720 208.540 ;
        RECT 83.500 207.840 83.640 209.900 ;
        RECT 89.480 209.880 89.620 211.260 ;
        RECT 84.360 209.560 84.620 209.880 ;
        RECT 89.420 209.560 89.680 209.880 ;
        RECT 83.900 208.540 84.160 208.860 ;
        RECT 83.440 207.520 83.700 207.840 ;
        RECT 83.960 206.140 84.100 208.540 ;
        RECT 84.420 207.160 84.560 209.560 ;
        RECT 88.960 209.220 89.220 209.540 ;
        RECT 84.360 206.840 84.620 207.160 ;
        RECT 84.820 206.500 85.080 206.820 ;
        RECT 83.900 205.820 84.160 206.140 ;
        RECT 84.880 205.120 85.020 206.500 ;
        RECT 84.820 204.800 85.080 205.120 ;
        RECT 89.020 204.440 89.160 209.220 ;
        RECT 97.460 208.005 99.000 208.375 ;
        RECT 92.180 207.180 92.440 207.500 ;
        RECT 91.720 206.500 91.980 206.820 ;
        RECT 88.960 204.120 89.220 204.440 ;
        RECT 91.260 204.120 91.520 204.440 ;
        RECT 84.360 203.780 84.620 204.100 ;
        RECT 82.520 201.400 82.780 201.720 ;
        RECT 82.980 201.060 83.240 201.380 ;
        RECT 82.520 199.360 82.780 199.680 ;
        RECT 82.060 196.640 82.320 196.960 ;
        RECT 78.840 195.280 79.100 195.600 ;
        RECT 81.140 195.280 81.400 195.600 ;
        RECT 77.920 193.920 78.180 194.240 ;
        RECT 78.380 193.920 78.640 194.240 ;
        RECT 73.780 193.240 74.040 193.560 ;
        RECT 73.320 190.520 73.580 190.840 ;
        RECT 73.840 190.500 73.980 193.240 ;
        RECT 78.900 193.220 79.040 195.280 ;
        RECT 79.300 194.940 79.560 195.260 ;
        RECT 79.360 194.240 79.500 194.940 ;
        RECT 80.035 194.405 81.575 194.775 ;
        RECT 79.300 193.920 79.560 194.240 ;
        RECT 78.840 192.900 79.100 193.220 ;
        RECT 77.920 192.220 78.180 192.540 ;
        RECT 81.600 192.450 81.860 192.540 ;
        RECT 82.120 192.450 82.260 196.640 ;
        RECT 82.580 196.620 82.720 199.360 ;
        RECT 83.040 198.660 83.180 201.060 ;
        RECT 82.980 198.340 83.240 198.660 ;
        RECT 82.520 196.300 82.780 196.620 ;
        RECT 81.600 192.310 82.260 192.450 ;
        RECT 81.600 192.220 81.860 192.310 ;
        RECT 77.460 190.520 77.720 190.840 ;
        RECT 73.780 190.180 74.040 190.500 ;
        RECT 72.400 189.840 72.660 190.160 ;
        RECT 73.320 189.840 73.580 190.160 ;
        RECT 71.940 185.080 72.200 185.400 ;
        RECT 72.460 185.060 72.600 189.840 ;
        RECT 73.380 188.800 73.520 189.840 ;
        RECT 73.320 188.480 73.580 188.800 ;
        RECT 73.840 188.120 73.980 190.180 ;
        RECT 76.540 189.500 76.800 189.820 ;
        RECT 72.860 187.800 73.120 188.120 ;
        RECT 73.780 187.800 74.040 188.120 ;
        RECT 75.160 187.800 75.420 188.120 ;
        RECT 72.400 184.740 72.660 185.060 ;
        RECT 72.920 184.380 73.060 187.800 ;
        RECT 74.230 187.265 74.510 187.635 ;
        RECT 74.240 187.120 74.500 187.265 ;
        RECT 75.220 184.720 75.360 187.800 ;
        RECT 76.600 187.100 76.740 189.500 ;
        RECT 77.520 188.800 77.660 190.520 ;
        RECT 77.460 188.480 77.720 188.800 ;
        RECT 76.990 187.265 77.270 187.635 ;
        RECT 77.060 187.100 77.200 187.265 ;
        RECT 76.540 186.780 76.800 187.100 ;
        RECT 77.000 186.780 77.260 187.100 ;
        RECT 76.600 185.740 76.740 186.780 ;
        RECT 76.540 185.420 76.800 185.740 ;
        RECT 75.160 184.400 75.420 184.720 ;
        RECT 71.020 184.060 71.280 184.380 ;
        RECT 72.860 184.060 73.120 184.380 ;
        RECT 70.560 182.020 70.820 182.340 ;
        RECT 68.720 179.640 68.980 179.960 ;
        RECT 71.080 177.920 71.220 184.060 ;
        RECT 71.480 182.020 71.740 182.340 ;
        RECT 71.020 177.600 71.280 177.920 ;
        RECT 68.260 177.490 68.520 177.580 ;
        RECT 67.860 177.350 68.520 177.490 ;
        RECT 67.340 166.720 67.600 167.040 ;
        RECT 67.860 152.760 68.000 177.350 ;
        RECT 68.260 177.260 68.520 177.350 ;
        RECT 68.260 176.580 68.520 176.900 ;
        RECT 68.320 174.180 68.460 176.580 ;
        RECT 68.260 173.860 68.520 174.180 ;
        RECT 68.320 172.480 68.460 173.860 ;
        RECT 69.180 173.520 69.440 173.840 ;
        RECT 68.260 172.160 68.520 172.480 ;
        RECT 68.260 168.080 68.520 168.400 ;
        RECT 68.320 167.040 68.460 168.080 ;
        RECT 69.240 167.120 69.380 173.520 ;
        RECT 70.100 173.180 70.360 173.500 ;
        RECT 70.160 168.860 70.300 173.180 ;
        RECT 71.080 170.780 71.220 177.600 ;
        RECT 71.540 174.520 71.680 182.020 ;
        RECT 71.940 179.300 72.200 179.620 ;
        RECT 72.000 174.860 72.140 179.300 ;
        RECT 72.400 176.920 72.660 177.240 ;
        RECT 72.460 175.200 72.600 176.920 ;
        RECT 72.400 174.880 72.660 175.200 ;
        RECT 71.940 174.540 72.200 174.860 ;
        RECT 71.480 174.200 71.740 174.520 ;
        RECT 72.920 173.500 73.060 184.060 ;
        RECT 75.220 183.020 75.360 184.400 ;
        RECT 75.160 182.700 75.420 183.020 ;
        RECT 76.540 182.930 76.800 183.020 ;
        RECT 76.140 182.790 76.800 182.930 ;
        RECT 76.140 177.920 76.280 182.790 ;
        RECT 76.540 182.700 76.800 182.790 ;
        RECT 77.060 182.195 77.200 186.780 ;
        RECT 77.980 182.660 78.120 192.220 ;
        RECT 78.840 191.200 79.100 191.520 ;
        RECT 78.900 188.800 79.040 191.200 ;
        RECT 79.300 189.500 79.560 189.820 ;
        RECT 78.380 188.480 78.640 188.800 ;
        RECT 78.840 188.480 79.100 188.800 ;
        RECT 78.440 187.440 78.580 188.480 ;
        RECT 78.380 187.120 78.640 187.440 ;
        RECT 78.440 185.740 78.580 187.120 ;
        RECT 79.360 186.160 79.500 189.500 ;
        RECT 80.035 188.965 81.575 189.335 ;
        RECT 82.520 187.800 82.780 188.120 ;
        RECT 82.060 187.460 82.320 187.780 ;
        RECT 80.680 186.780 80.940 187.100 ;
        RECT 78.900 186.020 79.500 186.160 ;
        RECT 78.380 185.420 78.640 185.740 ;
        RECT 77.980 182.520 78.580 182.660 ;
        RECT 76.990 181.825 77.270 182.195 ;
        RECT 78.440 180.640 78.580 182.520 ;
        RECT 78.380 180.320 78.640 180.640 ;
        RECT 76.080 177.600 76.340 177.920 ;
        RECT 73.320 173.860 73.580 174.180 ;
        RECT 74.240 173.860 74.500 174.180 ;
        RECT 72.860 173.180 73.120 173.500 ;
        RECT 73.380 172.480 73.520 173.860 ;
        RECT 74.300 173.500 74.440 173.860 ;
        RECT 74.240 173.180 74.500 173.500 ;
        RECT 73.320 172.160 73.580 172.480 ;
        RECT 74.300 172.390 74.440 173.180 ;
        RECT 76.140 172.480 76.280 177.600 ;
        RECT 77.920 177.260 78.180 177.580 ;
        RECT 76.540 173.860 76.800 174.180 ;
        RECT 76.600 172.480 76.740 173.860 ;
        RECT 73.840 172.250 74.440 172.390 ;
        RECT 72.400 171.480 72.660 171.800 ;
        RECT 71.020 170.460 71.280 170.780 ;
        RECT 72.460 169.080 72.600 171.480 ;
        RECT 72.860 171.140 73.120 171.460 ;
        RECT 70.160 168.720 71.680 168.860 ;
        RECT 72.400 168.760 72.660 169.080 ;
        RECT 68.260 166.720 68.520 167.040 ;
        RECT 68.780 166.980 69.380 167.120 ;
        RECT 67.800 152.440 68.060 152.760 ;
        RECT 61.820 152.100 62.080 152.420 ;
        RECT 64.580 152.100 64.840 152.420 ;
        RECT 66.420 152.160 66.680 152.420 ;
        RECT 66.420 152.100 67.540 152.160 ;
        RECT 61.820 149.040 62.080 149.360 ;
        RECT 61.880 147.660 62.020 149.040 ;
        RECT 62.615 148.165 64.155 148.535 ;
        RECT 61.820 147.340 62.080 147.660 ;
        RECT 58.140 146.660 58.400 146.980 ;
        RECT 57.680 144.960 57.940 145.280 ;
        RECT 57.740 141.540 57.880 144.960 ;
        RECT 58.200 144.260 58.340 146.660 ;
        RECT 59.970 146.465 60.250 146.835 ;
        RECT 60.040 146.300 60.180 146.465 ;
        RECT 59.980 146.210 60.240 146.300 ;
        RECT 59.980 146.070 60.640 146.210 ;
        RECT 59.980 145.980 60.240 146.070 ;
        RECT 58.140 143.940 58.400 144.260 ;
        RECT 59.060 143.600 59.320 143.920 ;
        RECT 57.680 141.220 57.940 141.540 ;
        RECT 59.120 139.160 59.260 143.600 ;
        RECT 60.500 139.840 60.640 146.070 ;
        RECT 61.360 145.980 61.620 146.300 ;
        RECT 61.820 145.980 62.080 146.300 ;
        RECT 61.420 145.280 61.560 145.980 ;
        RECT 61.360 144.960 61.620 145.280 ;
        RECT 61.880 144.940 62.020 145.980 ;
        RECT 61.820 144.620 62.080 144.940 ;
        RECT 64.640 143.580 64.780 152.100 ;
        RECT 66.480 152.020 67.540 152.100 ;
        RECT 65.500 151.420 65.760 151.740 ;
        RECT 65.040 147.000 65.300 147.320 ;
        RECT 65.100 145.280 65.240 147.000 ;
        RECT 65.040 144.960 65.300 145.280 ;
        RECT 65.040 144.280 65.300 144.600 ;
        RECT 60.900 143.260 61.160 143.580 ;
        RECT 61.820 143.260 62.080 143.580 ;
        RECT 64.580 143.260 64.840 143.580 ;
        RECT 60.960 142.220 61.100 143.260 ;
        RECT 60.900 141.900 61.160 142.220 ;
        RECT 61.880 141.540 62.020 143.260 ;
        RECT 62.615 142.725 64.155 143.095 ;
        RECT 61.820 141.220 62.080 141.540 ;
        RECT 59.980 139.520 60.240 139.840 ;
        RECT 60.440 139.520 60.700 139.840 ;
        RECT 60.040 139.240 60.180 139.520 ;
        RECT 64.640 139.500 64.780 143.260 ;
        RECT 65.100 142.560 65.240 144.280 ;
        RECT 65.040 142.240 65.300 142.560 ;
        RECT 65.560 141.880 65.700 151.420 ;
        RECT 67.400 147.320 67.540 152.020 ;
        RECT 67.340 147.000 67.600 147.320 ;
        RECT 66.880 146.835 67.140 146.980 ;
        RECT 66.870 146.465 67.150 146.835 ;
        RECT 65.960 145.980 66.220 146.300 ;
        RECT 66.880 145.980 67.140 146.300 ;
        RECT 65.500 141.560 65.760 141.880 ;
        RECT 65.560 139.500 65.700 141.560 ;
        RECT 57.680 138.840 57.940 139.160 ;
        RECT 59.060 138.840 59.320 139.160 ;
        RECT 60.040 139.100 60.640 139.240 ;
        RECT 64.580 139.180 64.840 139.500 ;
        RECT 65.500 139.180 65.760 139.500 ;
        RECT 57.220 136.800 57.480 137.120 ;
        RECT 57.220 135.780 57.480 136.100 ;
        RECT 57.280 134.400 57.420 135.780 ;
        RECT 57.740 135.760 57.880 138.840 ;
        RECT 59.120 136.440 59.260 138.840 ;
        RECT 59.980 138.500 60.240 138.820 ;
        RECT 59.060 136.120 59.320 136.440 ;
        RECT 59.520 135.780 59.780 136.100 ;
        RECT 57.680 135.440 57.940 135.760 ;
        RECT 59.580 135.420 59.720 135.780 ;
        RECT 60.040 135.760 60.180 138.500 ;
        RECT 60.500 138.140 60.640 139.100 ;
        RECT 60.440 137.820 60.700 138.140 ;
        RECT 60.500 136.780 60.640 137.820 ;
        RECT 62.615 137.285 64.155 137.655 ;
        RECT 60.900 136.800 61.160 137.120 ;
        RECT 60.440 136.460 60.700 136.780 ;
        RECT 59.980 135.440 60.240 135.760 ;
        RECT 59.520 135.100 59.780 135.420 ;
        RECT 57.220 134.080 57.480 134.400 ;
        RECT 56.760 131.360 57.020 131.680 ;
        RECT 56.300 131.020 56.560 131.340 ;
        RECT 55.380 130.680 55.640 131.000 ;
        RECT 57.280 130.320 57.420 134.080 ;
        RECT 60.960 133.720 61.100 136.800 ;
        RECT 64.640 136.440 64.780 139.180 ;
        RECT 66.020 138.050 66.160 145.980 ;
        RECT 66.940 144.940 67.080 145.980 ;
        RECT 66.880 144.620 67.140 144.940 ;
        RECT 66.880 138.050 67.140 138.140 ;
        RECT 66.020 137.910 67.140 138.050 ;
        RECT 66.880 137.820 67.140 137.910 ;
        RECT 62.280 136.120 62.540 136.440 ;
        RECT 64.580 136.120 64.840 136.440 ;
        RECT 62.340 135.420 62.480 136.120 ;
        RECT 61.360 135.100 61.620 135.420 ;
        RECT 62.280 135.100 62.540 135.420 ;
        RECT 60.900 133.400 61.160 133.720 ;
        RECT 57.680 132.720 57.940 133.040 ;
        RECT 57.740 131.340 57.880 132.720 ;
        RECT 57.680 131.020 57.940 131.340 ;
        RECT 57.740 130.660 57.880 131.020 ;
        RECT 57.680 130.340 57.940 130.660 ;
        RECT 57.220 130.000 57.480 130.320 ;
        RECT 59.060 129.660 59.320 129.980 ;
        RECT 60.440 129.660 60.700 129.980 ;
        RECT 59.120 128.620 59.260 129.660 ;
        RECT 59.060 128.300 59.320 128.620 ;
        RECT 60.500 128.280 60.640 129.660 ;
        RECT 60.440 127.960 60.700 128.280 ;
        RECT 49.400 127.620 49.660 127.940 ;
        RECT 54.920 127.620 55.180 127.940 ;
        RECT 45.260 126.940 45.520 127.260 ;
        RECT 43.420 125.920 43.680 126.240 ;
        RECT 41.580 124.900 41.840 125.220 ;
        RECT 45.320 124.880 45.460 126.940 ;
        RECT 45.260 124.560 45.520 124.880 ;
        RECT 47.560 124.220 47.820 124.540 ;
        RECT 45.190 123.685 46.730 124.055 ;
        RECT 47.620 122.840 47.760 124.220 ;
        RECT 49.460 123.180 49.600 127.620 ;
        RECT 60.960 127.600 61.100 133.400 ;
        RECT 61.420 131.680 61.560 135.100 ;
        RECT 62.615 131.845 64.155 132.215 ;
        RECT 61.360 131.360 61.620 131.680 ;
        RECT 64.640 127.940 64.780 136.120 ;
        RECT 65.960 132.380 66.220 132.700 ;
        RECT 66.020 131.680 66.160 132.380 ;
        RECT 65.960 131.360 66.220 131.680 ;
        RECT 66.420 129.660 66.680 129.980 ;
        RECT 64.580 127.620 64.840 127.940 ;
        RECT 54.460 127.280 54.720 127.600 ;
        RECT 60.900 127.280 61.160 127.600 ;
        RECT 54.520 123.520 54.660 127.280 ;
        RECT 59.060 126.940 59.320 127.260 ;
        RECT 59.120 124.880 59.260 126.940 ;
        RECT 62.615 126.405 64.155 126.775 ;
        RECT 64.640 125.220 64.780 127.620 ;
        RECT 65.040 127.280 65.300 127.600 ;
        RECT 65.100 126.240 65.240 127.280 ;
        RECT 65.040 125.920 65.300 126.240 ;
        RECT 66.480 125.560 66.620 129.660 ;
        RECT 66.940 128.960 67.080 137.820 ;
        RECT 67.860 137.120 68.000 152.440 ;
        RECT 68.260 148.700 68.520 149.020 ;
        RECT 68.320 146.980 68.460 148.700 ;
        RECT 68.780 148.000 68.920 166.980 ;
        RECT 69.180 166.040 69.440 166.360 ;
        RECT 69.240 164.320 69.380 166.040 ;
        RECT 71.540 165.340 71.680 168.720 ;
        RECT 71.480 165.020 71.740 165.340 ;
        RECT 69.180 164.000 69.440 164.320 ;
        RECT 70.560 162.980 70.820 163.300 ;
        RECT 70.620 160.580 70.760 162.980 ;
        RECT 71.540 162.960 71.680 165.020 ;
        RECT 72.920 162.960 73.060 171.140 ;
        RECT 73.320 170.460 73.580 170.780 ;
        RECT 73.380 167.040 73.520 170.460 ;
        RECT 73.320 166.720 73.580 167.040 ;
        RECT 73.320 166.040 73.580 166.360 ;
        RECT 71.480 162.640 71.740 162.960 ;
        RECT 71.940 162.640 72.200 162.960 ;
        RECT 72.860 162.640 73.120 162.960 ;
        RECT 71.540 160.920 71.680 162.640 ;
        RECT 71.480 160.600 71.740 160.920 ;
        RECT 70.560 160.260 70.820 160.580 ;
        RECT 70.620 158.880 70.760 160.260 ;
        RECT 72.000 159.900 72.140 162.640 ;
        RECT 71.940 159.580 72.200 159.900 ;
        RECT 70.560 158.560 70.820 158.880 ;
        RECT 72.000 157.860 72.140 159.580 ;
        RECT 72.920 158.880 73.060 162.640 ;
        RECT 72.860 158.560 73.120 158.880 ;
        RECT 71.940 157.540 72.200 157.860 ;
        RECT 73.380 157.715 73.520 166.040 ;
        RECT 73.310 157.345 73.590 157.715 ;
        RECT 71.020 156.860 71.280 157.180 ;
        RECT 71.080 156.160 71.220 156.860 ;
        RECT 71.020 155.840 71.280 156.160 ;
        RECT 73.380 155.560 73.520 157.345 ;
        RECT 73.840 156.160 73.980 172.250 ;
        RECT 74.700 172.160 74.960 172.480 ;
        RECT 76.080 172.160 76.340 172.480 ;
        RECT 76.540 172.160 76.800 172.480 ;
        RECT 74.240 171.480 74.500 171.800 ;
        RECT 74.300 169.420 74.440 171.480 ;
        RECT 74.760 170.780 74.900 172.160 ;
        RECT 77.980 171.800 78.120 177.260 ;
        RECT 78.440 174.520 78.580 180.320 ;
        RECT 78.900 179.280 79.040 186.020 ;
        RECT 79.300 184.740 79.560 185.060 ;
        RECT 78.840 178.960 79.100 179.280 ;
        RECT 79.360 177.240 79.500 184.740 ;
        RECT 80.740 184.720 80.880 186.780 ;
        RECT 80.680 184.400 80.940 184.720 ;
        RECT 80.035 183.525 81.575 183.895 ;
        RECT 82.120 182.680 82.260 187.460 ;
        RECT 82.580 185.060 82.720 187.800 ;
        RECT 82.520 184.740 82.780 185.060 ;
        RECT 82.060 182.360 82.320 182.680 ;
        RECT 80.035 178.085 81.575 178.455 ;
        RECT 79.300 176.920 79.560 177.240 ;
        RECT 82.120 176.220 82.260 182.360 ;
        RECT 82.520 178.960 82.780 179.280 ;
        RECT 82.580 177.920 82.720 178.960 ;
        RECT 82.520 177.600 82.780 177.920 ;
        RECT 78.840 176.075 79.100 176.220 ;
        RECT 78.830 175.705 79.110 176.075 ;
        RECT 82.060 175.900 82.320 176.220 ;
        RECT 82.120 174.520 82.260 175.900 ;
        RECT 78.380 174.200 78.640 174.520 ;
        RECT 82.060 174.200 82.320 174.520 ;
        RECT 82.520 173.180 82.780 173.500 ;
        RECT 80.035 172.645 81.575 173.015 ;
        RECT 82.060 172.160 82.320 172.480 ;
        RECT 77.460 171.480 77.720 171.800 ;
        RECT 77.920 171.480 78.180 171.800 ;
        RECT 79.300 171.480 79.560 171.800 ;
        RECT 76.540 171.140 76.800 171.460 ;
        RECT 75.620 170.800 75.880 171.120 ;
        RECT 74.700 170.460 74.960 170.780 ;
        RECT 74.240 169.100 74.500 169.420 ;
        RECT 74.300 166.700 74.440 169.100 ;
        RECT 75.160 167.740 75.420 168.060 ;
        RECT 75.220 166.700 75.360 167.740 ;
        RECT 74.240 166.380 74.500 166.700 ;
        RECT 75.160 166.380 75.420 166.700 ;
        RECT 74.700 165.700 74.960 166.020 ;
        RECT 75.160 165.700 75.420 166.020 ;
        RECT 74.240 164.000 74.500 164.320 ;
        RECT 74.300 160.580 74.440 164.000 ;
        RECT 74.760 161.260 74.900 165.700 ;
        RECT 75.220 164.320 75.360 165.700 ;
        RECT 75.160 164.000 75.420 164.320 ;
        RECT 75.220 161.600 75.360 164.000 ;
        RECT 75.160 161.280 75.420 161.600 ;
        RECT 74.700 160.940 74.960 161.260 ;
        RECT 74.240 160.260 74.500 160.580 ;
        RECT 74.300 157.180 74.440 160.260 ;
        RECT 74.240 156.860 74.500 157.180 ;
        RECT 73.780 155.840 74.040 156.160 ;
        RECT 73.380 155.420 73.980 155.560 ;
        RECT 73.840 154.460 73.980 155.420 ;
        RECT 73.320 154.140 73.580 154.460 ;
        RECT 73.780 154.140 74.040 154.460 ;
        RECT 73.380 152.420 73.520 154.140 ;
        RECT 74.760 152.420 74.900 160.940 ;
        RECT 75.160 160.600 75.420 160.920 ;
        RECT 75.220 160.435 75.360 160.600 ;
        RECT 75.150 160.065 75.430 160.435 ;
        RECT 75.220 158.200 75.360 160.065 ;
        RECT 75.680 158.880 75.820 170.800 ;
        RECT 76.600 170.780 76.740 171.140 ;
        RECT 76.540 170.460 76.800 170.780 ;
        RECT 76.080 168.760 76.340 169.080 ;
        RECT 76.140 165.680 76.280 168.760 ;
        RECT 76.080 165.360 76.340 165.680 ;
        RECT 76.140 160.580 76.280 165.360 ;
        RECT 76.600 160.580 76.740 170.460 ;
        RECT 77.000 169.100 77.260 169.420 ;
        RECT 77.060 163.300 77.200 169.100 ;
        RECT 77.520 165.340 77.660 171.480 ;
        RECT 77.460 165.020 77.720 165.340 ;
        RECT 77.980 164.320 78.120 171.480 ;
        RECT 78.380 167.740 78.640 168.060 ;
        RECT 77.920 164.000 78.180 164.320 ;
        RECT 78.440 163.640 78.580 167.740 ;
        RECT 79.360 167.040 79.500 171.480 ;
        RECT 80.035 167.205 81.575 167.575 ;
        RECT 79.300 166.720 79.560 167.040 ;
        RECT 78.380 163.320 78.640 163.640 ;
        RECT 77.000 162.980 77.260 163.300 ;
        RECT 77.000 161.280 77.260 161.600 ;
        RECT 77.060 160.920 77.200 161.280 ;
        RECT 77.000 160.600 77.260 160.920 ;
        RECT 76.080 160.260 76.340 160.580 ;
        RECT 76.540 160.260 76.800 160.580 ;
        RECT 75.620 158.560 75.880 158.880 ;
        RECT 75.160 157.880 75.420 158.200 ;
        RECT 75.680 155.140 75.820 158.560 ;
        RECT 75.620 154.820 75.880 155.140 ;
        RECT 75.160 154.140 75.420 154.460 ;
        RECT 73.320 152.100 73.580 152.420 ;
        RECT 74.240 152.100 74.500 152.420 ;
        RECT 74.700 152.100 74.960 152.420 ;
        RECT 72.400 151.420 72.660 151.740 ;
        RECT 73.780 151.420 74.040 151.740 ;
        RECT 68.720 147.680 68.980 148.000 ;
        RECT 68.260 146.660 68.520 146.980 ;
        RECT 70.100 146.660 70.360 146.980 ;
        RECT 70.160 145.280 70.300 146.660 ;
        RECT 70.100 144.960 70.360 145.280 ;
        RECT 72.460 144.940 72.600 151.420 ;
        RECT 73.840 150.120 73.980 151.420 ;
        RECT 74.300 150.720 74.440 152.100 ;
        RECT 74.240 150.400 74.500 150.720 ;
        RECT 73.840 149.980 74.440 150.120 ;
        RECT 72.400 144.620 72.660 144.940 ;
        RECT 72.860 137.820 73.120 138.140 ;
        RECT 73.320 137.820 73.580 138.140 ;
        RECT 67.800 136.800 68.060 137.120 ;
        RECT 67.860 136.520 68.000 136.800 ;
        RECT 67.860 136.380 68.920 136.520 ;
        RECT 72.920 136.440 73.060 137.820 ;
        RECT 73.380 137.120 73.520 137.820 ;
        RECT 73.320 136.800 73.580 137.120 ;
        RECT 67.800 135.440 68.060 135.760 ;
        RECT 67.860 134.360 68.000 135.440 ;
        RECT 68.260 134.360 68.520 134.400 ;
        RECT 67.860 134.220 68.520 134.360 ;
        RECT 68.260 134.080 68.520 134.220 ;
        RECT 68.780 133.800 68.920 136.380 ;
        RECT 72.860 136.120 73.120 136.440 ;
        RECT 72.400 135.100 72.660 135.420 ;
        RECT 73.780 135.100 74.040 135.420 ;
        RECT 69.180 134.080 69.440 134.400 ;
        RECT 67.860 133.660 68.920 133.800 ;
        RECT 67.860 133.380 68.000 133.660 ;
        RECT 67.800 133.060 68.060 133.380 ;
        RECT 69.240 132.700 69.380 134.080 ;
        RECT 72.460 133.720 72.600 135.100 ;
        RECT 73.840 134.400 73.980 135.100 ;
        RECT 73.780 134.080 74.040 134.400 ;
        RECT 74.300 134.360 74.440 149.980 ;
        RECT 74.300 134.220 74.900 134.360 ;
        RECT 72.400 133.400 72.660 133.720 ;
        RECT 73.840 133.040 73.980 134.080 ;
        RECT 74.760 133.040 74.900 134.220 ;
        RECT 75.220 134.060 75.360 154.140 ;
        RECT 75.610 153.945 75.890 154.315 ;
        RECT 75.680 150.040 75.820 153.945 ;
        RECT 76.140 152.080 76.280 160.260 ;
        RECT 76.600 157.180 76.740 160.260 ;
        RECT 78.440 159.900 78.580 163.320 ;
        RECT 80.035 161.765 81.575 162.135 ;
        RECT 82.120 161.000 82.260 172.160 ;
        RECT 82.580 166.360 82.720 173.180 ;
        RECT 83.040 172.480 83.180 198.340 ;
        RECT 83.440 188.315 83.700 188.460 ;
        RECT 83.430 187.945 83.710 188.315 ;
        RECT 83.500 179.620 83.640 187.945 ;
        RECT 83.900 187.010 84.160 187.100 ;
        RECT 84.420 187.010 84.560 203.780 ;
        RECT 84.820 200.380 85.080 200.700 ;
        RECT 84.880 199.680 85.020 200.380 ;
        RECT 84.820 199.360 85.080 199.680 ;
        RECT 89.020 196.280 89.160 204.120 ;
        RECT 91.320 202.400 91.460 204.120 ;
        RECT 91.260 202.080 91.520 202.400 ;
        RECT 91.780 201.800 91.920 206.500 ;
        RECT 92.240 203.420 92.380 207.180 ;
        RECT 99.140 206.820 99.280 211.260 ;
        RECT 104.660 210.560 104.800 211.940 ;
        RECT 107.820 211.260 108.080 211.580 ;
        RECT 108.740 211.260 109.000 211.580 ;
        RECT 116.560 211.260 116.820 211.580 ;
        RECT 127.600 211.260 127.860 211.580 ;
        RECT 137.720 211.260 137.980 211.580 ;
        RECT 104.600 210.240 104.860 210.560 ;
        RECT 107.880 210.220 108.020 211.260 ;
        RECT 107.820 209.900 108.080 210.220 ;
        RECT 100.000 209.560 100.260 209.880 ;
        RECT 100.060 207.840 100.200 209.560 ;
        RECT 105.520 208.540 105.780 208.860 ;
        RECT 100.000 207.520 100.260 207.840 ;
        RECT 99.080 206.500 99.340 206.820 ;
        RECT 105.580 206.480 105.720 208.540 ;
        RECT 108.800 206.480 108.940 211.260 ;
        RECT 114.880 210.725 116.420 211.095 ;
        RECT 116.620 210.560 116.760 211.260 ;
        RECT 116.560 210.240 116.820 210.560 ;
        RECT 122.540 209.560 122.800 209.880 ;
        RECT 124.840 209.560 125.100 209.880 ;
        RECT 111.500 208.880 111.760 209.200 ;
        RECT 110.580 206.500 110.840 206.820 ;
        RECT 105.520 206.160 105.780 206.480 ;
        RECT 108.740 206.160 109.000 206.480 ;
        RECT 93.100 205.820 93.360 206.140 ;
        RECT 99.080 205.820 99.340 206.140 ;
        RECT 110.120 205.820 110.380 206.140 ;
        RECT 93.160 205.120 93.300 205.820 ;
        RECT 93.100 204.800 93.360 205.120 ;
        RECT 92.180 203.100 92.440 203.420 ;
        RECT 92.640 203.100 92.900 203.420 ;
        RECT 91.320 201.660 91.920 201.800 ;
        RECT 88.960 195.960 89.220 196.280 ;
        RECT 86.200 193.920 86.460 194.240 ;
        RECT 86.260 191.180 86.400 193.920 ;
        RECT 89.020 193.560 89.160 195.960 ;
        RECT 88.960 193.240 89.220 193.560 ;
        RECT 89.020 191.520 89.160 193.240 ;
        RECT 86.660 191.200 86.920 191.520 ;
        RECT 88.960 191.200 89.220 191.520 ;
        RECT 86.200 190.860 86.460 191.180 ;
        RECT 86.260 188.460 86.400 190.860 ;
        RECT 84.820 188.140 85.080 188.460 ;
        RECT 86.200 188.140 86.460 188.460 ;
        RECT 83.900 186.870 84.560 187.010 ;
        RECT 83.900 186.780 84.160 186.870 ;
        RECT 83.960 182.340 84.100 186.780 ;
        RECT 84.880 185.740 85.020 188.140 ;
        RECT 84.820 185.420 85.080 185.740 ;
        RECT 83.900 182.020 84.160 182.340 ;
        RECT 83.960 181.660 84.100 182.020 ;
        RECT 83.900 181.340 84.160 181.660 ;
        RECT 86.720 180.640 86.860 191.200 ;
        RECT 87.580 186.955 87.840 187.100 ;
        RECT 87.570 186.585 87.850 186.955 ;
        RECT 90.340 185.760 90.600 186.080 ;
        RECT 87.580 185.080 87.840 185.400 ;
        RECT 87.640 180.640 87.780 185.080 ;
        RECT 88.960 182.700 89.220 183.020 ;
        RECT 86.660 180.320 86.920 180.640 ;
        RECT 87.580 180.320 87.840 180.640 ;
        RECT 83.440 179.300 83.700 179.620 ;
        RECT 87.580 178.620 87.840 178.940 ;
        RECT 87.640 177.920 87.780 178.620 ;
        RECT 87.580 177.600 87.840 177.920 ;
        RECT 83.440 176.920 83.700 177.240 ;
        RECT 82.980 172.160 83.240 172.480 ;
        RECT 83.500 168.400 83.640 176.920 ;
        RECT 85.280 174.200 85.540 174.520 ;
        RECT 85.340 172.480 85.480 174.200 ;
        RECT 85.280 172.390 85.540 172.480 ;
        RECT 84.880 172.250 85.540 172.390 ;
        RECT 83.440 168.080 83.700 168.400 ;
        RECT 82.520 166.040 82.780 166.360 ;
        RECT 82.520 162.300 82.780 162.620 ;
        RECT 81.200 160.860 82.260 161.000 ;
        RECT 82.580 160.920 82.720 162.300 ;
        RECT 81.200 160.580 81.340 160.860 ;
        RECT 82.520 160.600 82.780 160.920 ;
        RECT 83.440 160.830 83.700 160.920 ;
        RECT 83.040 160.690 83.700 160.830 ;
        RECT 81.140 160.260 81.400 160.580 ;
        RECT 81.600 160.435 81.860 160.580 ;
        RECT 80.680 159.920 80.940 160.240 ;
        RECT 78.380 159.580 78.640 159.900 ;
        RECT 80.740 158.960 80.880 159.920 ;
        RECT 81.200 159.900 81.340 160.260 ;
        RECT 81.590 160.065 81.870 160.435 ;
        RECT 81.660 159.900 81.800 160.065 ;
        RECT 81.140 159.580 81.400 159.900 ;
        RECT 81.600 159.580 81.860 159.900 ;
        RECT 83.040 158.960 83.180 160.690 ;
        RECT 83.440 160.600 83.700 160.690 ;
        RECT 83.900 160.600 84.160 160.920 ;
        RECT 83.960 158.960 84.100 160.600 ;
        RECT 78.380 158.560 78.640 158.880 ;
        RECT 80.740 158.820 83.180 158.960 ;
        RECT 83.500 158.820 84.100 158.960 ;
        RECT 84.880 158.880 85.020 172.250 ;
        RECT 85.280 172.160 85.540 172.250 ;
        RECT 89.020 172.140 89.160 182.700 ;
        RECT 89.880 179.300 90.140 179.620 ;
        RECT 89.940 175.200 90.080 179.300 ;
        RECT 90.400 175.200 90.540 185.760 ;
        RECT 90.800 184.060 91.060 184.380 ;
        RECT 90.860 182.340 91.000 184.060 ;
        RECT 90.800 182.020 91.060 182.340 ;
        RECT 90.860 177.920 91.000 182.020 ;
        RECT 90.800 177.600 91.060 177.920 ;
        RECT 89.880 174.880 90.140 175.200 ;
        RECT 90.340 174.880 90.600 175.200 ;
        RECT 90.400 172.480 90.540 174.880 ;
        RECT 91.320 174.180 91.460 201.660 ;
        RECT 92.240 199.000 92.380 203.100 ;
        RECT 92.700 199.340 92.840 203.100 ;
        RECT 97.460 202.565 99.000 202.935 ;
        RECT 99.140 202.060 99.280 205.820 ;
        RECT 106.900 203.440 107.160 203.760 ;
        RECT 99.540 203.100 99.800 203.420 ;
        RECT 99.080 201.740 99.340 202.060 ;
        RECT 92.640 199.020 92.900 199.340 ;
        RECT 92.180 198.680 92.440 199.000 ;
        RECT 99.140 197.980 99.280 201.740 ;
        RECT 94.020 197.660 94.280 197.980 ;
        RECT 99.080 197.660 99.340 197.980 ;
        RECT 93.560 192.220 93.820 192.540 ;
        RECT 92.180 190.860 92.440 191.180 ;
        RECT 92.240 188.120 92.380 190.860 ;
        RECT 92.640 189.840 92.900 190.160 ;
        RECT 92.700 188.120 92.840 189.840 ;
        RECT 92.180 187.800 92.440 188.120 ;
        RECT 92.640 187.800 92.900 188.120 ;
        RECT 92.640 186.780 92.900 187.100 ;
        RECT 91.720 181.340 91.980 181.660 ;
        RECT 91.260 173.860 91.520 174.180 ;
        RECT 90.340 172.160 90.600 172.480 ;
        RECT 88.960 171.820 89.220 172.140 ;
        RECT 85.280 168.420 85.540 168.740 ;
        RECT 85.340 162.620 85.480 168.420 ;
        RECT 91.320 168.060 91.460 173.860 ;
        RECT 91.260 167.740 91.520 168.060 ;
        RECT 90.800 162.640 91.060 162.960 ;
        RECT 85.280 162.300 85.540 162.620 ;
        RECT 90.860 160.580 91.000 162.640 ;
        RECT 86.660 160.260 86.920 160.580 ;
        RECT 90.800 160.260 91.060 160.580 ;
        RECT 78.440 157.180 78.580 158.560 ;
        RECT 83.500 157.600 83.640 158.820 ;
        RECT 84.820 158.560 85.080 158.880 ;
        RECT 83.040 157.460 83.640 157.600 ;
        RECT 84.360 157.540 84.620 157.860 ;
        RECT 85.740 157.540 86.000 157.860 ;
        RECT 76.540 156.860 76.800 157.180 ;
        RECT 78.380 156.860 78.640 157.180 ;
        RECT 78.440 152.420 78.580 156.860 ;
        RECT 80.035 156.325 81.575 156.695 ;
        RECT 83.040 155.820 83.180 157.460 ;
        RECT 83.440 156.860 83.700 157.180 ;
        RECT 83.500 155.820 83.640 156.860 ;
        RECT 84.420 155.820 84.560 157.540 ;
        RECT 85.800 156.160 85.940 157.540 ;
        RECT 85.740 155.840 86.000 156.160 ;
        RECT 82.980 155.500 83.240 155.820 ;
        RECT 83.440 155.500 83.700 155.820 ;
        RECT 84.360 155.500 84.620 155.820 ;
        RECT 86.200 155.500 86.460 155.820 ;
        RECT 82.520 152.440 82.780 152.760 ;
        RECT 78.380 152.100 78.640 152.420 ;
        RECT 76.080 151.760 76.340 152.080 ;
        RECT 76.540 151.420 76.800 151.740 ;
        RECT 76.600 150.720 76.740 151.420 ;
        RECT 80.035 150.885 81.575 151.255 ;
        RECT 76.540 150.400 76.800 150.720 ;
        RECT 75.620 149.720 75.880 150.040 ;
        RECT 79.300 149.380 79.560 149.700 ;
        RECT 77.920 147.340 78.180 147.660 ;
        RECT 77.460 146.320 77.720 146.640 ;
        RECT 77.520 145.280 77.660 146.320 ;
        RECT 77.980 146.300 78.120 147.340 ;
        RECT 78.840 146.660 79.100 146.980 ;
        RECT 77.920 145.980 78.180 146.300 ;
        RECT 78.380 145.980 78.640 146.300 ;
        RECT 77.460 144.960 77.720 145.280 ;
        RECT 76.540 141.220 76.800 141.540 ;
        RECT 77.460 141.220 77.720 141.540 ;
        RECT 75.620 140.540 75.880 140.860 ;
        RECT 75.680 136.635 75.820 140.540 ;
        RECT 76.600 139.500 76.740 141.220 ;
        RECT 77.000 140.540 77.260 140.860 ;
        RECT 76.540 139.180 76.800 139.500 ;
        RECT 76.080 137.820 76.340 138.140 ;
        RECT 76.140 137.120 76.280 137.820 ;
        RECT 76.080 136.800 76.340 137.120 ;
        RECT 75.610 136.265 75.890 136.635 ;
        RECT 75.680 135.760 75.820 136.265 ;
        RECT 77.060 135.760 77.200 140.540 ;
        RECT 77.520 139.500 77.660 141.220 ;
        RECT 77.460 139.180 77.720 139.500 ;
        RECT 77.980 138.480 78.120 145.980 ;
        RECT 78.440 145.280 78.580 145.980 ;
        RECT 78.380 144.960 78.640 145.280 ;
        RECT 78.900 144.600 79.040 146.660 ;
        RECT 79.360 146.300 79.500 149.380 ;
        RECT 82.580 146.980 82.720 152.440 ;
        RECT 83.500 151.740 83.640 155.500 ;
        RECT 84.820 154.820 85.080 155.140 ;
        RECT 84.880 153.440 85.020 154.820 ;
        RECT 84.820 153.120 85.080 153.440 ;
        RECT 86.260 152.420 86.400 155.500 ;
        RECT 86.200 152.100 86.460 152.420 ;
        RECT 83.440 151.420 83.700 151.740 ;
        RECT 83.500 146.980 83.640 151.420 ;
        RECT 82.520 146.890 82.780 146.980 ;
        RECT 82.520 146.750 83.180 146.890 ;
        RECT 82.520 146.660 82.780 146.750 ;
        RECT 79.300 145.980 79.560 146.300 ;
        RECT 78.840 144.280 79.100 144.600 ;
        RECT 78.380 143.940 78.640 144.260 ;
        RECT 78.440 138.820 78.580 143.940 ;
        RECT 78.380 138.500 78.640 138.820 ;
        RECT 77.920 138.160 78.180 138.480 ;
        RECT 77.980 135.955 78.120 138.160 ;
        RECT 75.620 135.440 75.880 135.760 ;
        RECT 77.000 135.440 77.260 135.760 ;
        RECT 77.910 135.585 78.190 135.955 ;
        RECT 78.440 135.760 78.580 138.500 ;
        RECT 78.380 135.440 78.640 135.760 ;
        RECT 76.080 135.100 76.340 135.420 ;
        RECT 75.160 133.740 75.420 134.060 ;
        RECT 76.140 133.380 76.280 135.100 ;
        RECT 76.080 133.060 76.340 133.380 ;
        RECT 73.780 132.720 74.040 133.040 ;
        RECT 74.700 132.720 74.960 133.040 ;
        RECT 69.180 132.380 69.440 132.700 ;
        RECT 73.840 130.320 73.980 132.720 ;
        RECT 73.780 130.000 74.040 130.320 ;
        RECT 74.760 129.980 74.900 132.720 ;
        RECT 77.060 132.700 77.200 135.440 ;
        RECT 77.000 132.380 77.260 132.700 ;
        RECT 78.900 131.340 79.040 144.280 ;
        RECT 79.360 139.840 79.500 145.980 ;
        RECT 80.035 145.445 81.575 145.815 ;
        RECT 82.060 144.280 82.320 144.600 ;
        RECT 80.035 140.005 81.575 140.375 ;
        RECT 79.300 139.520 79.560 139.840 ;
        RECT 82.120 139.500 82.260 144.280 ;
        RECT 83.040 143.920 83.180 146.750 ;
        RECT 83.440 146.660 83.700 146.980 ;
        RECT 82.980 143.600 83.240 143.920 ;
        RECT 82.060 139.180 82.320 139.500 ;
        RECT 79.300 138.840 79.560 139.160 ;
        RECT 80.220 138.840 80.480 139.160 ;
        RECT 78.840 131.020 79.100 131.340 ;
        RECT 75.620 130.680 75.880 131.000 ;
        RECT 75.160 130.340 75.420 130.660 ;
        RECT 75.680 130.400 75.820 130.680 ;
        RECT 74.700 129.660 74.960 129.980 ;
        RECT 75.220 128.960 75.360 130.340 ;
        RECT 75.680 130.260 76.280 130.400 ;
        RECT 76.140 129.980 76.280 130.260 ;
        RECT 76.080 129.660 76.340 129.980 ;
        RECT 66.880 128.640 67.140 128.960 ;
        RECT 75.160 128.640 75.420 128.960 ;
        RECT 78.900 128.620 79.040 131.020 ;
        RECT 79.360 130.320 79.500 138.840 ;
        RECT 80.280 138.390 80.420 138.840 ;
        RECT 81.140 138.390 81.400 138.480 ;
        RECT 80.280 138.250 81.400 138.390 ;
        RECT 80.280 136.100 80.420 138.250 ;
        RECT 81.140 138.160 81.400 138.250 ;
        RECT 82.520 137.820 82.780 138.140 ;
        RECT 82.060 136.460 82.320 136.780 ;
        RECT 80.220 135.780 80.480 136.100 ;
        RECT 80.035 134.565 81.575 134.935 ;
        RECT 82.120 130.660 82.260 136.460 ;
        RECT 82.580 135.760 82.720 137.820 ;
        RECT 82.520 135.440 82.780 135.760 ;
        RECT 83.040 135.160 83.180 143.600 ;
        RECT 83.500 143.580 83.640 146.660 ;
        RECT 86.260 145.280 86.400 152.100 ;
        RECT 86.720 146.980 86.860 160.260 ;
        RECT 91.780 158.200 91.920 181.340 ;
        RECT 92.170 179.105 92.450 179.475 ;
        RECT 92.240 178.940 92.380 179.105 ;
        RECT 92.180 178.620 92.440 178.940 ;
        RECT 92.180 176.580 92.440 176.900 ;
        RECT 92.240 174.520 92.380 176.580 ;
        RECT 92.180 174.200 92.440 174.520 ;
        RECT 92.240 172.480 92.380 174.200 ;
        RECT 92.180 172.160 92.440 172.480 ;
        RECT 92.700 166.360 92.840 186.780 ;
        RECT 93.100 174.200 93.360 174.520 ;
        RECT 93.160 169.760 93.300 174.200 ;
        RECT 93.100 169.440 93.360 169.760 ;
        RECT 92.640 166.040 92.900 166.360 ;
        RECT 92.180 163.320 92.440 163.640 ;
        RECT 92.240 160.920 92.380 163.320 ;
        RECT 93.620 163.300 93.760 192.220 ;
        RECT 94.080 190.500 94.220 197.660 ;
        RECT 97.460 197.125 99.000 197.495 ;
        RECT 99.140 195.600 99.280 197.660 ;
        RECT 99.080 195.280 99.340 195.600 ;
        RECT 98.620 193.240 98.880 193.560 ;
        RECT 96.780 192.220 97.040 192.540 ;
        RECT 98.680 192.450 98.820 193.240 ;
        RECT 98.680 192.310 99.280 192.450 ;
        RECT 96.840 191.180 96.980 192.220 ;
        RECT 97.460 191.685 99.000 192.055 ;
        RECT 96.780 190.860 97.040 191.180 ;
        RECT 94.020 190.180 94.280 190.500 ;
        RECT 99.140 190.240 99.280 192.310 ;
        RECT 95.400 189.840 95.660 190.160 ;
        RECT 97.700 189.840 97.960 190.160 ;
        RECT 98.680 190.100 99.280 190.240 ;
        RECT 94.480 187.800 94.740 188.120 ;
        RECT 94.940 187.800 95.200 188.120 ;
        RECT 94.540 183.020 94.680 187.800 ;
        RECT 95.000 187.635 95.140 187.800 ;
        RECT 94.930 187.265 95.210 187.635 ;
        RECT 94.480 182.700 94.740 183.020 ;
        RECT 94.480 180.320 94.740 180.640 ;
        RECT 94.540 179.620 94.680 180.320 ;
        RECT 94.480 179.300 94.740 179.620 ;
        RECT 94.020 176.920 94.280 177.240 ;
        RECT 94.080 174.520 94.220 176.920 ;
        RECT 94.480 175.900 94.740 176.220 ;
        RECT 94.020 174.200 94.280 174.520 ;
        RECT 94.540 173.500 94.680 175.900 ;
        RECT 94.480 173.180 94.740 173.500 ;
        RECT 94.540 172.480 94.680 173.180 ;
        RECT 94.480 172.160 94.740 172.480 ;
        RECT 95.460 169.420 95.600 189.840 ;
        RECT 97.760 188.800 97.900 189.840 ;
        RECT 97.700 188.480 97.960 188.800 ;
        RECT 98.680 187.780 98.820 190.100 ;
        RECT 99.080 189.500 99.340 189.820 ;
        RECT 98.620 187.460 98.880 187.780 ;
        RECT 99.140 187.100 99.280 189.500 ;
        RECT 96.320 186.780 96.580 187.100 ;
        RECT 99.080 186.780 99.340 187.100 ;
        RECT 96.380 179.620 96.520 186.780 ;
        RECT 97.460 186.245 99.000 186.615 ;
        RECT 99.600 185.400 99.740 203.100 ;
        RECT 100.460 201.060 100.720 201.380 ;
        RECT 100.520 199.680 100.660 201.060 ;
        RECT 101.840 200.380 102.100 200.700 ;
        RECT 100.460 199.360 100.720 199.680 ;
        RECT 100.000 199.020 100.260 199.340 ;
        RECT 101.380 199.195 101.640 199.340 ;
        RECT 100.060 196.960 100.200 199.020 ;
        RECT 101.370 198.825 101.650 199.195 ;
        RECT 101.900 198.660 102.040 200.380 ;
        RECT 106.440 198.680 106.700 199.000 ;
        RECT 101.840 198.340 102.100 198.660 ;
        RECT 106.500 196.960 106.640 198.680 ;
        RECT 100.000 196.640 100.260 196.960 ;
        RECT 104.600 196.640 104.860 196.960 ;
        RECT 106.440 196.640 106.700 196.960 ;
        RECT 104.660 195.260 104.800 196.640 ;
        RECT 106.440 195.280 106.700 195.600 ;
        RECT 100.920 194.940 101.180 195.260 ;
        RECT 102.300 194.940 102.560 195.260 ;
        RECT 104.600 194.940 104.860 195.260 ;
        RECT 105.520 194.940 105.780 195.260 ;
        RECT 100.980 193.560 101.120 194.940 ;
        RECT 102.360 194.240 102.500 194.940 ;
        RECT 102.300 193.920 102.560 194.240 ;
        RECT 101.440 193.560 102.960 193.640 ;
        RECT 100.920 193.240 101.180 193.560 ;
        RECT 101.380 193.500 102.960 193.560 ;
        RECT 101.380 193.240 101.640 193.500 ;
        RECT 100.000 192.220 100.260 192.540 ;
        RECT 100.460 192.220 100.720 192.540 ;
        RECT 100.060 188.120 100.200 192.220 ;
        RECT 100.520 188.120 100.660 192.220 ;
        RECT 100.000 187.800 100.260 188.120 ;
        RECT 100.460 187.800 100.720 188.120 ;
        RECT 100.980 188.030 101.120 193.240 ;
        RECT 102.300 192.900 102.560 193.220 ;
        RECT 102.360 190.840 102.500 192.900 ;
        RECT 102.300 190.520 102.560 190.840 ;
        RECT 102.360 188.120 102.500 190.520 ;
        RECT 102.820 188.120 102.960 193.500 ;
        RECT 103.220 190.180 103.480 190.500 ;
        RECT 101.840 188.030 102.100 188.120 ;
        RECT 100.980 187.890 102.100 188.030 ;
        RECT 101.840 187.800 102.100 187.890 ;
        RECT 102.300 187.800 102.560 188.120 ;
        RECT 102.760 187.800 103.020 188.120 ;
        RECT 99.540 185.080 99.800 185.400 ;
        RECT 99.080 184.400 99.340 184.720 ;
        RECT 96.780 181.340 97.040 181.660 ;
        RECT 96.840 179.960 96.980 181.340 ;
        RECT 97.460 180.805 99.000 181.175 ;
        RECT 99.140 180.210 99.280 184.400 ;
        RECT 98.680 180.070 99.280 180.210 ;
        RECT 96.780 179.640 97.040 179.960 ;
        RECT 96.320 179.300 96.580 179.620 ;
        RECT 96.380 177.240 96.520 179.300 ;
        RECT 96.840 177.240 96.980 179.640 ;
        RECT 98.680 179.620 98.820 180.070 ;
        RECT 98.620 179.300 98.880 179.620 ;
        RECT 96.320 176.920 96.580 177.240 ;
        RECT 96.780 176.920 97.040 177.240 ;
        RECT 97.460 175.365 99.000 175.735 ;
        RECT 99.080 173.180 99.340 173.500 ;
        RECT 97.460 169.925 99.000 170.295 ;
        RECT 95.400 169.100 95.660 169.420 ;
        RECT 99.140 169.160 99.280 173.180 ;
        RECT 99.540 170.460 99.800 170.780 ;
        RECT 98.220 169.020 99.280 169.160 ;
        RECT 98.220 168.740 98.360 169.020 ;
        RECT 95.400 168.420 95.660 168.740 ;
        RECT 96.780 168.420 97.040 168.740 ;
        RECT 98.160 168.420 98.420 168.740 ;
        RECT 98.620 168.420 98.880 168.740 ;
        RECT 95.460 166.700 95.600 168.420 ;
        RECT 95.400 166.380 95.660 166.700 ;
        RECT 95.860 166.040 96.120 166.360 ;
        RECT 96.320 166.040 96.580 166.360 ;
        RECT 95.400 165.020 95.660 165.340 ;
        RECT 93.560 162.980 93.820 163.300 ;
        RECT 92.180 160.600 92.440 160.920 ;
        RECT 93.560 160.260 93.820 160.580 ;
        RECT 93.100 159.580 93.360 159.900 ;
        RECT 91.720 157.880 91.980 158.200 ;
        RECT 92.640 157.880 92.900 158.200 ;
        RECT 88.040 157.540 88.300 157.860 ;
        RECT 92.700 157.715 92.840 157.880 ;
        RECT 87.580 157.200 87.840 157.520 ;
        RECT 87.640 155.480 87.780 157.200 ;
        RECT 88.100 155.480 88.240 157.540 ;
        RECT 89.420 157.200 89.680 157.520 ;
        RECT 90.340 157.200 90.600 157.520 ;
        RECT 92.630 157.345 92.910 157.715 ;
        RECT 89.480 155.820 89.620 157.200 ;
        RECT 89.420 155.500 89.680 155.820 ;
        RECT 90.400 155.480 90.540 157.200 ;
        RECT 91.260 155.500 91.520 155.820 ;
        RECT 87.580 155.160 87.840 155.480 ;
        RECT 88.040 155.160 88.300 155.480 ;
        RECT 90.340 155.160 90.600 155.480 ;
        RECT 91.320 154.800 91.460 155.500 ;
        RECT 91.260 154.480 91.520 154.800 ;
        RECT 88.040 154.140 88.300 154.460 ;
        RECT 87.120 152.955 87.380 153.100 ;
        RECT 87.110 152.585 87.390 152.955 ;
        RECT 88.100 152.275 88.240 154.140 ;
        RECT 91.320 152.420 91.460 154.480 ;
        RECT 88.030 151.905 88.310 152.275 ;
        RECT 91.260 152.100 91.520 152.420 ;
        RECT 86.660 146.660 86.920 146.980 ;
        RECT 88.960 146.320 89.220 146.640 ;
        RECT 89.020 145.280 89.160 146.320 ;
        RECT 86.200 144.960 86.460 145.280 ;
        RECT 88.960 144.960 89.220 145.280 ;
        RECT 93.160 144.600 93.300 159.580 ;
        RECT 93.620 158.880 93.760 160.260 ;
        RECT 93.560 158.560 93.820 158.880 ;
        RECT 95.460 158.280 95.600 165.020 ;
        RECT 95.920 163.980 96.060 166.040 ;
        RECT 96.380 164.320 96.520 166.040 ;
        RECT 96.320 164.000 96.580 164.320 ;
        RECT 95.860 163.660 96.120 163.980 ;
        RECT 96.840 160.920 96.980 168.420 ;
        RECT 98.220 167.040 98.360 168.420 ;
        RECT 98.680 167.040 98.820 168.420 ;
        RECT 98.160 166.720 98.420 167.040 ;
        RECT 98.620 166.720 98.880 167.040 ;
        RECT 97.460 164.485 99.000 164.855 ;
        RECT 99.140 163.300 99.280 169.020 ;
        RECT 99.600 168.740 99.740 170.460 ;
        RECT 100.920 168.760 101.180 169.080 ;
        RECT 101.900 168.860 102.040 187.800 ;
        RECT 102.290 187.520 102.570 187.635 ;
        RECT 102.820 187.520 102.960 187.800 ;
        RECT 102.290 187.380 102.960 187.520 ;
        RECT 102.290 187.265 102.570 187.380 ;
        RECT 103.280 187.100 103.420 190.180 ;
        RECT 103.680 187.800 103.940 188.120 ;
        RECT 103.220 186.780 103.480 187.100 ;
        RECT 103.280 185.740 103.420 186.780 ;
        RECT 103.740 186.080 103.880 187.800 ;
        RECT 104.140 186.780 104.400 187.100 ;
        RECT 103.680 185.760 103.940 186.080 ;
        RECT 103.220 185.420 103.480 185.740 ;
        RECT 104.200 185.400 104.340 186.780 ;
        RECT 104.140 185.080 104.400 185.400 ;
        RECT 103.680 184.740 103.940 185.060 ;
        RECT 102.760 182.700 103.020 183.020 ;
        RECT 102.300 182.020 102.560 182.340 ;
        RECT 99.540 168.420 99.800 168.740 ;
        RECT 100.000 168.420 100.260 168.740 ;
        RECT 100.060 166.700 100.200 168.420 ;
        RECT 100.000 166.380 100.260 166.700 ;
        RECT 99.080 162.980 99.340 163.300 ;
        RECT 100.000 162.640 100.260 162.960 ;
        RECT 96.780 160.600 97.040 160.920 ;
        RECT 97.460 159.045 99.000 159.415 ;
        RECT 95.460 158.140 96.520 158.280 ;
        RECT 95.400 157.540 95.660 157.860 ;
        RECT 94.480 154.820 94.740 155.140 ;
        RECT 93.560 152.100 93.820 152.420 ;
        RECT 94.020 152.330 94.280 152.420 ;
        RECT 94.540 152.330 94.680 154.820 ;
        RECT 94.940 154.480 95.200 154.800 ;
        RECT 94.020 152.190 94.680 152.330 ;
        RECT 94.020 152.100 94.280 152.190 ;
        RECT 93.620 150.040 93.760 152.100 ;
        RECT 94.540 150.040 94.680 152.190 ;
        RECT 95.000 150.720 95.140 154.480 ;
        RECT 95.460 153.440 95.600 157.540 ;
        RECT 95.860 156.860 96.120 157.180 ;
        RECT 95.920 156.160 96.060 156.860 ;
        RECT 95.860 155.840 96.120 156.160 ;
        RECT 95.860 154.820 96.120 155.140 ;
        RECT 95.400 153.120 95.660 153.440 ;
        RECT 95.920 152.420 96.060 154.820 ;
        RECT 96.380 154.460 96.520 158.140 ;
        RECT 99.080 157.880 99.340 158.200 ;
        RECT 98.160 157.540 98.420 157.860 ;
        RECT 98.220 156.160 98.360 157.540 ;
        RECT 98.160 155.840 98.420 156.160 ;
        RECT 96.320 154.140 96.580 154.460 ;
        RECT 95.860 152.100 96.120 152.420 ;
        RECT 96.380 151.740 96.520 154.140 ;
        RECT 97.460 153.605 99.000 153.975 ;
        RECT 98.160 153.120 98.420 153.440 ;
        RECT 97.230 152.585 97.510 152.955 ;
        RECT 97.300 151.740 97.440 152.585 ;
        RECT 97.700 152.275 97.960 152.420 ;
        RECT 97.690 151.905 97.970 152.275 ;
        RECT 96.320 151.420 96.580 151.740 ;
        RECT 97.240 151.420 97.500 151.740 ;
        RECT 98.220 150.720 98.360 153.120 ;
        RECT 94.940 150.400 95.200 150.720 ;
        RECT 98.160 150.400 98.420 150.720 ;
        RECT 93.560 149.720 93.820 150.040 ;
        RECT 94.480 149.720 94.740 150.040 ;
        RECT 93.620 146.640 93.760 149.720 ;
        RECT 94.540 147.660 94.680 149.720 ;
        RECT 95.000 149.020 95.140 150.400 ;
        RECT 99.140 149.700 99.280 157.880 ;
        RECT 99.080 149.380 99.340 149.700 ;
        RECT 94.940 148.700 95.200 149.020 ;
        RECT 94.480 147.340 94.740 147.660 ;
        RECT 93.560 146.320 93.820 146.640 ;
        RECT 95.000 145.280 95.140 148.700 ;
        RECT 97.460 148.165 99.000 148.535 ;
        RECT 100.060 147.320 100.200 162.640 ;
        RECT 100.980 152.420 101.120 168.760 ;
        RECT 101.440 168.720 102.040 168.860 ;
        RECT 101.440 157.860 101.580 168.720 ;
        RECT 101.840 161.280 102.100 161.600 ;
        RECT 101.900 158.200 102.040 161.280 ;
        RECT 101.840 157.880 102.100 158.200 ;
        RECT 101.380 157.540 101.640 157.860 ;
        RECT 101.380 156.860 101.640 157.180 ;
        RECT 101.440 154.460 101.580 156.860 ;
        RECT 101.900 156.160 102.040 157.880 ;
        RECT 101.840 155.840 102.100 156.160 ;
        RECT 101.840 155.160 102.100 155.480 ;
        RECT 101.380 154.140 101.640 154.460 ;
        RECT 100.920 152.100 101.180 152.420 ;
        RECT 101.900 149.700 102.040 155.160 ;
        RECT 102.360 153.440 102.500 182.020 ;
        RECT 102.820 180.640 102.960 182.700 ;
        RECT 103.740 182.660 103.880 184.740 ;
        RECT 103.740 182.520 104.340 182.660 ;
        RECT 102.760 180.320 103.020 180.640 ;
        RECT 103.220 179.300 103.480 179.620 ;
        RECT 103.280 177.920 103.420 179.300 ;
        RECT 103.220 177.600 103.480 177.920 ;
        RECT 103.220 176.580 103.480 176.900 ;
        RECT 103.280 173.840 103.420 176.580 ;
        RECT 103.220 173.520 103.480 173.840 ;
        RECT 102.760 170.460 103.020 170.780 ;
        RECT 102.820 167.040 102.960 170.460 ;
        RECT 102.760 166.720 103.020 167.040 ;
        RECT 104.200 166.270 104.340 182.520 ;
        RECT 104.660 176.220 104.800 194.940 ;
        RECT 105.060 185.420 105.320 185.740 ;
        RECT 105.120 179.620 105.260 185.420 ;
        RECT 105.580 182.680 105.720 194.940 ;
        RECT 106.500 193.220 106.640 195.280 ;
        RECT 106.440 192.900 106.700 193.220 ;
        RECT 105.520 182.360 105.780 182.680 ;
        RECT 105.060 179.300 105.320 179.620 ;
        RECT 104.600 175.900 104.860 176.220 ;
        RECT 104.660 166.360 104.800 175.900 ;
        RECT 105.120 175.200 105.260 179.300 ;
        RECT 106.500 179.190 106.640 192.900 ;
        RECT 106.960 183.360 107.100 203.440 ;
        RECT 110.180 201.380 110.320 205.820 ;
        RECT 110.640 203.420 110.780 206.500 ;
        RECT 110.580 203.100 110.840 203.420 ;
        RECT 110.640 201.720 110.780 203.100 ;
        RECT 110.580 201.400 110.840 201.720 ;
        RECT 108.280 201.060 108.540 201.380 ;
        RECT 110.120 201.060 110.380 201.380 ;
        RECT 108.340 197.980 108.480 201.060 ;
        RECT 108.280 197.660 108.540 197.980 ;
        RECT 108.340 191.520 108.480 197.660 ;
        RECT 111.560 195.260 111.700 208.880 ;
        RECT 111.960 208.540 112.220 208.860 ;
        RECT 112.880 208.540 113.140 208.860 ;
        RECT 111.500 194.940 111.760 195.260 ;
        RECT 110.120 193.240 110.380 193.560 ;
        RECT 108.280 191.200 108.540 191.520 ;
        RECT 109.660 185.420 109.920 185.740 ;
        RECT 109.720 184.720 109.860 185.420 ;
        RECT 110.180 184.970 110.320 193.240 ;
        RECT 111.040 192.900 111.300 193.220 ;
        RECT 111.100 191.520 111.240 192.900 ;
        RECT 111.040 191.200 111.300 191.520 ;
        RECT 112.020 185.740 112.160 208.540 ;
        RECT 112.940 206.820 113.080 208.540 ;
        RECT 122.600 207.840 122.740 209.560 ;
        RECT 123.000 208.540 123.260 208.860 ;
        RECT 122.540 207.520 122.800 207.840 ;
        RECT 112.880 206.500 113.140 206.820 ;
        RECT 114.880 205.285 116.420 205.655 ;
        RECT 112.420 204.120 112.680 204.440 ;
        RECT 112.480 202.400 112.620 204.120 ;
        RECT 112.420 202.080 112.680 202.400 ;
        RECT 123.060 201.380 123.200 208.540 ;
        RECT 124.900 207.840 125.040 209.560 ;
        RECT 124.840 207.520 125.100 207.840 ;
        RECT 127.660 206.820 127.800 211.260 ;
        RECT 130.360 208.540 130.620 208.860 ;
        RECT 130.420 207.840 130.560 208.540 ;
        RECT 132.305 208.005 133.845 208.375 ;
        RECT 130.360 207.520 130.620 207.840 ;
        RECT 127.600 206.500 127.860 206.820 ;
        RECT 137.780 206.480 137.920 211.260 ;
        RECT 127.140 206.160 127.400 206.480 ;
        RECT 137.720 206.160 137.980 206.480 ;
        RECT 123.000 201.060 123.260 201.380 ;
        RECT 117.020 200.720 117.280 201.040 ;
        RECT 114.880 199.845 116.420 200.215 ;
        RECT 117.080 199.680 117.220 200.720 ;
        RECT 121.620 200.380 121.880 200.700 ;
        RECT 117.020 199.360 117.280 199.680 ;
        RECT 115.640 198.680 115.900 199.000 ;
        RECT 113.340 197.660 113.600 197.980 ;
        RECT 112.420 195.960 112.680 196.280 ;
        RECT 112.480 190.840 112.620 195.960 ;
        RECT 113.400 192.880 113.540 197.660 ;
        RECT 115.700 196.960 115.840 198.680 ;
        RECT 121.680 196.960 121.820 200.380 ;
        RECT 124.380 198.340 124.640 198.660 ;
        RECT 123.000 197.660 123.260 197.980 ;
        RECT 115.640 196.640 115.900 196.960 ;
        RECT 121.620 196.640 121.880 196.960 ;
        RECT 118.400 195.960 118.660 196.280 ;
        RECT 117.480 195.620 117.740 195.940 ;
        RECT 113.800 194.940 114.060 195.260 ;
        RECT 113.340 192.560 113.600 192.880 ;
        RECT 112.420 190.520 112.680 190.840 ;
        RECT 113.400 190.500 113.540 192.560 ;
        RECT 113.340 190.180 113.600 190.500 ;
        RECT 113.400 188.800 113.540 190.180 ;
        RECT 113.340 188.480 113.600 188.800 ;
        RECT 112.420 185.760 112.680 186.080 ;
        RECT 111.960 185.420 112.220 185.740 ;
        RECT 111.040 184.970 111.300 185.060 ;
        RECT 110.180 184.830 111.300 184.970 ;
        RECT 109.660 184.400 109.920 184.720 ;
        RECT 106.900 183.040 107.160 183.360 ;
        RECT 109.720 182.680 109.860 184.400 ;
        RECT 109.660 182.360 109.920 182.680 ;
        RECT 109.720 181.660 109.860 182.360 ;
        RECT 110.180 182.000 110.320 184.830 ;
        RECT 111.040 184.740 111.300 184.830 ;
        RECT 111.040 184.060 111.300 184.380 ;
        RECT 111.100 182.680 111.240 184.060 ;
        RECT 111.040 182.360 111.300 182.680 ;
        RECT 110.120 181.680 110.380 182.000 ;
        RECT 109.660 181.340 109.920 181.660 ;
        RECT 106.900 179.190 107.160 179.280 ;
        RECT 106.500 179.050 107.160 179.190 ;
        RECT 106.900 178.960 107.160 179.050 ;
        RECT 108.280 178.960 108.540 179.280 ;
        RECT 105.980 178.850 106.240 178.940 ;
        RECT 105.580 178.710 106.240 178.850 ;
        RECT 105.580 176.900 105.720 178.710 ;
        RECT 105.980 178.620 106.240 178.710 ;
        RECT 105.980 177.260 106.240 177.580 ;
        RECT 105.520 176.580 105.780 176.900 ;
        RECT 106.040 175.200 106.180 177.260 ;
        RECT 106.960 177.240 107.100 178.960 ;
        RECT 108.340 177.580 108.480 178.960 ;
        RECT 109.720 178.940 109.860 181.340 ;
        RECT 110.120 179.300 110.380 179.620 ;
        RECT 109.660 178.620 109.920 178.940 ;
        RECT 108.280 177.260 108.540 177.580 ;
        RECT 109.720 177.240 109.860 178.620 ;
        RECT 106.900 176.920 107.160 177.240 ;
        RECT 108.740 176.920 109.000 177.240 ;
        RECT 109.660 176.920 109.920 177.240 ;
        RECT 108.800 176.220 108.940 176.920 ;
        RECT 108.740 175.900 109.000 176.220 ;
        RECT 105.060 174.880 105.320 175.200 ;
        RECT 105.980 174.880 106.240 175.200 ;
        RECT 105.120 171.460 105.260 174.880 ;
        RECT 105.060 171.140 105.320 171.460 ;
        RECT 108.740 171.140 109.000 171.460 ;
        RECT 108.800 169.760 108.940 171.140 ;
        RECT 108.740 169.440 109.000 169.760 ;
        RECT 109.200 168.760 109.460 169.080 ;
        RECT 103.740 166.130 104.340 166.270 ;
        RECT 103.220 157.880 103.480 158.200 ;
        RECT 102.300 153.120 102.560 153.440 ;
        RECT 101.840 149.380 102.100 149.700 ;
        RECT 102.300 147.340 102.560 147.660 ;
        RECT 100.000 147.000 100.260 147.320 ;
        RECT 100.000 145.980 100.260 146.300 ;
        RECT 94.940 144.960 95.200 145.280 ;
        RECT 93.100 144.280 93.360 144.600 ;
        RECT 83.440 143.260 83.700 143.580 ;
        RECT 87.580 143.260 87.840 143.580 ;
        RECT 86.200 139.180 86.460 139.500 ;
        RECT 84.360 138.840 84.620 139.160 ;
        RECT 83.440 137.820 83.700 138.140 ;
        RECT 83.500 136.100 83.640 137.820 ;
        RECT 84.420 136.440 84.560 138.840 ;
        RECT 86.260 138.140 86.400 139.180 ;
        RECT 87.640 139.160 87.780 143.260 ;
        RECT 97.460 142.725 99.000 143.095 ;
        RECT 94.480 141.560 94.740 141.880 ;
        RECT 89.880 139.520 90.140 139.840 ;
        RECT 89.940 139.160 90.080 139.520 ;
        RECT 87.580 138.840 87.840 139.160 ;
        RECT 89.420 138.840 89.680 139.160 ;
        RECT 89.880 138.840 90.140 139.160 ;
        RECT 86.200 137.820 86.460 138.140 ;
        RECT 88.960 137.820 89.220 138.140 ;
        RECT 89.020 136.440 89.160 137.820 ;
        RECT 84.360 136.120 84.620 136.440 ;
        RECT 88.960 136.120 89.220 136.440 ;
        RECT 83.440 135.780 83.700 136.100 ;
        RECT 84.820 135.840 85.080 136.100 ;
        RECT 83.960 135.780 85.080 135.840 ;
        RECT 83.960 135.700 85.020 135.780 ;
        RECT 83.960 135.420 84.100 135.700 ;
        RECT 82.580 135.020 83.180 135.160 ;
        RECT 82.060 130.340 82.320 130.660 ;
        RECT 79.300 130.000 79.560 130.320 ;
        RECT 79.360 128.960 79.500 130.000 ;
        RECT 80.035 129.125 81.575 129.495 ;
        RECT 82.580 128.960 82.720 135.020 ;
        RECT 83.430 134.905 83.710 135.275 ;
        RECT 83.900 135.100 84.160 135.420 ;
        RECT 84.360 135.100 84.620 135.420 ;
        RECT 82.980 132.380 83.240 132.700 ;
        RECT 83.040 131.680 83.180 132.380 ;
        RECT 82.980 131.360 83.240 131.680 ;
        RECT 79.300 128.640 79.560 128.960 ;
        RECT 82.520 128.640 82.780 128.960 ;
        RECT 78.840 128.300 79.100 128.620 ;
        RECT 82.580 128.280 82.720 128.640 ;
        RECT 83.500 128.280 83.640 134.905 ;
        RECT 84.420 131.340 84.560 135.100 ;
        RECT 89.480 134.360 89.620 138.840 ;
        RECT 92.180 138.160 92.440 138.480 ;
        RECT 89.870 136.265 90.150 136.635 ;
        RECT 89.940 136.100 90.080 136.265 ;
        RECT 89.880 135.780 90.140 136.100 ;
        RECT 92.240 135.420 92.380 138.160 ;
        RECT 93.560 137.820 93.820 138.140 ;
        RECT 93.620 136.100 93.760 137.820 ;
        RECT 94.540 136.440 94.680 141.560 ;
        RECT 100.060 141.540 100.200 145.980 ;
        RECT 102.360 143.920 102.500 147.340 ;
        RECT 103.280 144.940 103.420 157.880 ;
        RECT 103.740 150.040 103.880 166.130 ;
        RECT 104.600 166.040 104.860 166.360 ;
        RECT 107.820 165.020 108.080 165.340 ;
        RECT 107.880 164.320 108.020 165.020 ;
        RECT 107.820 164.000 108.080 164.320 ;
        RECT 106.440 162.300 106.700 162.620 ;
        RECT 106.500 161.600 106.640 162.300 ;
        RECT 106.440 161.280 106.700 161.600 ;
        RECT 105.060 158.220 105.320 158.540 ;
        RECT 105.120 150.040 105.260 158.220 ;
        RECT 109.260 157.180 109.400 168.760 ;
        RECT 110.180 157.860 110.320 179.300 ;
        RECT 111.100 174.180 111.240 182.360 ;
        RECT 111.960 179.640 112.220 179.960 ;
        RECT 111.040 173.860 111.300 174.180 ;
        RECT 110.580 167.740 110.840 168.060 ;
        RECT 110.640 166.020 110.780 167.740 ;
        RECT 111.100 166.360 111.240 173.860 ;
        RECT 112.020 169.420 112.160 179.640 ;
        RECT 112.480 177.920 112.620 185.760 ;
        RECT 113.340 184.740 113.600 185.060 ;
        RECT 113.400 183.360 113.540 184.740 ;
        RECT 113.340 183.040 113.600 183.360 ;
        RECT 113.860 182.875 114.000 194.940 ;
        RECT 114.880 194.405 116.420 194.775 ;
        RECT 116.560 193.240 116.820 193.560 ;
        RECT 116.620 190.840 116.760 193.240 ;
        RECT 117.540 192.880 117.680 195.620 ;
        RECT 118.460 193.130 118.600 195.960 ;
        RECT 121.680 195.850 121.820 196.640 ;
        RECT 121.220 195.710 121.820 195.850 ;
        RECT 120.700 193.920 120.960 194.240 ;
        RECT 119.320 193.130 119.580 193.220 ;
        RECT 118.000 192.990 119.580 193.130 ;
        RECT 117.480 192.560 117.740 192.880 ;
        RECT 116.560 190.520 116.820 190.840 ;
        RECT 114.880 188.965 116.420 189.335 ;
        RECT 116.620 188.800 116.760 190.520 ;
        RECT 118.000 190.500 118.140 192.990 ;
        RECT 119.320 192.900 119.580 192.990 ;
        RECT 120.760 192.960 120.900 193.920 ;
        RECT 121.220 193.560 121.360 195.710 ;
        RECT 121.620 194.940 121.880 195.260 ;
        RECT 121.680 194.240 121.820 194.940 ;
        RECT 121.620 193.920 121.880 194.240 ;
        RECT 121.160 193.240 121.420 193.560 ;
        RECT 120.760 192.820 121.820 192.960 ;
        RECT 120.700 192.220 120.960 192.540 ;
        RECT 120.760 190.840 120.900 192.220 ;
        RECT 120.700 190.520 120.960 190.840 ;
        RECT 117.940 190.180 118.200 190.500 ;
        RECT 120.240 190.180 120.500 190.500 ;
        RECT 116.560 188.480 116.820 188.800 ;
        RECT 118.000 188.460 118.140 190.180 ;
        RECT 117.940 188.140 118.200 188.460 ;
        RECT 117.020 187.120 117.280 187.440 ;
        RECT 114.260 185.420 114.520 185.740 ;
        RECT 113.790 182.505 114.070 182.875 ;
        RECT 113.340 182.020 113.600 182.340 ;
        RECT 113.400 179.620 113.540 182.020 ;
        RECT 113.860 180.640 114.000 182.505 ;
        RECT 113.800 180.320 114.060 180.640 ;
        RECT 113.340 179.300 113.600 179.620 ;
        RECT 112.420 177.600 112.680 177.920 ;
        RECT 113.400 176.640 113.540 179.300 ;
        RECT 112.480 176.500 113.540 176.640 ;
        RECT 111.960 169.100 112.220 169.420 ;
        RECT 112.480 166.700 112.620 176.500 ;
        RECT 112.880 175.900 113.140 176.220 ;
        RECT 112.940 175.200 113.080 175.900 ;
        RECT 114.320 175.200 114.460 185.420 ;
        RECT 116.560 184.060 116.820 184.380 ;
        RECT 114.880 183.525 116.420 183.895 ;
        RECT 116.620 182.000 116.760 184.060 ;
        RECT 117.080 183.020 117.220 187.120 ;
        RECT 117.480 186.780 117.740 187.100 ;
        RECT 117.020 182.700 117.280 183.020 ;
        RECT 116.560 181.680 116.820 182.000 ;
        RECT 116.620 179.620 116.760 181.680 ;
        RECT 117.080 181.660 117.220 182.700 ;
        RECT 117.020 181.340 117.280 181.660 ;
        RECT 116.560 179.300 116.820 179.620 ;
        RECT 114.880 178.085 116.420 178.455 ;
        RECT 117.020 177.260 117.280 177.580 ;
        RECT 112.880 174.880 113.140 175.200 ;
        RECT 114.260 174.880 114.520 175.200 ;
        RECT 113.340 173.860 113.600 174.180 ;
        RECT 113.400 172.480 113.540 173.860 ;
        RECT 113.340 172.160 113.600 172.480 ;
        RECT 113.400 168.740 113.540 172.160 ;
        RECT 114.320 171.800 114.460 174.880 ;
        RECT 117.080 174.180 117.220 177.260 ;
        RECT 117.540 177.240 117.680 186.780 ;
        RECT 120.300 186.080 120.440 190.180 ;
        RECT 121.680 189.820 121.820 192.820 ;
        RECT 121.160 189.500 121.420 189.820 ;
        RECT 121.620 189.500 121.880 189.820 ;
        RECT 120.240 185.760 120.500 186.080 ;
        RECT 119.320 185.080 119.580 185.400 ;
        RECT 118.860 184.060 119.120 184.380 ;
        RECT 118.920 183.020 119.060 184.060 ;
        RECT 118.860 182.700 119.120 183.020 ;
        RECT 119.380 179.620 119.520 185.080 ;
        RECT 121.220 185.060 121.360 189.500 ;
        RECT 121.680 186.160 121.820 189.500 ;
        RECT 123.060 188.315 123.200 197.660 ;
        RECT 124.440 193.560 124.580 198.340 ;
        RECT 124.380 193.470 124.640 193.560 ;
        RECT 124.380 193.330 125.040 193.470 ;
        RECT 124.380 193.240 124.640 193.330 ;
        RECT 123.920 192.560 124.180 192.880 ;
        RECT 122.990 187.945 123.270 188.315 ;
        RECT 121.680 186.020 122.280 186.160 ;
        RECT 121.620 185.080 121.880 185.400 ;
        RECT 121.160 184.740 121.420 185.060 ;
        RECT 119.780 184.060 120.040 184.380 ;
        RECT 119.840 183.020 119.980 184.060 ;
        RECT 121.220 183.360 121.360 184.740 ;
        RECT 121.160 183.040 121.420 183.360 ;
        RECT 119.780 182.700 120.040 183.020 ;
        RECT 119.840 180.300 119.980 182.700 ;
        RECT 121.680 182.680 121.820 185.080 ;
        RECT 121.620 182.360 121.880 182.680 ;
        RECT 120.700 182.020 120.960 182.340 ;
        RECT 119.780 179.980 120.040 180.300 ;
        RECT 119.320 179.300 119.580 179.620 ;
        RECT 117.940 178.620 118.200 178.940 ;
        RECT 117.480 176.920 117.740 177.240 ;
        RECT 117.540 175.200 117.680 176.920 ;
        RECT 117.480 174.880 117.740 175.200 ;
        RECT 118.000 174.600 118.140 178.620 ;
        RECT 120.760 176.560 120.900 182.020 ;
        RECT 121.680 179.960 121.820 182.360 ;
        RECT 122.140 180.640 122.280 186.020 ;
        RECT 123.980 184.720 124.120 192.560 ;
        RECT 124.380 192.220 124.640 192.540 ;
        RECT 124.440 190.500 124.580 192.220 ;
        RECT 124.380 190.180 124.640 190.500 ;
        RECT 124.900 185.400 125.040 193.330 ;
        RECT 126.220 193.240 126.480 193.560 ;
        RECT 126.280 191.520 126.420 193.240 ;
        RECT 126.220 191.200 126.480 191.520 ;
        RECT 125.300 190.180 125.560 190.500 ;
        RECT 124.840 185.080 125.100 185.400 ;
        RECT 123.920 184.400 124.180 184.720 ;
        RECT 123.000 182.360 123.260 182.680 ;
        RECT 123.060 181.660 123.200 182.360 ;
        RECT 123.000 181.340 123.260 181.660 ;
        RECT 122.080 180.320 122.340 180.640 ;
        RECT 122.540 180.320 122.800 180.640 ;
        RECT 121.620 179.640 121.880 179.960 ;
        RECT 122.140 177.920 122.280 180.320 ;
        RECT 122.080 177.600 122.340 177.920 ;
        RECT 122.600 177.580 122.740 180.320 ;
        RECT 123.060 179.960 123.200 181.340 ;
        RECT 123.000 179.640 123.260 179.960 ;
        RECT 123.460 178.620 123.720 178.940 ;
        RECT 122.540 177.260 122.800 177.580 ;
        RECT 123.520 177.240 123.660 178.620 ;
        RECT 123.460 176.920 123.720 177.240 ;
        RECT 120.700 176.240 120.960 176.560 ;
        RECT 119.320 175.900 119.580 176.220 ;
        RECT 119.380 175.200 119.520 175.900 ;
        RECT 119.320 174.880 119.580 175.200 ;
        RECT 117.540 174.460 118.140 174.600 ;
        RECT 117.020 173.860 117.280 174.180 ;
        RECT 116.560 173.180 116.820 173.500 ;
        RECT 114.880 172.645 116.420 173.015 ;
        RECT 116.620 171.800 116.760 173.180 ;
        RECT 114.260 171.480 114.520 171.800 ;
        RECT 116.560 171.480 116.820 171.800 ;
        RECT 113.340 168.420 113.600 168.740 ;
        RECT 114.320 168.060 114.460 171.480 ;
        RECT 114.720 170.460 114.980 170.780 ;
        RECT 114.780 169.760 114.920 170.460 ;
        RECT 114.720 169.440 114.980 169.760 ;
        RECT 116.100 168.595 116.360 168.740 ;
        RECT 116.090 168.225 116.370 168.595 ;
        RECT 117.540 168.310 117.680 174.460 ;
        RECT 120.760 174.180 120.900 176.240 ;
        RECT 118.860 173.860 119.120 174.180 ;
        RECT 120.700 173.860 120.960 174.180 ;
        RECT 118.920 172.480 119.060 173.860 ;
        RECT 118.860 172.160 119.120 172.480 ;
        RECT 117.940 171.820 118.200 172.140 ;
        RECT 118.000 168.860 118.140 171.820 ;
        RECT 118.920 169.760 119.060 172.160 ;
        RECT 119.780 171.480 120.040 171.800 ;
        RECT 118.860 169.440 119.120 169.760 ;
        RECT 118.000 168.740 119.060 168.860 ;
        RECT 119.840 168.740 119.980 171.480 ;
        RECT 118.000 168.720 119.120 168.740 ;
        RECT 118.860 168.420 119.120 168.720 ;
        RECT 119.780 168.420 120.040 168.740 ;
        RECT 117.940 168.310 118.200 168.400 ;
        RECT 117.540 168.170 118.200 168.310 ;
        RECT 117.940 168.080 118.200 168.170 ;
        RECT 114.260 167.740 114.520 168.060 ;
        RECT 116.560 167.740 116.820 168.060 ;
        RECT 114.880 167.205 116.420 167.575 ;
        RECT 116.620 167.040 116.760 167.740 ;
        RECT 116.560 166.720 116.820 167.040 ;
        RECT 112.420 166.380 112.680 166.700 ;
        RECT 111.040 166.040 111.300 166.360 ;
        RECT 118.000 166.020 118.140 168.080 ;
        RECT 110.580 165.700 110.840 166.020 ;
        RECT 111.960 165.700 112.220 166.020 ;
        RECT 117.940 165.700 118.200 166.020 ;
        RECT 111.040 165.360 111.300 165.680 ;
        RECT 110.120 157.540 110.380 157.860 ;
        RECT 109.200 156.860 109.460 157.180 ;
        RECT 109.260 155.480 109.400 156.860 ;
        RECT 107.820 155.160 108.080 155.480 ;
        RECT 109.200 155.160 109.460 155.480 ;
        RECT 105.520 154.820 105.780 155.140 ;
        RECT 103.680 149.720 103.940 150.040 ;
        RECT 105.060 149.720 105.320 150.040 ;
        RECT 103.680 148.700 103.940 149.020 ;
        RECT 103.220 144.620 103.480 144.940 ;
        RECT 102.300 143.600 102.560 143.920 ;
        RECT 100.000 141.220 100.260 141.540 ;
        RECT 102.360 139.500 102.500 143.600 ;
        RECT 103.280 141.880 103.420 144.620 ;
        RECT 103.740 144.600 103.880 148.700 ;
        RECT 103.680 144.280 103.940 144.600 ;
        RECT 103.220 141.560 103.480 141.880 ;
        RECT 102.760 140.540 103.020 140.860 ;
        RECT 96.780 139.180 97.040 139.500 ;
        RECT 102.300 139.180 102.560 139.500 ;
        RECT 96.840 137.120 96.980 139.180 ;
        RECT 98.620 138.560 98.880 138.820 ;
        RECT 98.620 138.500 99.280 138.560 ;
        RECT 101.380 138.500 101.640 138.820 ;
        RECT 98.680 138.420 99.280 138.500 ;
        RECT 97.460 137.285 99.000 137.655 ;
        RECT 96.780 136.800 97.040 137.120 ;
        RECT 96.320 136.460 96.580 136.780 ;
        RECT 94.480 136.120 94.740 136.440 ;
        RECT 93.560 135.780 93.820 136.100 ;
        RECT 94.540 135.420 94.680 136.120 ;
        RECT 92.180 135.100 92.440 135.420 ;
        RECT 94.480 135.100 94.740 135.420 ;
        RECT 89.020 134.220 89.620 134.360 ;
        RECT 89.020 134.060 89.160 134.220 ;
        RECT 88.960 133.740 89.220 134.060 ;
        RECT 84.360 131.020 84.620 131.340 ;
        RECT 85.280 130.340 85.540 130.660 ;
        RECT 84.820 130.000 85.080 130.320 ;
        RECT 84.880 128.960 85.020 130.000 ;
        RECT 85.340 129.980 85.480 130.340 ;
        RECT 85.280 129.660 85.540 129.980 ;
        RECT 86.200 129.660 86.460 129.980 ;
        RECT 84.820 128.640 85.080 128.960 ;
        RECT 85.340 128.620 85.480 129.660 ;
        RECT 86.260 128.960 86.400 129.660 ;
        RECT 86.200 128.640 86.460 128.960 ;
        RECT 85.280 128.300 85.540 128.620 ;
        RECT 67.340 127.960 67.600 128.280 ;
        RECT 82.520 127.960 82.780 128.280 ;
        RECT 83.440 127.960 83.700 128.280 ;
        RECT 67.400 126.240 67.540 127.960 ;
        RECT 82.580 127.600 82.720 127.960 ;
        RECT 82.520 127.280 82.780 127.600 ;
        RECT 89.020 127.260 89.160 133.740 ;
        RECT 90.340 132.380 90.600 132.700 ;
        RECT 89.420 129.660 89.680 129.980 ;
        RECT 89.480 128.960 89.620 129.660 ;
        RECT 89.420 128.640 89.680 128.960 ;
        RECT 90.400 128.620 90.540 132.380 ;
        RECT 90.340 128.300 90.600 128.620 ;
        RECT 92.640 127.620 92.900 127.940 ;
        RECT 88.960 126.940 89.220 127.260 ;
        RECT 91.260 126.940 91.520 127.260 ;
        RECT 67.340 125.920 67.600 126.240 ;
        RECT 91.320 125.560 91.460 126.940 ;
        RECT 92.700 126.240 92.840 127.620 ;
        RECT 92.640 125.920 92.900 126.240 ;
        RECT 66.420 125.240 66.680 125.560 ;
        RECT 91.260 125.240 91.520 125.560 ;
        RECT 96.380 125.220 96.520 136.460 ;
        RECT 97.460 131.845 99.000 132.215 ;
        RECT 99.140 131.680 99.280 138.420 ;
        RECT 101.440 133.720 101.580 138.500 ;
        RECT 101.380 133.400 101.640 133.720 ;
        RECT 99.080 131.360 99.340 131.680 ;
        RECT 99.140 128.280 99.280 131.360 ;
        RECT 102.360 130.660 102.500 139.180 ;
        RECT 102.820 138.820 102.960 140.540 ;
        RECT 102.760 138.500 103.020 138.820 ;
        RECT 103.280 138.480 103.420 141.560 ;
        RECT 103.740 141.540 103.880 144.280 ;
        RECT 105.060 143.260 105.320 143.580 ;
        RECT 105.120 142.560 105.260 143.260 ;
        RECT 105.060 142.240 105.320 142.560 ;
        RECT 105.580 141.960 105.720 154.820 ;
        RECT 107.880 150.040 108.020 155.160 ;
        RECT 108.740 154.140 109.000 154.460 ;
        RECT 108.800 150.720 108.940 154.140 ;
        RECT 111.100 153.100 111.240 165.360 ;
        RECT 112.020 161.600 112.160 165.700 ;
        RECT 119.320 165.020 119.580 165.340 ;
        RECT 114.880 161.765 116.420 162.135 ;
        RECT 111.960 161.280 112.220 161.600 ;
        RECT 114.880 156.325 116.420 156.695 ;
        RECT 111.040 152.780 111.300 153.100 ;
        RECT 109.200 151.760 109.460 152.080 ;
        RECT 109.260 150.720 109.400 151.760 ;
        RECT 111.100 150.720 111.240 152.780 ;
        RECT 118.860 152.440 119.120 152.760 ;
        RECT 114.880 150.885 116.420 151.255 ;
        RECT 108.740 150.400 109.000 150.720 ;
        RECT 109.200 150.400 109.460 150.720 ;
        RECT 111.040 150.400 111.300 150.720 ;
        RECT 107.820 149.720 108.080 150.040 ;
        RECT 108.280 149.720 108.540 150.040 ;
        RECT 108.340 148.000 108.480 149.720 ;
        RECT 109.660 148.700 109.920 149.020 ;
        RECT 110.120 148.700 110.380 149.020 ;
        RECT 108.280 147.680 108.540 148.000 ;
        RECT 109.720 147.660 109.860 148.700 ;
        RECT 109.660 147.340 109.920 147.660 ;
        RECT 105.120 141.820 105.720 141.960 ;
        RECT 103.680 141.280 103.940 141.540 ;
        RECT 103.680 141.220 104.340 141.280 ;
        RECT 103.740 141.140 104.340 141.220 ;
        RECT 103.220 138.160 103.480 138.480 ;
        RECT 104.200 133.720 104.340 141.140 ;
        RECT 105.120 139.840 105.260 141.820 ;
        RECT 105.520 141.220 105.780 141.540 ;
        RECT 105.980 141.220 106.240 141.540 ;
        RECT 107.820 141.220 108.080 141.540 ;
        RECT 105.580 140.860 105.720 141.220 ;
        RECT 105.520 140.540 105.780 140.860 ;
        RECT 105.060 139.520 105.320 139.840 ;
        RECT 105.580 139.160 105.720 140.540 ;
        RECT 106.040 139.840 106.180 141.220 ;
        RECT 107.880 139.840 108.020 141.220 ;
        RECT 109.720 140.860 109.860 147.340 ;
        RECT 110.180 141.540 110.320 148.700 ;
        RECT 110.580 146.890 110.840 146.980 ;
        RECT 111.100 146.890 111.240 150.400 ;
        RECT 113.340 150.060 113.600 150.380 ;
        RECT 111.500 149.720 111.760 150.040 ;
        RECT 111.560 147.320 111.700 149.720 ;
        RECT 111.500 147.000 111.760 147.320 ;
        RECT 113.400 146.980 113.540 150.060 ;
        RECT 114.720 149.720 114.980 150.040 ;
        RECT 114.780 148.000 114.920 149.720 ;
        RECT 116.560 148.700 116.820 149.020 ;
        RECT 114.720 147.680 114.980 148.000 ;
        RECT 110.580 146.750 111.240 146.890 ;
        RECT 110.580 146.660 110.840 146.750 ;
        RECT 113.340 146.660 113.600 146.980 ;
        RECT 116.620 146.640 116.760 148.700 ;
        RECT 117.940 146.660 118.200 146.980 ;
        RECT 111.500 146.320 111.760 146.640 ;
        RECT 116.560 146.320 116.820 146.640 ;
        RECT 111.560 141.540 111.700 146.320 ;
        RECT 114.880 145.445 116.420 145.815 ;
        RECT 116.560 144.280 116.820 144.600 ;
        RECT 110.120 141.220 110.380 141.540 ;
        RECT 111.500 141.220 111.760 141.540 ;
        RECT 108.280 140.540 108.540 140.860 ;
        RECT 109.660 140.540 109.920 140.860 ;
        RECT 105.980 139.520 106.240 139.840 ;
        RECT 107.820 139.520 108.080 139.840 ;
        RECT 105.520 138.840 105.780 139.160 ;
        RECT 106.440 137.820 106.700 138.140 ;
        RECT 104.140 133.400 104.400 133.720 ;
        RECT 104.600 133.400 104.860 133.720 ;
        RECT 104.200 131.000 104.340 133.400 ;
        RECT 104.660 131.340 104.800 133.400 ;
        RECT 106.500 133.040 106.640 137.820 ;
        RECT 108.340 136.780 108.480 140.540 ;
        RECT 110.120 138.500 110.380 138.820 ;
        RECT 108.280 136.460 108.540 136.780 ;
        RECT 106.900 135.440 107.160 135.760 ;
        RECT 106.960 133.720 107.100 135.440 ;
        RECT 108.340 133.720 108.480 136.460 ;
        RECT 110.180 135.420 110.320 138.500 ;
        RECT 111.560 135.760 111.700 141.220 ;
        RECT 113.800 140.540 114.060 140.860 ;
        RECT 113.860 139.840 114.000 140.540 ;
        RECT 114.880 140.005 116.420 140.375 ;
        RECT 116.620 139.840 116.760 144.280 ;
        RECT 113.800 139.520 114.060 139.840 ;
        RECT 116.560 139.520 116.820 139.840 ;
        RECT 118.000 138.820 118.140 146.660 ;
        RECT 118.920 141.280 119.060 152.440 ;
        RECT 119.380 146.980 119.520 165.020 ;
        RECT 120.760 150.380 120.900 173.860 ;
        RECT 122.540 173.180 122.800 173.500 ;
        RECT 122.600 168.740 122.740 173.180 ;
        RECT 123.520 172.480 123.660 176.920 ;
        RECT 123.460 172.160 123.720 172.480 ;
        RECT 124.380 171.480 124.640 171.800 ;
        RECT 123.000 171.140 123.260 171.460 ;
        RECT 121.160 168.420 121.420 168.740 ;
        RECT 122.540 168.420 122.800 168.740 ;
        RECT 121.220 165.340 121.360 168.420 ;
        RECT 121.160 165.020 121.420 165.340 ;
        RECT 123.060 152.760 123.200 171.140 ;
        RECT 124.440 169.760 124.580 171.480 ;
        RECT 124.380 169.440 124.640 169.760 ;
        RECT 124.900 166.700 125.040 185.080 ;
        RECT 125.360 182.760 125.500 190.180 ;
        RECT 125.760 184.740 126.020 185.060 ;
        RECT 125.820 184.120 125.960 184.740 ;
        RECT 125.820 183.980 126.420 184.120 ;
        RECT 126.680 184.060 126.940 184.380 ;
        RECT 125.750 182.760 126.030 182.875 ;
        RECT 125.360 182.620 126.030 182.760 ;
        RECT 125.750 182.505 126.030 182.620 ;
        RECT 125.760 182.360 126.020 182.505 ;
        RECT 125.300 175.900 125.560 176.220 ;
        RECT 125.360 175.200 125.500 175.900 ;
        RECT 125.300 174.880 125.560 175.200 ;
        RECT 125.820 174.180 125.960 182.360 ;
        RECT 126.280 182.000 126.420 183.980 ;
        RECT 126.740 183.360 126.880 184.060 ;
        RECT 126.680 183.040 126.940 183.360 ;
        RECT 126.220 181.680 126.480 182.000 ;
        RECT 125.760 173.860 126.020 174.180 ;
        RECT 124.840 166.380 125.100 166.700 ;
        RECT 124.900 158.540 125.040 166.380 ;
        RECT 127.200 166.360 127.340 206.160 ;
        RECT 129.440 205.820 129.700 206.140 ;
        RECT 127.600 201.060 127.860 201.380 ;
        RECT 127.660 199.340 127.800 201.060 ;
        RECT 127.600 199.020 127.860 199.340 ;
        RECT 127.660 193.220 127.800 199.020 ;
        RECT 129.500 199.000 129.640 205.820 ;
        RECT 132.305 202.565 133.845 202.935 ;
        RECT 129.440 198.680 129.700 199.000 ;
        RECT 132.305 197.125 133.845 197.495 ;
        RECT 130.820 193.240 131.080 193.560 ;
        RECT 127.600 192.900 127.860 193.220 ;
        RECT 127.660 185.400 127.800 192.900 ;
        RECT 129.440 192.220 129.700 192.540 ;
        RECT 129.500 191.520 129.640 192.220 ;
        RECT 130.880 191.520 131.020 193.240 ;
        RECT 131.280 192.220 131.540 192.540 ;
        RECT 129.440 191.200 129.700 191.520 ;
        RECT 130.820 191.200 131.080 191.520 ;
        RECT 131.340 190.500 131.480 192.220 ;
        RECT 132.305 191.685 133.845 192.055 ;
        RECT 130.360 190.180 130.620 190.500 ;
        RECT 131.280 190.180 131.540 190.500 ;
        RECT 127.600 185.080 127.860 185.400 ;
        RECT 129.900 184.400 130.160 184.720 ;
        RECT 129.960 183.360 130.100 184.400 ;
        RECT 129.900 183.040 130.160 183.360 ;
        RECT 129.900 179.640 130.160 179.960 ;
        RECT 127.600 178.620 127.860 178.940 ;
        RECT 127.660 177.920 127.800 178.620 ;
        RECT 127.600 177.600 127.860 177.920 ;
        RECT 129.960 172.480 130.100 179.640 ;
        RECT 130.420 176.560 130.560 190.180 ;
        RECT 132.305 186.245 133.845 186.615 ;
        RECT 134.500 184.060 134.760 184.380 ;
        RECT 132.305 180.805 133.845 181.175 ;
        RECT 134.560 179.620 134.700 184.060 ;
        RECT 134.500 179.300 134.760 179.620 ;
        RECT 130.360 176.240 130.620 176.560 ;
        RECT 132.305 175.365 133.845 175.735 ;
        RECT 129.900 172.160 130.160 172.480 ;
        RECT 132.305 169.925 133.845 170.295 ;
        RECT 146.520 168.595 146.660 215.190 ;
        RECT 149.725 210.725 151.265 211.095 ;
        RECT 149.725 205.285 151.265 205.655 ;
        RECT 149.725 199.845 151.265 200.215 ;
        RECT 149.725 194.405 151.265 194.775 ;
        RECT 149.725 188.965 151.265 189.335 ;
        RECT 149.725 183.525 151.265 183.895 ;
        RECT 149.725 178.085 151.265 178.455 ;
        RECT 149.725 172.645 151.265 173.015 ;
        RECT 146.450 168.225 146.730 168.595 ;
        RECT 149.725 167.205 151.265 167.575 ;
        RECT 127.140 166.040 127.400 166.360 ;
        RECT 132.305 164.485 133.845 164.855 ;
        RECT 149.725 161.765 151.265 162.135 ;
        RECT 132.305 159.045 133.845 159.415 ;
        RECT 124.840 158.220 125.100 158.540 ;
        RECT 149.725 156.325 151.265 156.695 ;
        RECT 132.305 153.605 133.845 153.975 ;
        RECT 123.000 152.440 123.260 152.760 ;
        RECT 120.700 150.060 120.960 150.380 ;
        RECT 123.060 150.040 123.200 152.440 ;
        RECT 149.725 150.885 151.265 151.255 ;
        RECT 123.000 149.720 123.260 150.040 ;
        RECT 132.305 148.165 133.845 148.535 ;
        RECT 119.320 146.660 119.580 146.980 ;
        RECT 149.725 145.445 151.265 145.815 ;
        RECT 119.780 143.260 120.040 143.580 ;
        RECT 118.460 141.200 119.060 141.280 ;
        RECT 119.840 141.200 119.980 143.260 ;
        RECT 132.305 142.725 133.845 143.095 ;
        RECT 118.400 141.140 119.060 141.200 ;
        RECT 118.400 140.880 118.660 141.140 ;
        RECT 119.780 140.880 120.040 141.200 ;
        RECT 117.940 138.500 118.200 138.820 ;
        RECT 111.500 135.440 111.760 135.760 ;
        RECT 110.120 135.100 110.380 135.420 ;
        RECT 110.180 133.720 110.320 135.100 ;
        RECT 114.880 134.565 116.420 134.935 ;
        RECT 106.900 133.400 107.160 133.720 ;
        RECT 108.280 133.400 108.540 133.720 ;
        RECT 110.120 133.400 110.380 133.720 ;
        RECT 106.440 132.720 106.700 133.040 ;
        RECT 112.880 132.380 113.140 132.700 ;
        RECT 104.600 131.020 104.860 131.340 ;
        RECT 104.140 130.680 104.400 131.000 ;
        RECT 112.940 130.660 113.080 132.380 ;
        RECT 118.460 131.680 118.600 140.880 ;
        RECT 149.725 140.005 151.265 140.375 ;
        RECT 132.305 137.285 133.845 137.655 ;
        RECT 149.725 134.565 151.265 134.935 ;
        RECT 132.305 131.845 133.845 132.215 ;
        RECT 118.400 131.360 118.660 131.680 ;
        RECT 102.300 130.340 102.560 130.660 ;
        RECT 112.880 130.340 113.140 130.660 ;
        RECT 114.880 129.125 116.420 129.495 ;
        RECT 149.725 129.125 151.265 129.495 ;
        RECT 99.080 127.960 99.340 128.280 ;
        RECT 97.460 126.405 99.000 126.775 ;
        RECT 132.305 126.405 133.845 126.775 ;
        RECT 64.580 124.900 64.840 125.220 ;
        RECT 96.320 124.900 96.580 125.220 ;
        RECT 59.060 124.560 59.320 124.880 ;
        RECT 80.035 123.685 81.575 124.055 ;
        RECT 114.880 123.685 116.420 124.055 ;
        RECT 149.725 123.685 151.265 124.055 ;
        RECT 54.460 123.200 54.720 123.520 ;
        RECT 49.400 122.860 49.660 123.180 ;
        RECT 47.560 122.520 47.820 122.840 ;
        RECT 27.770 120.965 29.310 121.335 ;
        RECT 62.615 120.965 64.155 121.335 ;
        RECT 97.460 120.965 99.000 121.335 ;
        RECT 132.305 120.965 133.845 121.335 ;
        RECT 45.190 118.245 46.730 118.615 ;
        RECT 80.035 118.245 81.575 118.615 ;
        RECT 114.880 118.245 116.420 118.615 ;
        RECT 149.725 118.245 151.265 118.615 ;
        RECT 27.770 115.525 29.310 115.895 ;
        RECT 62.615 115.525 64.155 115.895 ;
        RECT 97.460 115.525 99.000 115.895 ;
        RECT 132.305 115.525 133.845 115.895 ;
        RECT 45.190 112.805 46.730 113.175 ;
        RECT 80.035 112.805 81.575 113.175 ;
        RECT 114.880 112.805 116.420 113.175 ;
        RECT 149.725 112.805 151.265 113.175 ;
        RECT 27.770 110.085 29.310 110.455 ;
        RECT 62.615 110.085 64.155 110.455 ;
        RECT 97.460 110.085 99.000 110.455 ;
        RECT 132.305 110.085 133.845 110.455 ;
        RECT 45.190 107.365 46.730 107.735 ;
        RECT 80.035 107.365 81.575 107.735 ;
        RECT 114.880 107.365 116.420 107.735 ;
        RECT 149.725 107.365 151.265 107.735 ;
        RECT 27.770 104.645 29.310 105.015 ;
        RECT 62.615 104.645 64.155 105.015 ;
        RECT 97.460 104.645 99.000 105.015 ;
        RECT 132.305 104.645 133.845 105.015 ;
        RECT 45.190 101.925 46.730 102.295 ;
        RECT 80.035 101.925 81.575 102.295 ;
        RECT 114.880 101.925 116.420 102.295 ;
        RECT 149.725 101.925 151.265 102.295 ;
        RECT 27.770 99.205 29.310 99.575 ;
        RECT 62.615 99.205 64.155 99.575 ;
        RECT 97.460 99.205 99.000 99.575 ;
        RECT 132.305 99.205 133.845 99.575 ;
        RECT 45.190 96.485 46.730 96.855 ;
        RECT 80.035 96.485 81.575 96.855 ;
        RECT 114.880 96.485 116.420 96.855 ;
        RECT 149.725 96.485 151.265 96.855 ;
        RECT 27.770 93.765 29.310 94.135 ;
        RECT 62.615 93.765 64.155 94.135 ;
        RECT 97.460 93.765 99.000 94.135 ;
        RECT 132.305 93.765 133.845 94.135 ;
        RECT 45.190 91.045 46.730 91.415 ;
        RECT 80.035 91.045 81.575 91.415 ;
        RECT 114.880 91.045 116.420 91.415 ;
        RECT 149.725 91.045 151.265 91.415 ;
        RECT 27.770 88.325 29.310 88.695 ;
        RECT 62.615 88.325 64.155 88.695 ;
        RECT 97.460 88.325 99.000 88.695 ;
        RECT 132.305 88.325 133.845 88.695 ;
        RECT 45.190 85.605 46.730 85.975 ;
        RECT 80.035 85.605 81.575 85.975 ;
        RECT 114.880 85.605 116.420 85.975 ;
        RECT 149.725 85.605 151.265 85.975 ;
        RECT 27.770 82.885 29.310 83.255 ;
        RECT 62.615 82.885 64.155 83.255 ;
        RECT 97.460 82.885 99.000 83.255 ;
        RECT 132.305 82.885 133.845 83.255 ;
        RECT 45.190 80.165 46.730 80.535 ;
        RECT 80.035 80.165 81.575 80.535 ;
        RECT 114.880 80.165 116.420 80.535 ;
        RECT 149.725 80.165 151.265 80.535 ;
        RECT 27.770 77.445 29.310 77.815 ;
        RECT 62.615 77.445 64.155 77.815 ;
        RECT 97.460 77.445 99.000 77.815 ;
        RECT 132.305 77.445 133.845 77.815 ;
        RECT 45.190 74.725 46.730 75.095 ;
        RECT 80.035 74.725 81.575 75.095 ;
        RECT 114.880 74.725 116.420 75.095 ;
        RECT 149.725 74.725 151.265 75.095 ;
        RECT 54.930 54.700 77.070 59.620 ;
        RECT 62.000 49.240 62.940 49.700 ;
        RECT 64.680 49.250 65.590 49.750 ;
        RECT 78.760 49.110 79.750 49.690 ;
        RECT 81.010 48.920 82.950 51.960 ;
        RECT 95.020 50.660 105.690 60.270 ;
        RECT 117.160 54.670 134.820 58.500 ;
        RECT 78.760 48.340 82.950 48.920 ;
        RECT 124.230 48.840 125.170 49.300 ;
        RECT 126.910 48.850 127.820 49.350 ;
        RECT 140.990 48.710 141.980 49.290 ;
        RECT 143.240 48.520 145.180 51.560 ;
        RECT 78.760 48.330 79.750 48.340 ;
        RECT 78.750 47.530 79.740 48.110 ;
        RECT 81.010 47.510 82.950 48.340 ;
        RECT 140.990 47.940 145.180 48.520 ;
        RECT 140.990 47.930 141.980 47.940 ;
        RECT 64.630 47.305 65.640 47.330 ;
        RECT 77.540 47.305 78.230 47.360 ;
        RECT 81.030 47.330 82.050 47.510 ;
        RECT 64.630 46.875 78.505 47.305 ;
        RECT 64.630 46.860 65.640 46.875 ;
        RECT 62.000 44.600 62.940 45.060 ;
        RECT 64.680 44.580 65.590 45.080 ;
        RECT 64.630 42.735 65.640 42.770 ;
        RECT 66.425 42.735 66.855 46.875 ;
        RECT 77.540 46.820 78.230 46.875 ;
        RECT 78.750 46.750 82.050 47.330 ;
        RECT 140.980 47.130 141.970 47.710 ;
        RECT 143.240 47.110 145.180 47.940 ;
        RECT 78.740 45.960 79.730 46.540 ;
        RECT 81.030 45.740 82.050 46.750 ;
        RECT 126.860 46.905 127.870 46.930 ;
        RECT 139.770 46.905 140.460 46.960 ;
        RECT 143.260 46.930 144.280 47.110 ;
        RECT 126.860 46.475 140.735 46.905 ;
        RECT 126.860 46.460 127.870 46.475 ;
        RECT 78.750 45.160 82.050 45.740 ;
        RECT 78.770 44.370 79.760 44.950 ;
        RECT 81.030 44.170 82.050 45.160 ;
        RECT 124.230 44.200 125.170 44.660 ;
        RECT 126.910 44.180 127.820 44.680 ;
        RECT 78.760 43.590 82.050 44.170 ;
        RECT 78.770 42.790 79.760 43.370 ;
        RECT 64.630 42.305 66.855 42.735 ;
        RECT 81.030 42.590 82.050 43.590 ;
        RECT 75.030 42.570 75.890 42.580 ;
        RECT 73.620 42.450 75.890 42.570 ;
        RECT 64.630 42.300 65.640 42.305 ;
        RECT 62.010 40.030 62.950 40.490 ;
        RECT 64.670 40.010 65.580 40.510 ;
        RECT 64.630 38.145 65.640 38.190 ;
        RECT 66.425 38.145 66.855 42.305 ;
        RECT 73.610 41.990 75.890 42.450 ;
        RECT 78.760 42.030 82.050 42.590 ;
        RECT 78.760 42.010 79.750 42.030 ;
        RECT 73.620 41.840 75.890 41.990 ;
        RECT 73.590 39.770 74.540 40.150 ;
        RECT 64.615 37.715 66.855 38.145 ;
        RECT 75.030 38.020 75.890 41.840 ;
        RECT 78.770 41.210 79.760 41.790 ;
        RECT 78.760 40.995 79.750 41.010 ;
        RECT 81.030 40.995 82.050 42.030 ;
        RECT 106.955 41.740 108.745 43.470 ;
        RECT 126.860 42.335 127.870 42.370 ;
        RECT 128.655 42.335 129.085 46.475 ;
        RECT 139.770 46.420 140.460 46.475 ;
        RECT 140.980 46.350 144.280 46.930 ;
        RECT 140.970 45.560 141.960 46.140 ;
        RECT 143.260 45.340 144.280 46.350 ;
        RECT 140.980 44.760 144.280 45.340 ;
        RECT 141.000 43.970 141.990 44.550 ;
        RECT 143.260 43.770 144.280 44.760 ;
        RECT 140.990 43.190 144.280 43.770 ;
        RECT 141.000 42.390 141.990 42.970 ;
        RECT 126.860 41.905 129.085 42.335 ;
        RECT 143.260 42.190 144.280 43.190 ;
        RECT 137.260 42.170 138.120 42.180 ;
        RECT 135.850 42.050 138.120 42.170 ;
        RECT 126.860 41.900 127.870 41.905 ;
        RECT 78.760 40.435 82.050 40.995 ;
        RECT 78.760 40.430 79.750 40.435 ;
        RECT 78.750 39.630 79.740 40.210 ;
        RECT 78.760 39.425 79.750 39.430 ;
        RECT 81.030 39.425 82.050 40.435 ;
        RECT 78.760 38.870 82.050 39.425 ;
        RECT 78.760 38.850 79.750 38.870 ;
        RECT 78.760 38.050 79.750 38.630 ;
        RECT 62.030 35.490 62.940 35.890 ;
        RECT 64.690 35.440 65.590 35.890 ;
        RECT 64.760 35.110 65.790 35.160 ;
        RECT 66.425 35.110 66.855 37.715 ;
        RECT 73.600 37.290 75.890 38.020 ;
        RECT 64.750 34.680 66.855 35.110 ;
        RECT 73.580 35.060 74.540 35.670 ;
        RECT 64.760 34.640 65.790 34.680 ;
        RECT 75.030 33.490 75.890 37.290 ;
        RECT 78.760 37.825 79.750 37.840 ;
        RECT 81.030 37.825 82.050 38.870 ;
        RECT 95.110 38.060 96.110 39.160 ;
        RECT 78.760 37.270 82.050 37.825 ;
        RECT 78.760 37.260 79.750 37.270 ;
        RECT 78.770 36.470 79.760 37.050 ;
        RECT 81.030 36.260 82.050 37.270 ;
        RECT 95.360 36.700 95.900 38.060 ;
        RECT 97.400 38.040 98.400 39.140 ;
        RECT 99.690 38.020 100.690 39.120 ;
        RECT 101.950 38.040 102.950 39.140 ;
        RECT 104.240 38.040 105.240 39.140 ;
        RECT 99.920 36.700 100.460 38.020 ;
        RECT 104.470 36.700 105.010 38.040 ;
        RECT 78.760 35.680 82.050 36.260 ;
        RECT 78.770 34.900 79.760 35.480 ;
        RECT 81.030 34.670 82.050 35.680 ;
        RECT 95.330 35.460 105.150 36.700 ;
        RECT 78.760 34.110 82.050 34.670 ;
        RECT 78.760 34.090 81.690 34.110 ;
        RECT 78.760 33.810 79.700 33.850 ;
        RECT 78.760 33.770 79.720 33.810 ;
        RECT 59.530 30.960 64.390 33.110 ;
        RECT 73.530 32.760 75.890 33.490 ;
        RECT 78.730 33.250 79.750 33.770 ;
        RECT 75.030 31.850 75.890 32.760 ;
        RECT 78.750 31.850 79.750 33.250 ;
        RECT 75.030 31.550 84.770 31.850 ;
        RECT 54.960 30.310 55.960 30.420 ;
        RECT 51.990 29.440 55.960 30.310 ;
        RECT 51.990 21.815 52.860 29.440 ;
        RECT 54.960 28.510 55.960 29.440 ;
        RECT 59.530 28.760 60.875 30.960 ;
        RECT 63.420 30.950 64.390 30.960 ;
        RECT 73.580 30.520 74.540 31.040 ;
        RECT 75.030 30.950 90.920 31.550 ;
        RECT 75.030 30.590 84.770 30.950 ;
        RECT 66.585 30.215 67.240 30.230 ;
        RECT 66.585 29.645 69.925 30.215 ;
        RECT 66.585 29.635 67.240 29.645 ;
        RECT 64.260 29.300 65.290 29.340 ;
        RECT 66.200 29.300 67.280 29.340 ;
        RECT 64.260 28.820 67.280 29.300 ;
        RECT 59.530 28.590 60.870 28.760 ;
        RECT 57.840 27.790 62.690 28.590 ;
        RECT 66.760 27.870 67.280 28.820 ;
        RECT 69.355 28.090 69.925 29.645 ;
        RECT 75.030 28.850 75.890 30.590 ;
        RECT 73.560 28.120 75.890 28.850 ;
        RECT 55.540 25.000 55.800 26.520 ;
        RECT 57.840 25.420 58.120 27.790 ;
        RECT 60.120 25.420 60.400 26.520 ;
        RECT 62.410 25.420 62.690 27.790 ;
        RECT 64.710 25.420 64.990 26.520 ;
        RECT 60.130 25.000 60.390 25.420 ;
        RECT 64.720 25.000 64.980 25.420 ;
        RECT 55.540 23.840 64.980 25.000 ;
        RECT 55.560 23.790 64.950 23.840 ;
        RECT 66.520 22.580 67.520 27.870 ;
        RECT 69.140 23.520 70.140 28.090 ;
        RECT 73.590 26.000 74.540 26.440 ;
        RECT 90.320 23.705 90.920 30.950 ;
        RECT 106.985 29.840 108.715 41.740 ;
        RECT 124.240 39.630 125.180 40.090 ;
        RECT 126.900 39.610 127.810 40.110 ;
        RECT 126.860 37.745 127.870 37.790 ;
        RECT 128.655 37.745 129.085 41.905 ;
        RECT 135.840 41.590 138.120 42.050 ;
        RECT 140.990 41.630 144.280 42.190 ;
        RECT 140.990 41.610 141.980 41.630 ;
        RECT 135.850 41.440 138.120 41.590 ;
        RECT 135.820 39.370 136.770 39.750 ;
        RECT 126.845 37.315 129.085 37.745 ;
        RECT 137.260 37.620 138.120 41.440 ;
        RECT 141.000 40.810 141.990 41.390 ;
        RECT 140.990 40.595 141.980 40.610 ;
        RECT 143.260 40.595 144.280 41.630 ;
        RECT 140.990 40.035 144.280 40.595 ;
        RECT 140.990 40.030 141.980 40.035 ;
        RECT 140.980 39.230 141.970 39.810 ;
        RECT 140.990 39.025 141.980 39.030 ;
        RECT 143.260 39.025 144.280 40.035 ;
        RECT 140.990 38.470 144.280 39.025 ;
        RECT 140.990 38.450 141.980 38.470 ;
        RECT 140.990 37.650 141.980 38.230 ;
        RECT 124.260 35.090 125.170 35.490 ;
        RECT 126.920 35.040 127.820 35.490 ;
        RECT 126.990 34.710 128.020 34.760 ;
        RECT 128.655 34.710 129.085 37.315 ;
        RECT 135.830 36.890 138.120 37.620 ;
        RECT 126.980 34.280 129.085 34.710 ;
        RECT 135.810 34.660 136.770 35.270 ;
        RECT 126.990 34.240 128.020 34.280 ;
        RECT 137.260 33.090 138.120 36.890 ;
        RECT 140.990 37.425 141.980 37.440 ;
        RECT 143.260 37.425 144.280 38.470 ;
        RECT 140.990 36.870 144.280 37.425 ;
        RECT 140.990 36.860 141.980 36.870 ;
        RECT 141.000 36.070 141.990 36.650 ;
        RECT 143.260 35.860 144.280 36.870 ;
        RECT 140.990 35.280 144.280 35.860 ;
        RECT 141.000 34.500 141.990 35.080 ;
        RECT 143.260 34.270 144.280 35.280 ;
        RECT 140.990 33.710 144.280 34.270 ;
        RECT 140.990 33.690 143.920 33.710 ;
        RECT 140.990 33.410 141.930 33.450 ;
        RECT 140.990 33.370 141.950 33.410 ;
        RECT 121.760 30.560 126.620 32.710 ;
        RECT 135.760 32.360 138.120 33.090 ;
        RECT 140.960 32.850 141.980 33.370 ;
        RECT 137.260 31.450 138.120 32.360 ;
        RECT 140.980 31.450 141.980 32.850 ;
        RECT 137.260 31.150 147.000 31.450 ;
        RECT 106.985 29.830 113.910 29.840 ;
        RECT 117.190 29.830 118.190 30.020 ;
        RECT 106.985 29.070 118.190 29.830 ;
        RECT 106.985 29.050 111.750 29.070 ;
        RECT 107.225 26.410 108.095 29.050 ;
        RECT 117.190 28.110 118.190 29.070 ;
        RECT 121.760 28.360 123.105 30.560 ;
        RECT 125.650 30.550 126.620 30.560 ;
        RECT 135.810 30.120 136.770 30.640 ;
        RECT 137.260 30.550 151.130 31.150 ;
        RECT 137.260 30.190 147.000 30.550 ;
        RECT 128.815 29.815 129.470 29.830 ;
        RECT 128.815 29.245 132.155 29.815 ;
        RECT 128.815 29.235 129.470 29.245 ;
        RECT 126.490 28.900 127.520 28.940 ;
        RECT 128.430 28.900 129.510 28.940 ;
        RECT 126.490 28.420 129.510 28.900 ;
        RECT 121.760 28.190 123.100 28.360 ;
        RECT 120.070 27.390 124.920 28.190 ;
        RECT 128.990 27.470 129.510 28.420 ;
        RECT 131.585 27.690 132.155 29.245 ;
        RECT 137.260 28.450 138.120 30.190 ;
        RECT 135.790 27.720 138.120 28.450 ;
        RECT 107.205 25.590 108.115 26.410 ;
        RECT 107.225 25.565 108.095 25.590 ;
        RECT 117.770 24.600 118.030 26.120 ;
        RECT 120.070 25.020 120.350 27.390 ;
        RECT 122.350 25.020 122.630 26.120 ;
        RECT 124.640 25.020 124.920 27.390 ;
        RECT 126.940 25.020 127.220 26.120 ;
        RECT 122.360 24.600 122.620 25.020 ;
        RECT 126.950 24.600 127.210 25.020 ;
        RECT 69.130 23.320 70.140 23.520 ;
        RECT 69.030 22.720 70.140 23.320 ;
        RECT 90.300 23.155 90.940 23.705 ;
        RECT 117.770 23.440 127.210 24.600 ;
        RECT 117.790 23.390 127.180 23.440 ;
        RECT 90.320 23.130 90.920 23.155 ;
        RECT 51.990 20.945 60.930 21.815 ;
        RECT 55.150 10.850 64.860 18.920 ;
        RECT 66.730 9.340 67.330 22.580 ;
        RECT 69.130 22.520 70.140 22.720 ;
        RECT 61.300 8.740 67.330 9.340 ;
        RECT 56.435 5.380 56.985 5.400 ;
        RECT 61.300 5.380 61.900 8.740 ;
        RECT 69.450 7.975 70.050 22.520 ;
        RECT 128.750 22.180 129.750 27.470 ;
        RECT 131.370 23.120 132.370 27.690 ;
        RECT 135.820 25.600 136.770 26.040 ;
        RECT 73.660 10.790 84.410 18.850 ;
        RECT 94.350 11.450 105.980 18.660 ;
        RECT 117.190 13.030 127.820 18.860 ;
        RECT 69.430 7.425 70.070 7.975 ;
        RECT 69.450 7.400 70.050 7.425 ;
        RECT 128.970 7.165 129.570 22.180 ;
        RECT 131.360 22.120 132.370 23.120 ;
        RECT 131.570 20.610 132.170 22.120 ;
        RECT 150.530 20.735 151.130 30.550 ;
        RECT 134.505 20.610 135.055 20.630 ;
        RECT 131.570 20.010 135.080 20.610 ;
        RECT 150.510 20.185 151.150 20.735 ;
        RECT 150.530 20.160 151.130 20.185 ;
        RECT 134.505 19.990 135.055 20.010 ;
        RECT 135.840 13.390 146.360 18.670 ;
        RECT 128.950 6.615 129.590 7.165 ;
        RECT 128.970 6.590 129.570 6.615 ;
        RECT 56.410 4.780 61.900 5.380 ;
        RECT 56.435 4.760 56.985 4.780 ;
      LAYER via2 ;
        RECT 57.790 223.420 58.090 223.720 ;
        RECT 35.120 216.570 35.420 216.870 ;
        RECT 25.000 216.150 25.300 216.450 ;
        RECT 73.880 220.580 74.180 220.880 ;
        RECT 85.720 218.450 86.020 218.750 ;
        RECT 55.360 217.100 55.660 217.400 ;
        RECT 45.240 215.750 45.540 216.050 ;
        RECT 69.160 216.900 69.460 217.200 ;
        RECT 79.580 217.740 79.880 218.040 ;
        RECT 126.950 223.590 127.250 223.890 ;
        RECT 105.960 217.840 106.260 218.140 ;
        RECT 143.810 221.120 144.110 221.420 ;
        RECT 151.190 220.060 151.490 220.360 ;
        RECT 126.200 218.210 126.500 218.510 ;
        RECT 146.440 217.400 146.740 217.700 ;
        RECT 27.800 213.490 28.080 213.770 ;
        RECT 28.200 213.490 28.480 213.770 ;
        RECT 28.600 213.490 28.880 213.770 ;
        RECT 29.000 213.490 29.280 213.770 ;
        RECT 27.800 208.050 28.080 208.330 ;
        RECT 28.200 208.050 28.480 208.330 ;
        RECT 28.600 208.050 28.880 208.330 ;
        RECT 29.000 208.050 29.280 208.330 ;
        RECT 27.800 202.610 28.080 202.890 ;
        RECT 28.200 202.610 28.480 202.890 ;
        RECT 28.600 202.610 28.880 202.890 ;
        RECT 29.000 202.610 29.280 202.890 ;
        RECT 27.800 197.170 28.080 197.450 ;
        RECT 28.200 197.170 28.480 197.450 ;
        RECT 28.600 197.170 28.880 197.450 ;
        RECT 29.000 197.170 29.280 197.450 ;
        RECT 19.490 187.310 19.770 187.590 ;
        RECT 27.800 191.730 28.080 192.010 ;
        RECT 28.200 191.730 28.480 192.010 ;
        RECT 28.600 191.730 28.880 192.010 ;
        RECT 29.000 191.730 29.280 192.010 ;
        RECT 27.800 186.290 28.080 186.570 ;
        RECT 28.200 186.290 28.480 186.570 ;
        RECT 28.600 186.290 28.880 186.570 ;
        RECT 29.000 186.290 29.280 186.570 ;
        RECT 30.070 184.590 30.350 184.870 ;
        RECT 27.800 180.850 28.080 181.130 ;
        RECT 28.200 180.850 28.480 181.130 ;
        RECT 28.600 180.850 28.880 181.130 ;
        RECT 29.000 180.850 29.280 181.130 ;
        RECT 27.800 175.410 28.080 175.690 ;
        RECT 28.200 175.410 28.480 175.690 ;
        RECT 28.600 175.410 28.880 175.690 ;
        RECT 29.000 175.410 29.280 175.690 ;
        RECT 26.390 168.950 26.670 169.230 ;
        RECT 27.800 169.970 28.080 170.250 ;
        RECT 28.200 169.970 28.480 170.250 ;
        RECT 28.600 169.970 28.880 170.250 ;
        RECT 29.000 169.970 29.280 170.250 ;
        RECT 27.800 164.530 28.080 164.810 ;
        RECT 28.200 164.530 28.480 164.810 ;
        RECT 28.600 164.530 28.880 164.810 ;
        RECT 29.000 164.530 29.280 164.810 ;
        RECT 27.800 159.090 28.080 159.370 ;
        RECT 28.200 159.090 28.480 159.370 ;
        RECT 28.600 159.090 28.880 159.370 ;
        RECT 29.000 159.090 29.280 159.370 ;
        RECT 27.800 153.650 28.080 153.930 ;
        RECT 28.200 153.650 28.480 153.930 ;
        RECT 28.600 153.650 28.880 153.930 ;
        RECT 29.000 153.650 29.280 153.930 ;
        RECT 27.800 148.210 28.080 148.490 ;
        RECT 28.200 148.210 28.480 148.490 ;
        RECT 28.600 148.210 28.880 148.490 ;
        RECT 29.000 148.210 29.280 148.490 ;
        RECT 27.800 142.770 28.080 143.050 ;
        RECT 28.200 142.770 28.480 143.050 ;
        RECT 28.600 142.770 28.880 143.050 ;
        RECT 29.000 142.770 29.280 143.050 ;
        RECT 27.800 137.330 28.080 137.610 ;
        RECT 28.200 137.330 28.480 137.610 ;
        RECT 28.600 137.330 28.880 137.610 ;
        RECT 29.000 137.330 29.280 137.610 ;
        RECT 35.130 184.590 35.410 184.870 ;
        RECT 36.970 174.390 37.250 174.670 ;
        RECT 39.270 168.950 39.550 169.230 ;
        RECT 45.220 210.770 45.500 211.050 ;
        RECT 45.620 210.770 45.900 211.050 ;
        RECT 46.020 210.770 46.300 211.050 ;
        RECT 46.420 210.770 46.700 211.050 ;
        RECT 45.220 205.330 45.500 205.610 ;
        RECT 45.620 205.330 45.900 205.610 ;
        RECT 46.020 205.330 46.300 205.610 ;
        RECT 46.420 205.330 46.700 205.610 ;
        RECT 45.220 199.890 45.500 200.170 ;
        RECT 45.620 199.890 45.900 200.170 ;
        RECT 46.020 199.890 46.300 200.170 ;
        RECT 46.420 199.890 46.700 200.170 ;
        RECT 45.220 194.450 45.500 194.730 ;
        RECT 45.620 194.450 45.900 194.730 ;
        RECT 46.020 194.450 46.300 194.730 ;
        RECT 46.420 194.450 46.700 194.730 ;
        RECT 45.220 189.010 45.500 189.290 ;
        RECT 45.620 189.010 45.900 189.290 ;
        RECT 46.020 189.010 46.300 189.290 ;
        RECT 46.420 189.010 46.700 189.290 ;
        RECT 45.220 183.570 45.500 183.850 ;
        RECT 45.620 183.570 45.900 183.850 ;
        RECT 46.020 183.570 46.300 183.850 ;
        RECT 46.420 183.570 46.700 183.850 ;
        RECT 47.090 181.870 47.370 182.150 ;
        RECT 45.220 178.130 45.500 178.410 ;
        RECT 45.620 178.130 45.900 178.410 ;
        RECT 46.020 178.130 46.300 178.410 ;
        RECT 46.420 178.130 46.700 178.410 ;
        RECT 45.220 172.690 45.500 172.970 ;
        RECT 45.620 172.690 45.900 172.970 ;
        RECT 46.020 172.690 46.300 172.970 ;
        RECT 46.420 172.690 46.700 172.970 ;
        RECT 62.645 213.490 62.925 213.770 ;
        RECT 63.045 213.490 63.325 213.770 ;
        RECT 63.445 213.490 63.725 213.770 ;
        RECT 63.845 213.490 64.125 213.770 ;
        RECT 45.220 167.250 45.500 167.530 ;
        RECT 45.620 167.250 45.900 167.530 ;
        RECT 46.020 167.250 46.300 167.530 ;
        RECT 46.420 167.250 46.700 167.530 ;
        RECT 45.220 161.810 45.500 162.090 ;
        RECT 45.620 161.810 45.900 162.090 ;
        RECT 46.020 161.810 46.300 162.090 ;
        RECT 46.420 161.810 46.700 162.090 ;
        RECT 45.220 156.370 45.500 156.650 ;
        RECT 45.620 156.370 45.900 156.650 ;
        RECT 46.020 156.370 46.300 156.650 ;
        RECT 46.420 156.370 46.700 156.650 ;
        RECT 45.220 150.930 45.500 151.210 ;
        RECT 45.620 150.930 45.900 151.210 ;
        RECT 46.020 150.930 46.300 151.210 ;
        RECT 46.420 150.930 46.700 151.210 ;
        RECT 27.800 131.890 28.080 132.170 ;
        RECT 28.200 131.890 28.480 132.170 ;
        RECT 28.600 131.890 28.880 132.170 ;
        RECT 29.000 131.890 29.280 132.170 ;
        RECT 45.220 145.490 45.500 145.770 ;
        RECT 45.620 145.490 45.900 145.770 ;
        RECT 46.020 145.490 46.300 145.770 ;
        RECT 46.420 145.490 46.700 145.770 ;
        RECT 45.220 140.050 45.500 140.330 ;
        RECT 45.620 140.050 45.900 140.330 ;
        RECT 46.020 140.050 46.300 140.330 ;
        RECT 46.420 140.050 46.700 140.330 ;
        RECT 45.220 134.610 45.500 134.890 ;
        RECT 45.620 134.610 45.900 134.890 ;
        RECT 46.020 134.610 46.300 134.890 ;
        RECT 46.420 134.610 46.700 134.890 ;
        RECT 27.800 126.450 28.080 126.730 ;
        RECT 28.200 126.450 28.480 126.730 ;
        RECT 28.600 126.450 28.880 126.730 ;
        RECT 29.000 126.450 29.280 126.730 ;
        RECT 62.645 208.050 62.925 208.330 ;
        RECT 63.045 208.050 63.325 208.330 ;
        RECT 63.445 208.050 63.725 208.330 ;
        RECT 63.845 208.050 64.125 208.330 ;
        RECT 62.645 202.610 62.925 202.890 ;
        RECT 63.045 202.610 63.325 202.890 ;
        RECT 63.445 202.610 63.725 202.890 ;
        RECT 63.845 202.610 64.125 202.890 ;
        RECT 62.645 197.170 62.925 197.450 ;
        RECT 63.045 197.170 63.325 197.450 ;
        RECT 63.445 197.170 63.725 197.450 ;
        RECT 63.845 197.170 64.125 197.450 ;
        RECT 62.645 191.730 62.925 192.010 ;
        RECT 63.045 191.730 63.325 192.010 ;
        RECT 63.445 191.730 63.725 192.010 ;
        RECT 63.845 191.730 64.125 192.010 ;
        RECT 57.670 176.430 57.950 176.710 ;
        RECT 45.220 129.170 45.500 129.450 ;
        RECT 45.620 129.170 45.900 129.450 ;
        RECT 46.020 129.170 46.300 129.450 ;
        RECT 46.420 129.170 46.700 129.450 ;
        RECT 62.645 186.290 62.925 186.570 ;
        RECT 63.045 186.290 63.325 186.570 ;
        RECT 63.445 186.290 63.725 186.570 ;
        RECT 63.845 186.290 64.125 186.570 ;
        RECT 80.065 210.770 80.345 211.050 ;
        RECT 80.465 210.770 80.745 211.050 ;
        RECT 80.865 210.770 81.145 211.050 ;
        RECT 81.265 210.770 81.545 211.050 ;
        RECT 97.490 213.490 97.770 213.770 ;
        RECT 97.890 213.490 98.170 213.770 ;
        RECT 98.290 213.490 98.570 213.770 ;
        RECT 98.690 213.490 98.970 213.770 ;
        RECT 132.335 213.490 132.615 213.770 ;
        RECT 132.735 213.490 133.015 213.770 ;
        RECT 133.135 213.490 133.415 213.770 ;
        RECT 133.535 213.490 133.815 213.770 ;
        RECT 62.645 180.850 62.925 181.130 ;
        RECT 63.045 180.850 63.325 181.130 ;
        RECT 63.445 180.850 63.725 181.130 ;
        RECT 63.845 180.850 64.125 181.130 ;
        RECT 62.645 175.410 62.925 175.690 ;
        RECT 63.045 175.410 63.325 175.690 ;
        RECT 63.445 175.410 63.725 175.690 ;
        RECT 63.845 175.410 64.125 175.690 ;
        RECT 63.650 174.390 63.930 174.670 ;
        RECT 66.410 179.150 66.690 179.430 ;
        RECT 62.645 169.970 62.925 170.250 ;
        RECT 63.045 169.970 63.325 170.250 ;
        RECT 63.445 169.970 63.725 170.250 ;
        RECT 63.845 169.970 64.125 170.250 ;
        RECT 62.645 164.530 62.925 164.810 ;
        RECT 63.045 164.530 63.325 164.810 ;
        RECT 63.445 164.530 63.725 164.810 ;
        RECT 63.845 164.530 64.125 164.810 ;
        RECT 62.645 159.090 62.925 159.370 ;
        RECT 63.045 159.090 63.325 159.370 ;
        RECT 63.445 159.090 63.725 159.370 ;
        RECT 63.845 159.090 64.125 159.370 ;
        RECT 62.645 153.650 62.925 153.930 ;
        RECT 63.045 153.650 63.325 153.930 ;
        RECT 63.445 153.650 63.725 153.930 ;
        RECT 63.845 153.650 64.125 153.930 ;
        RECT 67.790 179.150 68.070 179.430 ;
        RECT 70.090 186.630 70.370 186.910 ;
        RECT 80.065 205.330 80.345 205.610 ;
        RECT 80.465 205.330 80.745 205.610 ;
        RECT 80.865 205.330 81.145 205.610 ;
        RECT 81.265 205.330 81.545 205.610 ;
        RECT 80.065 199.890 80.345 200.170 ;
        RECT 80.465 199.890 80.745 200.170 ;
        RECT 80.865 199.890 81.145 200.170 ;
        RECT 81.265 199.890 81.545 200.170 ;
        RECT 76.990 198.870 77.270 199.150 ;
        RECT 97.490 208.050 97.770 208.330 ;
        RECT 97.890 208.050 98.170 208.330 ;
        RECT 98.290 208.050 98.570 208.330 ;
        RECT 98.690 208.050 98.970 208.330 ;
        RECT 80.065 194.450 80.345 194.730 ;
        RECT 80.465 194.450 80.745 194.730 ;
        RECT 80.865 194.450 81.145 194.730 ;
        RECT 81.265 194.450 81.545 194.730 ;
        RECT 74.230 187.310 74.510 187.590 ;
        RECT 76.990 187.310 77.270 187.590 ;
        RECT 80.065 189.010 80.345 189.290 ;
        RECT 80.465 189.010 80.745 189.290 ;
        RECT 80.865 189.010 81.145 189.290 ;
        RECT 81.265 189.010 81.545 189.290 ;
        RECT 76.990 181.870 77.270 182.150 ;
        RECT 62.645 148.210 62.925 148.490 ;
        RECT 63.045 148.210 63.325 148.490 ;
        RECT 63.445 148.210 63.725 148.490 ;
        RECT 63.845 148.210 64.125 148.490 ;
        RECT 59.970 146.510 60.250 146.790 ;
        RECT 62.645 142.770 62.925 143.050 ;
        RECT 63.045 142.770 63.325 143.050 ;
        RECT 63.445 142.770 63.725 143.050 ;
        RECT 63.845 142.770 64.125 143.050 ;
        RECT 66.870 146.510 67.150 146.790 ;
        RECT 62.645 137.330 62.925 137.610 ;
        RECT 63.045 137.330 63.325 137.610 ;
        RECT 63.445 137.330 63.725 137.610 ;
        RECT 63.845 137.330 64.125 137.610 ;
        RECT 45.220 123.730 45.500 124.010 ;
        RECT 45.620 123.730 45.900 124.010 ;
        RECT 46.020 123.730 46.300 124.010 ;
        RECT 46.420 123.730 46.700 124.010 ;
        RECT 62.645 131.890 62.925 132.170 ;
        RECT 63.045 131.890 63.325 132.170 ;
        RECT 63.445 131.890 63.725 132.170 ;
        RECT 63.845 131.890 64.125 132.170 ;
        RECT 62.645 126.450 62.925 126.730 ;
        RECT 63.045 126.450 63.325 126.730 ;
        RECT 63.445 126.450 63.725 126.730 ;
        RECT 63.845 126.450 64.125 126.730 ;
        RECT 73.310 157.390 73.590 157.670 ;
        RECT 80.065 183.570 80.345 183.850 ;
        RECT 80.465 183.570 80.745 183.850 ;
        RECT 80.865 183.570 81.145 183.850 ;
        RECT 81.265 183.570 81.545 183.850 ;
        RECT 80.065 178.130 80.345 178.410 ;
        RECT 80.465 178.130 80.745 178.410 ;
        RECT 80.865 178.130 81.145 178.410 ;
        RECT 81.265 178.130 81.545 178.410 ;
        RECT 78.830 175.750 79.110 176.030 ;
        RECT 80.065 172.690 80.345 172.970 ;
        RECT 80.465 172.690 80.745 172.970 ;
        RECT 80.865 172.690 81.145 172.970 ;
        RECT 81.265 172.690 81.545 172.970 ;
        RECT 75.150 160.110 75.430 160.390 ;
        RECT 80.065 167.250 80.345 167.530 ;
        RECT 80.465 167.250 80.745 167.530 ;
        RECT 80.865 167.250 81.145 167.530 ;
        RECT 81.265 167.250 81.545 167.530 ;
        RECT 75.610 153.990 75.890 154.270 ;
        RECT 80.065 161.810 80.345 162.090 ;
        RECT 80.465 161.810 80.745 162.090 ;
        RECT 80.865 161.810 81.145 162.090 ;
        RECT 81.265 161.810 81.545 162.090 ;
        RECT 83.430 187.990 83.710 188.270 ;
        RECT 114.910 210.770 115.190 211.050 ;
        RECT 115.310 210.770 115.590 211.050 ;
        RECT 115.710 210.770 115.990 211.050 ;
        RECT 116.110 210.770 116.390 211.050 ;
        RECT 87.570 186.630 87.850 186.910 ;
        RECT 81.590 160.110 81.870 160.390 ;
        RECT 97.490 202.610 97.770 202.890 ;
        RECT 97.890 202.610 98.170 202.890 ;
        RECT 98.290 202.610 98.570 202.890 ;
        RECT 98.690 202.610 98.970 202.890 ;
        RECT 80.065 156.370 80.345 156.650 ;
        RECT 80.465 156.370 80.745 156.650 ;
        RECT 80.865 156.370 81.145 156.650 ;
        RECT 81.265 156.370 81.545 156.650 ;
        RECT 80.065 150.930 80.345 151.210 ;
        RECT 80.465 150.930 80.745 151.210 ;
        RECT 80.865 150.930 81.145 151.210 ;
        RECT 81.265 150.930 81.545 151.210 ;
        RECT 75.610 136.310 75.890 136.590 ;
        RECT 77.910 135.630 78.190 135.910 ;
        RECT 80.065 145.490 80.345 145.770 ;
        RECT 80.465 145.490 80.745 145.770 ;
        RECT 80.865 145.490 81.145 145.770 ;
        RECT 81.265 145.490 81.545 145.770 ;
        RECT 80.065 140.050 80.345 140.330 ;
        RECT 80.465 140.050 80.745 140.330 ;
        RECT 80.865 140.050 81.145 140.330 ;
        RECT 81.265 140.050 81.545 140.330 ;
        RECT 80.065 134.610 80.345 134.890 ;
        RECT 80.465 134.610 80.745 134.890 ;
        RECT 80.865 134.610 81.145 134.890 ;
        RECT 81.265 134.610 81.545 134.890 ;
        RECT 92.170 179.150 92.450 179.430 ;
        RECT 97.490 197.170 97.770 197.450 ;
        RECT 97.890 197.170 98.170 197.450 ;
        RECT 98.290 197.170 98.570 197.450 ;
        RECT 98.690 197.170 98.970 197.450 ;
        RECT 97.490 191.730 97.770 192.010 ;
        RECT 97.890 191.730 98.170 192.010 ;
        RECT 98.290 191.730 98.570 192.010 ;
        RECT 98.690 191.730 98.970 192.010 ;
        RECT 94.930 187.310 95.210 187.590 ;
        RECT 97.490 186.290 97.770 186.570 ;
        RECT 97.890 186.290 98.170 186.570 ;
        RECT 98.290 186.290 98.570 186.570 ;
        RECT 98.690 186.290 98.970 186.570 ;
        RECT 101.370 198.870 101.650 199.150 ;
        RECT 97.490 180.850 97.770 181.130 ;
        RECT 97.890 180.850 98.170 181.130 ;
        RECT 98.290 180.850 98.570 181.130 ;
        RECT 98.690 180.850 98.970 181.130 ;
        RECT 97.490 175.410 97.770 175.690 ;
        RECT 97.890 175.410 98.170 175.690 ;
        RECT 98.290 175.410 98.570 175.690 ;
        RECT 98.690 175.410 98.970 175.690 ;
        RECT 97.490 169.970 97.770 170.250 ;
        RECT 97.890 169.970 98.170 170.250 ;
        RECT 98.290 169.970 98.570 170.250 ;
        RECT 98.690 169.970 98.970 170.250 ;
        RECT 92.630 157.390 92.910 157.670 ;
        RECT 87.110 152.630 87.390 152.910 ;
        RECT 88.030 151.950 88.310 152.230 ;
        RECT 97.490 164.530 97.770 164.810 ;
        RECT 97.890 164.530 98.170 164.810 ;
        RECT 98.290 164.530 98.570 164.810 ;
        RECT 98.690 164.530 98.970 164.810 ;
        RECT 102.290 187.310 102.570 187.590 ;
        RECT 97.490 159.090 97.770 159.370 ;
        RECT 97.890 159.090 98.170 159.370 ;
        RECT 98.290 159.090 98.570 159.370 ;
        RECT 98.690 159.090 98.970 159.370 ;
        RECT 97.490 153.650 97.770 153.930 ;
        RECT 97.890 153.650 98.170 153.930 ;
        RECT 98.290 153.650 98.570 153.930 ;
        RECT 98.690 153.650 98.970 153.930 ;
        RECT 97.230 152.630 97.510 152.910 ;
        RECT 97.690 151.950 97.970 152.230 ;
        RECT 97.490 148.210 97.770 148.490 ;
        RECT 97.890 148.210 98.170 148.490 ;
        RECT 98.290 148.210 98.570 148.490 ;
        RECT 98.690 148.210 98.970 148.490 ;
        RECT 114.910 205.330 115.190 205.610 ;
        RECT 115.310 205.330 115.590 205.610 ;
        RECT 115.710 205.330 115.990 205.610 ;
        RECT 116.110 205.330 116.390 205.610 ;
        RECT 132.335 208.050 132.615 208.330 ;
        RECT 132.735 208.050 133.015 208.330 ;
        RECT 133.135 208.050 133.415 208.330 ;
        RECT 133.535 208.050 133.815 208.330 ;
        RECT 114.910 199.890 115.190 200.170 ;
        RECT 115.310 199.890 115.590 200.170 ;
        RECT 115.710 199.890 115.990 200.170 ;
        RECT 116.110 199.890 116.390 200.170 ;
        RECT 97.490 142.770 97.770 143.050 ;
        RECT 97.890 142.770 98.170 143.050 ;
        RECT 98.290 142.770 98.570 143.050 ;
        RECT 98.690 142.770 98.970 143.050 ;
        RECT 80.065 129.170 80.345 129.450 ;
        RECT 80.465 129.170 80.745 129.450 ;
        RECT 80.865 129.170 81.145 129.450 ;
        RECT 81.265 129.170 81.545 129.450 ;
        RECT 83.430 134.950 83.710 135.230 ;
        RECT 89.870 136.310 90.150 136.590 ;
        RECT 114.910 194.450 115.190 194.730 ;
        RECT 115.310 194.450 115.590 194.730 ;
        RECT 115.710 194.450 115.990 194.730 ;
        RECT 116.110 194.450 116.390 194.730 ;
        RECT 114.910 189.010 115.190 189.290 ;
        RECT 115.310 189.010 115.590 189.290 ;
        RECT 115.710 189.010 115.990 189.290 ;
        RECT 116.110 189.010 116.390 189.290 ;
        RECT 113.790 182.550 114.070 182.830 ;
        RECT 114.910 183.570 115.190 183.850 ;
        RECT 115.310 183.570 115.590 183.850 ;
        RECT 115.710 183.570 115.990 183.850 ;
        RECT 116.110 183.570 116.390 183.850 ;
        RECT 114.910 178.130 115.190 178.410 ;
        RECT 115.310 178.130 115.590 178.410 ;
        RECT 115.710 178.130 115.990 178.410 ;
        RECT 116.110 178.130 116.390 178.410 ;
        RECT 122.990 187.990 123.270 188.270 ;
        RECT 114.910 172.690 115.190 172.970 ;
        RECT 115.310 172.690 115.590 172.970 ;
        RECT 115.710 172.690 115.990 172.970 ;
        RECT 116.110 172.690 116.390 172.970 ;
        RECT 116.090 168.270 116.370 168.550 ;
        RECT 114.910 167.250 115.190 167.530 ;
        RECT 115.310 167.250 115.590 167.530 ;
        RECT 115.710 167.250 115.990 167.530 ;
        RECT 116.110 167.250 116.390 167.530 ;
        RECT 97.490 137.330 97.770 137.610 ;
        RECT 97.890 137.330 98.170 137.610 ;
        RECT 98.290 137.330 98.570 137.610 ;
        RECT 98.690 137.330 98.970 137.610 ;
        RECT 97.490 131.890 97.770 132.170 ;
        RECT 97.890 131.890 98.170 132.170 ;
        RECT 98.290 131.890 98.570 132.170 ;
        RECT 98.690 131.890 98.970 132.170 ;
        RECT 114.910 161.810 115.190 162.090 ;
        RECT 115.310 161.810 115.590 162.090 ;
        RECT 115.710 161.810 115.990 162.090 ;
        RECT 116.110 161.810 116.390 162.090 ;
        RECT 114.910 156.370 115.190 156.650 ;
        RECT 115.310 156.370 115.590 156.650 ;
        RECT 115.710 156.370 115.990 156.650 ;
        RECT 116.110 156.370 116.390 156.650 ;
        RECT 114.910 150.930 115.190 151.210 ;
        RECT 115.310 150.930 115.590 151.210 ;
        RECT 115.710 150.930 115.990 151.210 ;
        RECT 116.110 150.930 116.390 151.210 ;
        RECT 114.910 145.490 115.190 145.770 ;
        RECT 115.310 145.490 115.590 145.770 ;
        RECT 115.710 145.490 115.990 145.770 ;
        RECT 116.110 145.490 116.390 145.770 ;
        RECT 114.910 140.050 115.190 140.330 ;
        RECT 115.310 140.050 115.590 140.330 ;
        RECT 115.710 140.050 115.990 140.330 ;
        RECT 116.110 140.050 116.390 140.330 ;
        RECT 125.750 182.550 126.030 182.830 ;
        RECT 132.335 202.610 132.615 202.890 ;
        RECT 132.735 202.610 133.015 202.890 ;
        RECT 133.135 202.610 133.415 202.890 ;
        RECT 133.535 202.610 133.815 202.890 ;
        RECT 132.335 197.170 132.615 197.450 ;
        RECT 132.735 197.170 133.015 197.450 ;
        RECT 133.135 197.170 133.415 197.450 ;
        RECT 133.535 197.170 133.815 197.450 ;
        RECT 132.335 191.730 132.615 192.010 ;
        RECT 132.735 191.730 133.015 192.010 ;
        RECT 133.135 191.730 133.415 192.010 ;
        RECT 133.535 191.730 133.815 192.010 ;
        RECT 132.335 186.290 132.615 186.570 ;
        RECT 132.735 186.290 133.015 186.570 ;
        RECT 133.135 186.290 133.415 186.570 ;
        RECT 133.535 186.290 133.815 186.570 ;
        RECT 132.335 180.850 132.615 181.130 ;
        RECT 132.735 180.850 133.015 181.130 ;
        RECT 133.135 180.850 133.415 181.130 ;
        RECT 133.535 180.850 133.815 181.130 ;
        RECT 132.335 175.410 132.615 175.690 ;
        RECT 132.735 175.410 133.015 175.690 ;
        RECT 133.135 175.410 133.415 175.690 ;
        RECT 133.535 175.410 133.815 175.690 ;
        RECT 132.335 169.970 132.615 170.250 ;
        RECT 132.735 169.970 133.015 170.250 ;
        RECT 133.135 169.970 133.415 170.250 ;
        RECT 133.535 169.970 133.815 170.250 ;
        RECT 149.755 210.770 150.035 211.050 ;
        RECT 150.155 210.770 150.435 211.050 ;
        RECT 150.555 210.770 150.835 211.050 ;
        RECT 150.955 210.770 151.235 211.050 ;
        RECT 149.755 205.330 150.035 205.610 ;
        RECT 150.155 205.330 150.435 205.610 ;
        RECT 150.555 205.330 150.835 205.610 ;
        RECT 150.955 205.330 151.235 205.610 ;
        RECT 149.755 199.890 150.035 200.170 ;
        RECT 150.155 199.890 150.435 200.170 ;
        RECT 150.555 199.890 150.835 200.170 ;
        RECT 150.955 199.890 151.235 200.170 ;
        RECT 149.755 194.450 150.035 194.730 ;
        RECT 150.155 194.450 150.435 194.730 ;
        RECT 150.555 194.450 150.835 194.730 ;
        RECT 150.955 194.450 151.235 194.730 ;
        RECT 149.755 189.010 150.035 189.290 ;
        RECT 150.155 189.010 150.435 189.290 ;
        RECT 150.555 189.010 150.835 189.290 ;
        RECT 150.955 189.010 151.235 189.290 ;
        RECT 149.755 183.570 150.035 183.850 ;
        RECT 150.155 183.570 150.435 183.850 ;
        RECT 150.555 183.570 150.835 183.850 ;
        RECT 150.955 183.570 151.235 183.850 ;
        RECT 149.755 178.130 150.035 178.410 ;
        RECT 150.155 178.130 150.435 178.410 ;
        RECT 150.555 178.130 150.835 178.410 ;
        RECT 150.955 178.130 151.235 178.410 ;
        RECT 149.755 172.690 150.035 172.970 ;
        RECT 150.155 172.690 150.435 172.970 ;
        RECT 150.555 172.690 150.835 172.970 ;
        RECT 150.955 172.690 151.235 172.970 ;
        RECT 146.450 168.270 146.730 168.550 ;
        RECT 149.755 167.250 150.035 167.530 ;
        RECT 150.155 167.250 150.435 167.530 ;
        RECT 150.555 167.250 150.835 167.530 ;
        RECT 150.955 167.250 151.235 167.530 ;
        RECT 132.335 164.530 132.615 164.810 ;
        RECT 132.735 164.530 133.015 164.810 ;
        RECT 133.135 164.530 133.415 164.810 ;
        RECT 133.535 164.530 133.815 164.810 ;
        RECT 149.755 161.810 150.035 162.090 ;
        RECT 150.155 161.810 150.435 162.090 ;
        RECT 150.555 161.810 150.835 162.090 ;
        RECT 150.955 161.810 151.235 162.090 ;
        RECT 132.335 159.090 132.615 159.370 ;
        RECT 132.735 159.090 133.015 159.370 ;
        RECT 133.135 159.090 133.415 159.370 ;
        RECT 133.535 159.090 133.815 159.370 ;
        RECT 149.755 156.370 150.035 156.650 ;
        RECT 150.155 156.370 150.435 156.650 ;
        RECT 150.555 156.370 150.835 156.650 ;
        RECT 150.955 156.370 151.235 156.650 ;
        RECT 132.335 153.650 132.615 153.930 ;
        RECT 132.735 153.650 133.015 153.930 ;
        RECT 133.135 153.650 133.415 153.930 ;
        RECT 133.535 153.650 133.815 153.930 ;
        RECT 149.755 150.930 150.035 151.210 ;
        RECT 150.155 150.930 150.435 151.210 ;
        RECT 150.555 150.930 150.835 151.210 ;
        RECT 150.955 150.930 151.235 151.210 ;
        RECT 132.335 148.210 132.615 148.490 ;
        RECT 132.735 148.210 133.015 148.490 ;
        RECT 133.135 148.210 133.415 148.490 ;
        RECT 133.535 148.210 133.815 148.490 ;
        RECT 149.755 145.490 150.035 145.770 ;
        RECT 150.155 145.490 150.435 145.770 ;
        RECT 150.555 145.490 150.835 145.770 ;
        RECT 150.955 145.490 151.235 145.770 ;
        RECT 132.335 142.770 132.615 143.050 ;
        RECT 132.735 142.770 133.015 143.050 ;
        RECT 133.135 142.770 133.415 143.050 ;
        RECT 133.535 142.770 133.815 143.050 ;
        RECT 114.910 134.610 115.190 134.890 ;
        RECT 115.310 134.610 115.590 134.890 ;
        RECT 115.710 134.610 115.990 134.890 ;
        RECT 116.110 134.610 116.390 134.890 ;
        RECT 149.755 140.050 150.035 140.330 ;
        RECT 150.155 140.050 150.435 140.330 ;
        RECT 150.555 140.050 150.835 140.330 ;
        RECT 150.955 140.050 151.235 140.330 ;
        RECT 132.335 137.330 132.615 137.610 ;
        RECT 132.735 137.330 133.015 137.610 ;
        RECT 133.135 137.330 133.415 137.610 ;
        RECT 133.535 137.330 133.815 137.610 ;
        RECT 149.755 134.610 150.035 134.890 ;
        RECT 150.155 134.610 150.435 134.890 ;
        RECT 150.555 134.610 150.835 134.890 ;
        RECT 150.955 134.610 151.235 134.890 ;
        RECT 132.335 131.890 132.615 132.170 ;
        RECT 132.735 131.890 133.015 132.170 ;
        RECT 133.135 131.890 133.415 132.170 ;
        RECT 133.535 131.890 133.815 132.170 ;
        RECT 114.910 129.170 115.190 129.450 ;
        RECT 115.310 129.170 115.590 129.450 ;
        RECT 115.710 129.170 115.990 129.450 ;
        RECT 116.110 129.170 116.390 129.450 ;
        RECT 149.755 129.170 150.035 129.450 ;
        RECT 150.155 129.170 150.435 129.450 ;
        RECT 150.555 129.170 150.835 129.450 ;
        RECT 150.955 129.170 151.235 129.450 ;
        RECT 97.490 126.450 97.770 126.730 ;
        RECT 97.890 126.450 98.170 126.730 ;
        RECT 98.290 126.450 98.570 126.730 ;
        RECT 98.690 126.450 98.970 126.730 ;
        RECT 132.335 126.450 132.615 126.730 ;
        RECT 132.735 126.450 133.015 126.730 ;
        RECT 133.135 126.450 133.415 126.730 ;
        RECT 133.535 126.450 133.815 126.730 ;
        RECT 80.065 123.730 80.345 124.010 ;
        RECT 80.465 123.730 80.745 124.010 ;
        RECT 80.865 123.730 81.145 124.010 ;
        RECT 81.265 123.730 81.545 124.010 ;
        RECT 114.910 123.730 115.190 124.010 ;
        RECT 115.310 123.730 115.590 124.010 ;
        RECT 115.710 123.730 115.990 124.010 ;
        RECT 116.110 123.730 116.390 124.010 ;
        RECT 149.755 123.730 150.035 124.010 ;
        RECT 150.155 123.730 150.435 124.010 ;
        RECT 150.555 123.730 150.835 124.010 ;
        RECT 150.955 123.730 151.235 124.010 ;
        RECT 27.800 121.010 28.080 121.290 ;
        RECT 28.200 121.010 28.480 121.290 ;
        RECT 28.600 121.010 28.880 121.290 ;
        RECT 29.000 121.010 29.280 121.290 ;
        RECT 62.645 121.010 62.925 121.290 ;
        RECT 63.045 121.010 63.325 121.290 ;
        RECT 63.445 121.010 63.725 121.290 ;
        RECT 63.845 121.010 64.125 121.290 ;
        RECT 97.490 121.010 97.770 121.290 ;
        RECT 97.890 121.010 98.170 121.290 ;
        RECT 98.290 121.010 98.570 121.290 ;
        RECT 98.690 121.010 98.970 121.290 ;
        RECT 132.335 121.010 132.615 121.290 ;
        RECT 132.735 121.010 133.015 121.290 ;
        RECT 133.135 121.010 133.415 121.290 ;
        RECT 133.535 121.010 133.815 121.290 ;
        RECT 45.220 118.290 45.500 118.570 ;
        RECT 45.620 118.290 45.900 118.570 ;
        RECT 46.020 118.290 46.300 118.570 ;
        RECT 46.420 118.290 46.700 118.570 ;
        RECT 80.065 118.290 80.345 118.570 ;
        RECT 80.465 118.290 80.745 118.570 ;
        RECT 80.865 118.290 81.145 118.570 ;
        RECT 81.265 118.290 81.545 118.570 ;
        RECT 114.910 118.290 115.190 118.570 ;
        RECT 115.310 118.290 115.590 118.570 ;
        RECT 115.710 118.290 115.990 118.570 ;
        RECT 116.110 118.290 116.390 118.570 ;
        RECT 149.755 118.290 150.035 118.570 ;
        RECT 150.155 118.290 150.435 118.570 ;
        RECT 150.555 118.290 150.835 118.570 ;
        RECT 150.955 118.290 151.235 118.570 ;
        RECT 27.800 115.570 28.080 115.850 ;
        RECT 28.200 115.570 28.480 115.850 ;
        RECT 28.600 115.570 28.880 115.850 ;
        RECT 29.000 115.570 29.280 115.850 ;
        RECT 62.645 115.570 62.925 115.850 ;
        RECT 63.045 115.570 63.325 115.850 ;
        RECT 63.445 115.570 63.725 115.850 ;
        RECT 63.845 115.570 64.125 115.850 ;
        RECT 97.490 115.570 97.770 115.850 ;
        RECT 97.890 115.570 98.170 115.850 ;
        RECT 98.290 115.570 98.570 115.850 ;
        RECT 98.690 115.570 98.970 115.850 ;
        RECT 132.335 115.570 132.615 115.850 ;
        RECT 132.735 115.570 133.015 115.850 ;
        RECT 133.135 115.570 133.415 115.850 ;
        RECT 133.535 115.570 133.815 115.850 ;
        RECT 45.220 112.850 45.500 113.130 ;
        RECT 45.620 112.850 45.900 113.130 ;
        RECT 46.020 112.850 46.300 113.130 ;
        RECT 46.420 112.850 46.700 113.130 ;
        RECT 80.065 112.850 80.345 113.130 ;
        RECT 80.465 112.850 80.745 113.130 ;
        RECT 80.865 112.850 81.145 113.130 ;
        RECT 81.265 112.850 81.545 113.130 ;
        RECT 114.910 112.850 115.190 113.130 ;
        RECT 115.310 112.850 115.590 113.130 ;
        RECT 115.710 112.850 115.990 113.130 ;
        RECT 116.110 112.850 116.390 113.130 ;
        RECT 149.755 112.850 150.035 113.130 ;
        RECT 150.155 112.850 150.435 113.130 ;
        RECT 150.555 112.850 150.835 113.130 ;
        RECT 150.955 112.850 151.235 113.130 ;
        RECT 27.800 110.130 28.080 110.410 ;
        RECT 28.200 110.130 28.480 110.410 ;
        RECT 28.600 110.130 28.880 110.410 ;
        RECT 29.000 110.130 29.280 110.410 ;
        RECT 62.645 110.130 62.925 110.410 ;
        RECT 63.045 110.130 63.325 110.410 ;
        RECT 63.445 110.130 63.725 110.410 ;
        RECT 63.845 110.130 64.125 110.410 ;
        RECT 97.490 110.130 97.770 110.410 ;
        RECT 97.890 110.130 98.170 110.410 ;
        RECT 98.290 110.130 98.570 110.410 ;
        RECT 98.690 110.130 98.970 110.410 ;
        RECT 132.335 110.130 132.615 110.410 ;
        RECT 132.735 110.130 133.015 110.410 ;
        RECT 133.135 110.130 133.415 110.410 ;
        RECT 133.535 110.130 133.815 110.410 ;
        RECT 45.220 107.410 45.500 107.690 ;
        RECT 45.620 107.410 45.900 107.690 ;
        RECT 46.020 107.410 46.300 107.690 ;
        RECT 46.420 107.410 46.700 107.690 ;
        RECT 80.065 107.410 80.345 107.690 ;
        RECT 80.465 107.410 80.745 107.690 ;
        RECT 80.865 107.410 81.145 107.690 ;
        RECT 81.265 107.410 81.545 107.690 ;
        RECT 114.910 107.410 115.190 107.690 ;
        RECT 115.310 107.410 115.590 107.690 ;
        RECT 115.710 107.410 115.990 107.690 ;
        RECT 116.110 107.410 116.390 107.690 ;
        RECT 149.755 107.410 150.035 107.690 ;
        RECT 150.155 107.410 150.435 107.690 ;
        RECT 150.555 107.410 150.835 107.690 ;
        RECT 150.955 107.410 151.235 107.690 ;
        RECT 27.800 104.690 28.080 104.970 ;
        RECT 28.200 104.690 28.480 104.970 ;
        RECT 28.600 104.690 28.880 104.970 ;
        RECT 29.000 104.690 29.280 104.970 ;
        RECT 62.645 104.690 62.925 104.970 ;
        RECT 63.045 104.690 63.325 104.970 ;
        RECT 63.445 104.690 63.725 104.970 ;
        RECT 63.845 104.690 64.125 104.970 ;
        RECT 97.490 104.690 97.770 104.970 ;
        RECT 97.890 104.690 98.170 104.970 ;
        RECT 98.290 104.690 98.570 104.970 ;
        RECT 98.690 104.690 98.970 104.970 ;
        RECT 132.335 104.690 132.615 104.970 ;
        RECT 132.735 104.690 133.015 104.970 ;
        RECT 133.135 104.690 133.415 104.970 ;
        RECT 133.535 104.690 133.815 104.970 ;
        RECT 45.220 101.970 45.500 102.250 ;
        RECT 45.620 101.970 45.900 102.250 ;
        RECT 46.020 101.970 46.300 102.250 ;
        RECT 46.420 101.970 46.700 102.250 ;
        RECT 80.065 101.970 80.345 102.250 ;
        RECT 80.465 101.970 80.745 102.250 ;
        RECT 80.865 101.970 81.145 102.250 ;
        RECT 81.265 101.970 81.545 102.250 ;
        RECT 114.910 101.970 115.190 102.250 ;
        RECT 115.310 101.970 115.590 102.250 ;
        RECT 115.710 101.970 115.990 102.250 ;
        RECT 116.110 101.970 116.390 102.250 ;
        RECT 149.755 101.970 150.035 102.250 ;
        RECT 150.155 101.970 150.435 102.250 ;
        RECT 150.555 101.970 150.835 102.250 ;
        RECT 150.955 101.970 151.235 102.250 ;
        RECT 27.800 99.250 28.080 99.530 ;
        RECT 28.200 99.250 28.480 99.530 ;
        RECT 28.600 99.250 28.880 99.530 ;
        RECT 29.000 99.250 29.280 99.530 ;
        RECT 62.645 99.250 62.925 99.530 ;
        RECT 63.045 99.250 63.325 99.530 ;
        RECT 63.445 99.250 63.725 99.530 ;
        RECT 63.845 99.250 64.125 99.530 ;
        RECT 97.490 99.250 97.770 99.530 ;
        RECT 97.890 99.250 98.170 99.530 ;
        RECT 98.290 99.250 98.570 99.530 ;
        RECT 98.690 99.250 98.970 99.530 ;
        RECT 132.335 99.250 132.615 99.530 ;
        RECT 132.735 99.250 133.015 99.530 ;
        RECT 133.135 99.250 133.415 99.530 ;
        RECT 133.535 99.250 133.815 99.530 ;
        RECT 45.220 96.530 45.500 96.810 ;
        RECT 45.620 96.530 45.900 96.810 ;
        RECT 46.020 96.530 46.300 96.810 ;
        RECT 46.420 96.530 46.700 96.810 ;
        RECT 80.065 96.530 80.345 96.810 ;
        RECT 80.465 96.530 80.745 96.810 ;
        RECT 80.865 96.530 81.145 96.810 ;
        RECT 81.265 96.530 81.545 96.810 ;
        RECT 114.910 96.530 115.190 96.810 ;
        RECT 115.310 96.530 115.590 96.810 ;
        RECT 115.710 96.530 115.990 96.810 ;
        RECT 116.110 96.530 116.390 96.810 ;
        RECT 149.755 96.530 150.035 96.810 ;
        RECT 150.155 96.530 150.435 96.810 ;
        RECT 150.555 96.530 150.835 96.810 ;
        RECT 150.955 96.530 151.235 96.810 ;
        RECT 27.800 93.810 28.080 94.090 ;
        RECT 28.200 93.810 28.480 94.090 ;
        RECT 28.600 93.810 28.880 94.090 ;
        RECT 29.000 93.810 29.280 94.090 ;
        RECT 62.645 93.810 62.925 94.090 ;
        RECT 63.045 93.810 63.325 94.090 ;
        RECT 63.445 93.810 63.725 94.090 ;
        RECT 63.845 93.810 64.125 94.090 ;
        RECT 97.490 93.810 97.770 94.090 ;
        RECT 97.890 93.810 98.170 94.090 ;
        RECT 98.290 93.810 98.570 94.090 ;
        RECT 98.690 93.810 98.970 94.090 ;
        RECT 132.335 93.810 132.615 94.090 ;
        RECT 132.735 93.810 133.015 94.090 ;
        RECT 133.135 93.810 133.415 94.090 ;
        RECT 133.535 93.810 133.815 94.090 ;
        RECT 45.220 91.090 45.500 91.370 ;
        RECT 45.620 91.090 45.900 91.370 ;
        RECT 46.020 91.090 46.300 91.370 ;
        RECT 46.420 91.090 46.700 91.370 ;
        RECT 80.065 91.090 80.345 91.370 ;
        RECT 80.465 91.090 80.745 91.370 ;
        RECT 80.865 91.090 81.145 91.370 ;
        RECT 81.265 91.090 81.545 91.370 ;
        RECT 114.910 91.090 115.190 91.370 ;
        RECT 115.310 91.090 115.590 91.370 ;
        RECT 115.710 91.090 115.990 91.370 ;
        RECT 116.110 91.090 116.390 91.370 ;
        RECT 149.755 91.090 150.035 91.370 ;
        RECT 150.155 91.090 150.435 91.370 ;
        RECT 150.555 91.090 150.835 91.370 ;
        RECT 150.955 91.090 151.235 91.370 ;
        RECT 27.800 88.370 28.080 88.650 ;
        RECT 28.200 88.370 28.480 88.650 ;
        RECT 28.600 88.370 28.880 88.650 ;
        RECT 29.000 88.370 29.280 88.650 ;
        RECT 62.645 88.370 62.925 88.650 ;
        RECT 63.045 88.370 63.325 88.650 ;
        RECT 63.445 88.370 63.725 88.650 ;
        RECT 63.845 88.370 64.125 88.650 ;
        RECT 97.490 88.370 97.770 88.650 ;
        RECT 97.890 88.370 98.170 88.650 ;
        RECT 98.290 88.370 98.570 88.650 ;
        RECT 98.690 88.370 98.970 88.650 ;
        RECT 132.335 88.370 132.615 88.650 ;
        RECT 132.735 88.370 133.015 88.650 ;
        RECT 133.135 88.370 133.415 88.650 ;
        RECT 133.535 88.370 133.815 88.650 ;
        RECT 45.220 85.650 45.500 85.930 ;
        RECT 45.620 85.650 45.900 85.930 ;
        RECT 46.020 85.650 46.300 85.930 ;
        RECT 46.420 85.650 46.700 85.930 ;
        RECT 80.065 85.650 80.345 85.930 ;
        RECT 80.465 85.650 80.745 85.930 ;
        RECT 80.865 85.650 81.145 85.930 ;
        RECT 81.265 85.650 81.545 85.930 ;
        RECT 114.910 85.650 115.190 85.930 ;
        RECT 115.310 85.650 115.590 85.930 ;
        RECT 115.710 85.650 115.990 85.930 ;
        RECT 116.110 85.650 116.390 85.930 ;
        RECT 149.755 85.650 150.035 85.930 ;
        RECT 150.155 85.650 150.435 85.930 ;
        RECT 150.555 85.650 150.835 85.930 ;
        RECT 150.955 85.650 151.235 85.930 ;
        RECT 27.800 82.930 28.080 83.210 ;
        RECT 28.200 82.930 28.480 83.210 ;
        RECT 28.600 82.930 28.880 83.210 ;
        RECT 29.000 82.930 29.280 83.210 ;
        RECT 62.645 82.930 62.925 83.210 ;
        RECT 63.045 82.930 63.325 83.210 ;
        RECT 63.445 82.930 63.725 83.210 ;
        RECT 63.845 82.930 64.125 83.210 ;
        RECT 97.490 82.930 97.770 83.210 ;
        RECT 97.890 82.930 98.170 83.210 ;
        RECT 98.290 82.930 98.570 83.210 ;
        RECT 98.690 82.930 98.970 83.210 ;
        RECT 132.335 82.930 132.615 83.210 ;
        RECT 132.735 82.930 133.015 83.210 ;
        RECT 133.135 82.930 133.415 83.210 ;
        RECT 133.535 82.930 133.815 83.210 ;
        RECT 45.220 80.210 45.500 80.490 ;
        RECT 45.620 80.210 45.900 80.490 ;
        RECT 46.020 80.210 46.300 80.490 ;
        RECT 46.420 80.210 46.700 80.490 ;
        RECT 80.065 80.210 80.345 80.490 ;
        RECT 80.465 80.210 80.745 80.490 ;
        RECT 80.865 80.210 81.145 80.490 ;
        RECT 81.265 80.210 81.545 80.490 ;
        RECT 114.910 80.210 115.190 80.490 ;
        RECT 115.310 80.210 115.590 80.490 ;
        RECT 115.710 80.210 115.990 80.490 ;
        RECT 116.110 80.210 116.390 80.490 ;
        RECT 149.755 80.210 150.035 80.490 ;
        RECT 150.155 80.210 150.435 80.490 ;
        RECT 150.555 80.210 150.835 80.490 ;
        RECT 150.955 80.210 151.235 80.490 ;
        RECT 27.800 77.490 28.080 77.770 ;
        RECT 28.200 77.490 28.480 77.770 ;
        RECT 28.600 77.490 28.880 77.770 ;
        RECT 29.000 77.490 29.280 77.770 ;
        RECT 62.645 77.490 62.925 77.770 ;
        RECT 63.045 77.490 63.325 77.770 ;
        RECT 63.445 77.490 63.725 77.770 ;
        RECT 63.845 77.490 64.125 77.770 ;
        RECT 97.490 77.490 97.770 77.770 ;
        RECT 97.890 77.490 98.170 77.770 ;
        RECT 98.290 77.490 98.570 77.770 ;
        RECT 98.690 77.490 98.970 77.770 ;
        RECT 132.335 77.490 132.615 77.770 ;
        RECT 132.735 77.490 133.015 77.770 ;
        RECT 133.135 77.490 133.415 77.770 ;
        RECT 133.535 77.490 133.815 77.770 ;
        RECT 45.220 74.770 45.500 75.050 ;
        RECT 45.620 74.770 45.900 75.050 ;
        RECT 46.020 74.770 46.300 75.050 ;
        RECT 46.420 74.770 46.700 75.050 ;
        RECT 80.065 74.770 80.345 75.050 ;
        RECT 80.465 74.770 80.745 75.050 ;
        RECT 80.865 74.770 81.145 75.050 ;
        RECT 81.265 74.770 81.545 75.050 ;
        RECT 114.910 74.770 115.190 75.050 ;
        RECT 115.310 74.770 115.590 75.050 ;
        RECT 115.710 74.770 115.990 75.050 ;
        RECT 116.110 74.770 116.390 75.050 ;
        RECT 149.755 74.770 150.035 75.050 ;
        RECT 150.155 74.770 150.435 75.050 ;
        RECT 150.555 74.770 150.835 75.050 ;
        RECT 150.955 74.770 151.235 75.050 ;
        RECT 55.340 55.020 76.610 59.300 ;
        RECT 95.400 55.090 105.220 59.770 ;
        RECT 62.000 49.290 62.940 49.650 ;
        RECT 64.680 49.300 65.590 49.700 ;
        RECT 78.760 49.160 79.750 49.640 ;
        RECT 117.310 54.830 134.530 58.370 ;
        RECT 124.230 48.890 125.170 49.250 ;
        RECT 126.910 48.900 127.820 49.300 ;
        RECT 140.990 48.760 141.980 49.240 ;
        RECT 78.750 47.580 79.740 48.060 ;
        RECT 62.000 44.650 62.940 45.010 ;
        RECT 64.680 44.630 65.590 45.030 ;
        RECT 140.980 47.180 141.970 47.660 ;
        RECT 78.740 46.010 79.730 46.490 ;
        RECT 78.770 44.420 79.760 44.900 ;
        RECT 124.230 44.250 125.170 44.610 ;
        RECT 126.910 44.230 127.820 44.630 ;
        RECT 78.770 42.840 79.760 43.320 ;
        RECT 62.010 40.080 62.950 40.440 ;
        RECT 64.670 40.060 65.580 40.460 ;
        RECT 73.590 39.820 74.540 40.100 ;
        RECT 78.770 41.260 79.760 41.740 ;
        RECT 140.970 45.610 141.960 46.090 ;
        RECT 141.000 44.020 141.990 44.500 ;
        RECT 141.000 42.440 141.990 42.920 ;
        RECT 78.750 39.680 79.740 40.160 ;
        RECT 78.760 38.100 79.750 38.580 ;
        RECT 62.030 35.540 62.940 35.840 ;
        RECT 64.690 35.490 65.590 35.840 ;
        RECT 73.580 35.110 74.540 35.620 ;
        RECT 78.770 36.520 79.760 37.000 ;
        RECT 78.770 34.950 79.760 35.430 ;
        RECT 78.760 33.230 79.700 33.800 ;
        RECT 73.580 30.570 74.540 30.990 ;
        RECT 73.590 26.050 74.540 26.390 ;
        RECT 124.240 39.680 125.180 40.040 ;
        RECT 126.900 39.660 127.810 40.060 ;
        RECT 135.820 39.420 136.770 39.700 ;
        RECT 141.000 40.860 141.990 41.340 ;
        RECT 140.980 39.280 141.970 39.760 ;
        RECT 140.990 37.700 141.980 38.180 ;
        RECT 124.260 35.140 125.170 35.440 ;
        RECT 126.920 35.090 127.820 35.440 ;
        RECT 135.810 34.710 136.770 35.220 ;
        RECT 141.000 36.120 141.990 36.600 ;
        RECT 141.000 34.550 141.990 35.030 ;
        RECT 140.990 32.830 141.930 33.400 ;
        RECT 135.810 30.170 136.770 30.590 ;
        RECT 107.250 25.590 108.070 26.410 ;
        RECT 90.345 23.155 90.895 23.705 ;
        RECT 60.015 20.945 60.885 21.815 ;
        RECT 55.390 11.400 64.190 18.240 ;
        RECT 135.820 25.650 136.770 25.990 ;
        RECT 74.330 11.280 83.680 18.120 ;
        RECT 94.640 11.670 105.730 18.200 ;
        RECT 117.320 13.120 127.600 18.610 ;
        RECT 69.475 7.425 70.025 7.975 ;
        RECT 134.505 20.035 135.055 20.585 ;
        RECT 150.555 20.185 151.105 20.735 ;
        RECT 135.980 13.520 146.160 18.400 ;
        RECT 128.995 6.615 129.545 7.165 ;
        RECT 56.435 4.805 56.985 5.355 ;
      LAYER met3 ;
        RECT 57.765 223.720 58.115 223.745 ;
        RECT 59.990 223.720 60.370 223.730 ;
        RECT 57.765 223.420 60.370 223.720 ;
        RECT 74.950 223.580 75.330 223.900 ;
        RECT 126.925 223.890 127.275 223.915 ;
        RECT 129.530 223.890 129.910 223.900 ;
        RECT 126.925 223.590 129.910 223.890 ;
        RECT 57.765 223.395 58.115 223.420 ;
        RECT 59.990 223.410 60.370 223.420 ;
        RECT 70.220 221.860 70.540 221.900 ;
        RECT 35.120 221.560 70.540 221.860 ;
        RECT 24.990 218.480 25.310 218.860 ;
        RECT 25.000 216.475 25.300 218.480 ;
        RECT 35.120 216.895 35.420 221.560 ;
        RECT 70.220 221.520 70.540 221.560 ;
        RECT 73.870 221.480 74.190 221.860 ;
        RECT 73.880 220.905 74.180 221.480 ;
        RECT 73.855 220.555 74.205 220.905 ;
        RECT 74.990 219.890 75.290 223.580 ;
        RECT 126.925 223.565 127.275 223.590 ;
        RECT 129.530 223.580 129.910 223.590 ;
        RECT 143.800 222.460 144.120 222.840 ;
        RECT 143.810 221.445 144.110 222.460 ;
        RECT 151.180 222.240 151.500 222.620 ;
        RECT 143.785 221.095 144.135 221.445 ;
        RECT 151.190 220.385 151.490 222.240 ;
        RECT 60.600 219.590 75.290 219.890 ;
        RECT 105.950 219.810 106.270 220.190 ;
        RECT 151.165 220.035 151.515 220.385 ;
        RECT 55.335 217.400 55.685 217.425 ;
        RECT 60.600 217.400 60.900 219.590 ;
        RECT 85.695 218.750 86.045 218.775 ;
        RECT 87.150 218.750 87.530 218.760 ;
        RECT 85.695 218.450 87.530 218.750 ;
        RECT 85.695 218.425 86.045 218.450 ;
        RECT 87.150 218.440 87.530 218.450 ;
        RECT 105.960 218.165 106.260 219.810 ;
        RECT 126.190 219.230 126.510 219.610 ;
        RECT 126.200 218.535 126.500 219.230 ;
        RECT 126.175 218.185 126.525 218.535 ;
        RECT 79.555 218.040 79.905 218.065 ;
        RECT 83.810 218.040 84.130 218.080 ;
        RECT 79.555 217.740 84.130 218.040 ;
        RECT 105.935 217.815 106.285 218.165 ;
        RECT 79.555 217.715 79.905 217.740 ;
        RECT 83.810 217.700 84.130 217.740 ;
        RECT 146.415 217.700 146.765 217.725 ;
        RECT 153.620 217.700 154.000 217.710 ;
        RECT 35.095 216.545 35.445 216.895 ;
        RECT 24.975 216.125 25.325 216.475 ;
        RECT 45.240 216.075 45.540 217.200 ;
        RECT 55.335 217.100 60.900 217.400 ;
        RECT 146.415 217.400 154.000 217.700 ;
        RECT 146.415 217.375 146.765 217.400 ;
        RECT 153.620 217.390 154.000 217.400 ;
        RECT 69.135 217.200 69.485 217.225 ;
        RECT 72.020 217.200 72.340 217.240 ;
        RECT 55.335 217.075 55.685 217.100 ;
        RECT 69.135 216.900 72.340 217.200 ;
        RECT 69.135 216.875 69.485 216.900 ;
        RECT 72.020 216.860 72.340 216.900 ;
        RECT 45.215 215.725 45.565 216.075 ;
        RECT 27.750 213.465 29.330 213.795 ;
        RECT 62.595 213.465 64.175 213.795 ;
        RECT 97.440 213.465 99.020 213.795 ;
        RECT 132.285 213.465 133.865 213.795 ;
        RECT 45.170 210.745 46.750 211.075 ;
        RECT 80.015 210.745 81.595 211.075 ;
        RECT 114.860 210.745 116.440 211.075 ;
        RECT 149.705 210.745 151.285 211.075 ;
        RECT 27.750 208.025 29.330 208.355 ;
        RECT 62.595 208.025 64.175 208.355 ;
        RECT 97.440 208.025 99.020 208.355 ;
        RECT 132.285 208.025 133.865 208.355 ;
        RECT 45.170 205.305 46.750 205.635 ;
        RECT 80.015 205.305 81.595 205.635 ;
        RECT 114.860 205.305 116.440 205.635 ;
        RECT 149.705 205.305 151.285 205.635 ;
        RECT 27.750 202.585 29.330 202.915 ;
        RECT 62.595 202.585 64.175 202.915 ;
        RECT 97.440 202.585 99.020 202.915 ;
        RECT 132.285 202.585 133.865 202.915 ;
        RECT 45.170 199.865 46.750 200.195 ;
        RECT 80.015 199.865 81.595 200.195 ;
        RECT 114.860 199.865 116.440 200.195 ;
        RECT 149.705 199.865 151.285 200.195 ;
        RECT 76.965 199.160 77.295 199.175 ;
        RECT 101.345 199.160 101.675 199.175 ;
        RECT 76.965 198.860 101.675 199.160 ;
        RECT 76.965 198.845 77.295 198.860 ;
        RECT 101.345 198.845 101.675 198.860 ;
        RECT 27.750 197.145 29.330 197.475 ;
        RECT 62.595 197.145 64.175 197.475 ;
        RECT 97.440 197.145 99.020 197.475 ;
        RECT 132.285 197.145 133.865 197.475 ;
        RECT 45.170 194.425 46.750 194.755 ;
        RECT 80.015 194.425 81.595 194.755 ;
        RECT 114.860 194.425 116.440 194.755 ;
        RECT 149.705 194.425 151.285 194.755 ;
        RECT 27.750 191.705 29.330 192.035 ;
        RECT 62.595 191.705 64.175 192.035 ;
        RECT 97.440 191.705 99.020 192.035 ;
        RECT 132.285 191.705 133.865 192.035 ;
        RECT 45.170 188.985 46.750 189.315 ;
        RECT 80.015 188.985 81.595 189.315 ;
        RECT 114.860 188.985 116.440 189.315 ;
        RECT 149.705 188.985 151.285 189.315 ;
        RECT 83.405 188.280 83.735 188.295 ;
        RECT 122.965 188.280 123.295 188.295 ;
        RECT 83.405 187.980 123.295 188.280 ;
        RECT 83.405 187.965 83.735 187.980 ;
        RECT 122.965 187.965 123.295 187.980 ;
        RECT 19.465 187.600 19.795 187.615 ;
        RECT 74.205 187.600 74.535 187.615 ;
        RECT 19.465 187.300 74.535 187.600 ;
        RECT 19.465 187.285 19.795 187.300 ;
        RECT 74.205 187.285 74.535 187.300 ;
        RECT 76.965 187.600 77.295 187.615 ;
        RECT 94.905 187.600 95.235 187.615 ;
        RECT 102.265 187.600 102.595 187.615 ;
        RECT 76.965 187.300 95.235 187.600 ;
        RECT 76.965 187.285 77.295 187.300 ;
        RECT 94.905 187.285 95.235 187.300 ;
        RECT 96.070 187.300 102.595 187.600 ;
        RECT 70.065 186.920 70.395 186.935 ;
        RECT 87.545 186.920 87.875 186.935 ;
        RECT 96.070 186.920 96.370 187.300 ;
        RECT 102.265 187.285 102.595 187.300 ;
        RECT 70.065 186.620 96.370 186.920 ;
        RECT 70.065 186.605 70.395 186.620 ;
        RECT 87.545 186.605 87.875 186.620 ;
        RECT 27.750 186.265 29.330 186.595 ;
        RECT 62.595 186.265 64.175 186.595 ;
        RECT 97.440 186.265 99.020 186.595 ;
        RECT 132.285 186.265 133.865 186.595 ;
        RECT 30.045 184.880 30.375 184.895 ;
        RECT 35.105 184.880 35.435 184.895 ;
        RECT 30.045 184.580 35.435 184.880 ;
        RECT 30.045 184.565 30.375 184.580 ;
        RECT 35.105 184.565 35.435 184.580 ;
        RECT 45.170 183.545 46.750 183.875 ;
        RECT 80.015 183.545 81.595 183.875 ;
        RECT 114.860 183.545 116.440 183.875 ;
        RECT 149.705 183.545 151.285 183.875 ;
        RECT 113.765 182.840 114.095 182.855 ;
        RECT 125.725 182.840 126.055 182.855 ;
        RECT 113.765 182.540 126.055 182.840 ;
        RECT 113.765 182.525 114.095 182.540 ;
        RECT 125.725 182.525 126.055 182.540 ;
        RECT 47.065 182.160 47.395 182.175 ;
        RECT 76.965 182.160 77.295 182.175 ;
        RECT 47.065 181.860 77.295 182.160 ;
        RECT 47.065 181.845 47.395 181.860 ;
        RECT 76.965 181.845 77.295 181.860 ;
        RECT 27.750 180.825 29.330 181.155 ;
        RECT 62.595 180.825 64.175 181.155 ;
        RECT 97.440 180.825 99.020 181.155 ;
        RECT 132.285 180.825 133.865 181.155 ;
        RECT 66.385 179.440 66.715 179.455 ;
        RECT 67.765 179.440 68.095 179.455 ;
        RECT 92.145 179.440 92.475 179.455 ;
        RECT 66.385 179.140 92.475 179.440 ;
        RECT 66.385 179.125 66.715 179.140 ;
        RECT 67.765 179.125 68.095 179.140 ;
        RECT 92.145 179.125 92.475 179.140 ;
        RECT 45.170 178.105 46.750 178.435 ;
        RECT 80.015 178.105 81.595 178.435 ;
        RECT 114.860 178.105 116.440 178.435 ;
        RECT 149.705 178.105 151.285 178.435 ;
        RECT 57.645 176.720 57.975 176.735 ;
        RECT 57.645 176.420 70.610 176.720 ;
        RECT 57.645 176.405 57.975 176.420 ;
        RECT 70.310 176.040 70.610 176.420 ;
        RECT 75.790 176.040 76.170 176.050 ;
        RECT 78.805 176.040 79.135 176.055 ;
        RECT 70.310 175.740 79.135 176.040 ;
        RECT 75.790 175.730 76.170 175.740 ;
        RECT 78.805 175.725 79.135 175.740 ;
        RECT 27.750 175.385 29.330 175.715 ;
        RECT 62.595 175.385 64.175 175.715 ;
        RECT 97.440 175.385 99.020 175.715 ;
        RECT 132.285 175.385 133.865 175.715 ;
        RECT 36.945 174.680 37.275 174.695 ;
        RECT 63.625 174.680 63.955 174.695 ;
        RECT 36.945 174.380 63.955 174.680 ;
        RECT 36.945 174.365 37.275 174.380 ;
        RECT 63.625 174.365 63.955 174.380 ;
        RECT 45.170 172.665 46.750 172.995 ;
        RECT 80.015 172.665 81.595 172.995 ;
        RECT 114.860 172.665 116.440 172.995 ;
        RECT 149.705 172.665 151.285 172.995 ;
        RECT 27.750 169.945 29.330 170.275 ;
        RECT 62.595 169.945 64.175 170.275 ;
        RECT 97.440 169.945 99.020 170.275 ;
        RECT 132.285 169.945 133.865 170.275 ;
        RECT 26.365 169.240 26.695 169.255 ;
        RECT 39.245 169.240 39.575 169.255 ;
        RECT 26.365 168.940 39.575 169.240 ;
        RECT 26.365 168.925 26.695 168.940 ;
        RECT 39.245 168.925 39.575 168.940 ;
        RECT 116.065 168.560 116.395 168.575 ;
        RECT 146.425 168.560 146.755 168.575 ;
        RECT 116.065 168.260 146.755 168.560 ;
        RECT 116.065 168.245 116.395 168.260 ;
        RECT 146.425 168.245 146.755 168.260 ;
        RECT 45.170 167.225 46.750 167.555 ;
        RECT 80.015 167.225 81.595 167.555 ;
        RECT 114.860 167.225 116.440 167.555 ;
        RECT 149.705 167.225 151.285 167.555 ;
        RECT 27.750 164.505 29.330 164.835 ;
        RECT 62.595 164.505 64.175 164.835 ;
        RECT 97.440 164.505 99.020 164.835 ;
        RECT 132.285 164.505 133.865 164.835 ;
        RECT 45.170 161.785 46.750 162.115 ;
        RECT 80.015 161.785 81.595 162.115 ;
        RECT 114.860 161.785 116.440 162.115 ;
        RECT 149.705 161.785 151.285 162.115 ;
        RECT 75.125 160.400 75.455 160.415 ;
        RECT 81.565 160.400 81.895 160.415 ;
        RECT 75.125 160.100 81.895 160.400 ;
        RECT 75.125 160.085 75.455 160.100 ;
        RECT 81.565 160.085 81.895 160.100 ;
        RECT 27.750 159.065 29.330 159.395 ;
        RECT 62.595 159.065 64.175 159.395 ;
        RECT 97.440 159.065 99.020 159.395 ;
        RECT 132.285 159.065 133.865 159.395 ;
        RECT 73.285 157.680 73.615 157.695 ;
        RECT 92.605 157.680 92.935 157.695 ;
        RECT 73.285 157.380 92.935 157.680 ;
        RECT 73.285 157.365 73.615 157.380 ;
        RECT 92.605 157.365 92.935 157.380 ;
        RECT 45.170 156.345 46.750 156.675 ;
        RECT 80.015 156.345 81.595 156.675 ;
        RECT 114.860 156.345 116.440 156.675 ;
        RECT 149.705 156.345 151.285 156.675 ;
        RECT 75.585 154.290 75.915 154.295 ;
        RECT 75.585 154.280 76.170 154.290 ;
        RECT 75.585 153.980 76.370 154.280 ;
        RECT 75.585 153.970 76.170 153.980 ;
        RECT 75.585 153.965 75.915 153.970 ;
        RECT 27.750 153.625 29.330 153.955 ;
        RECT 62.595 153.625 64.175 153.955 ;
        RECT 97.440 153.625 99.020 153.955 ;
        RECT 132.285 153.625 133.865 153.955 ;
        RECT 87.085 152.920 87.415 152.935 ;
        RECT 97.205 152.920 97.535 152.935 ;
        RECT 87.085 152.620 97.535 152.920 ;
        RECT 87.085 152.605 87.415 152.620 ;
        RECT 97.205 152.605 97.535 152.620 ;
        RECT 88.005 152.240 88.335 152.255 ;
        RECT 97.665 152.240 97.995 152.255 ;
        RECT 88.005 151.940 97.995 152.240 ;
        RECT 88.005 151.925 88.335 151.940 ;
        RECT 97.665 151.925 97.995 151.940 ;
        RECT 45.170 150.905 46.750 151.235 ;
        RECT 80.015 150.905 81.595 151.235 ;
        RECT 114.860 150.905 116.440 151.235 ;
        RECT 149.705 150.905 151.285 151.235 ;
        RECT 27.750 148.185 29.330 148.515 ;
        RECT 62.595 148.185 64.175 148.515 ;
        RECT 97.440 148.185 99.020 148.515 ;
        RECT 132.285 148.185 133.865 148.515 ;
        RECT 59.945 146.800 60.275 146.815 ;
        RECT 66.845 146.800 67.175 146.815 ;
        RECT 59.945 146.500 67.175 146.800 ;
        RECT 59.945 146.485 60.275 146.500 ;
        RECT 66.845 146.485 67.175 146.500 ;
        RECT 45.170 145.465 46.750 145.795 ;
        RECT 80.015 145.465 81.595 145.795 ;
        RECT 114.860 145.465 116.440 145.795 ;
        RECT 149.705 145.465 151.285 145.795 ;
        RECT 27.750 142.745 29.330 143.075 ;
        RECT 62.595 142.745 64.175 143.075 ;
        RECT 97.440 142.745 99.020 143.075 ;
        RECT 132.285 142.745 133.865 143.075 ;
        RECT 45.170 140.025 46.750 140.355 ;
        RECT 80.015 140.025 81.595 140.355 ;
        RECT 114.860 140.025 116.440 140.355 ;
        RECT 149.705 140.025 151.285 140.355 ;
        RECT 27.750 137.305 29.330 137.635 ;
        RECT 62.595 137.305 64.175 137.635 ;
        RECT 97.440 137.305 99.020 137.635 ;
        RECT 132.285 137.305 133.865 137.635 ;
        RECT 75.585 136.600 75.915 136.615 ;
        RECT 89.845 136.600 90.175 136.615 ;
        RECT 75.585 136.300 90.175 136.600 ;
        RECT 75.585 136.285 75.915 136.300 ;
        RECT 89.845 136.285 90.175 136.300 ;
        RECT 77.885 135.920 78.215 135.935 ;
        RECT 77.885 135.620 83.490 135.920 ;
        RECT 77.885 135.605 78.215 135.620 ;
        RECT 83.190 135.255 83.490 135.620 ;
        RECT 83.190 134.940 83.735 135.255 ;
        RECT 83.405 134.925 83.735 134.940 ;
        RECT 45.170 134.585 46.750 134.915 ;
        RECT 80.015 134.585 81.595 134.915 ;
        RECT 114.860 134.585 116.440 134.915 ;
        RECT 149.705 134.585 151.285 134.915 ;
        RECT 27.750 131.865 29.330 132.195 ;
        RECT 62.595 131.865 64.175 132.195 ;
        RECT 97.440 131.865 99.020 132.195 ;
        RECT 132.285 131.865 133.865 132.195 ;
        RECT 45.170 129.145 46.750 129.475 ;
        RECT 80.015 129.145 81.595 129.475 ;
        RECT 114.860 129.145 116.440 129.475 ;
        RECT 149.705 129.145 151.285 129.475 ;
        RECT 27.750 126.425 29.330 126.755 ;
        RECT 62.595 126.425 64.175 126.755 ;
        RECT 97.440 126.425 99.020 126.755 ;
        RECT 132.285 126.425 133.865 126.755 ;
        RECT 45.170 123.705 46.750 124.035 ;
        RECT 80.015 123.705 81.595 124.035 ;
        RECT 114.860 123.705 116.440 124.035 ;
        RECT 149.705 123.705 151.285 124.035 ;
        RECT 27.750 120.985 29.330 121.315 ;
        RECT 62.595 120.985 64.175 121.315 ;
        RECT 97.440 120.985 99.020 121.315 ;
        RECT 132.285 120.985 133.865 121.315 ;
        RECT 45.170 118.265 46.750 118.595 ;
        RECT 80.015 118.265 81.595 118.595 ;
        RECT 114.860 118.265 116.440 118.595 ;
        RECT 149.705 118.265 151.285 118.595 ;
        RECT 27.750 115.545 29.330 115.875 ;
        RECT 62.595 115.545 64.175 115.875 ;
        RECT 97.440 115.545 99.020 115.875 ;
        RECT 132.285 115.545 133.865 115.875 ;
        RECT 45.170 112.825 46.750 113.155 ;
        RECT 80.015 112.825 81.595 113.155 ;
        RECT 114.860 112.825 116.440 113.155 ;
        RECT 149.705 112.825 151.285 113.155 ;
        RECT 27.750 110.105 29.330 110.435 ;
        RECT 62.595 110.105 64.175 110.435 ;
        RECT 97.440 110.105 99.020 110.435 ;
        RECT 132.285 110.105 133.865 110.435 ;
        RECT 45.170 107.385 46.750 107.715 ;
        RECT 80.015 107.385 81.595 107.715 ;
        RECT 114.860 107.385 116.440 107.715 ;
        RECT 149.705 107.385 151.285 107.715 ;
        RECT 27.750 104.665 29.330 104.995 ;
        RECT 62.595 104.665 64.175 104.995 ;
        RECT 97.440 104.665 99.020 104.995 ;
        RECT 132.285 104.665 133.865 104.995 ;
        RECT 45.170 101.945 46.750 102.275 ;
        RECT 80.015 101.945 81.595 102.275 ;
        RECT 114.860 101.945 116.440 102.275 ;
        RECT 149.705 101.945 151.285 102.275 ;
        RECT 27.750 99.225 29.330 99.555 ;
        RECT 62.595 99.225 64.175 99.555 ;
        RECT 97.440 99.225 99.020 99.555 ;
        RECT 132.285 99.225 133.865 99.555 ;
        RECT 45.170 96.505 46.750 96.835 ;
        RECT 80.015 96.505 81.595 96.835 ;
        RECT 114.860 96.505 116.440 96.835 ;
        RECT 149.705 96.505 151.285 96.835 ;
        RECT 27.750 93.785 29.330 94.115 ;
        RECT 62.595 93.785 64.175 94.115 ;
        RECT 97.440 93.785 99.020 94.115 ;
        RECT 132.285 93.785 133.865 94.115 ;
        RECT 45.170 91.065 46.750 91.395 ;
        RECT 80.015 91.065 81.595 91.395 ;
        RECT 114.860 91.065 116.440 91.395 ;
        RECT 149.705 91.065 151.285 91.395 ;
        RECT 27.750 88.345 29.330 88.675 ;
        RECT 62.595 88.345 64.175 88.675 ;
        RECT 97.440 88.345 99.020 88.675 ;
        RECT 132.285 88.345 133.865 88.675 ;
        RECT 45.170 85.625 46.750 85.955 ;
        RECT 80.015 85.625 81.595 85.955 ;
        RECT 114.860 85.625 116.440 85.955 ;
        RECT 149.705 85.625 151.285 85.955 ;
        RECT 27.750 82.905 29.330 83.235 ;
        RECT 62.595 82.905 64.175 83.235 ;
        RECT 97.440 82.905 99.020 83.235 ;
        RECT 132.285 82.905 133.865 83.235 ;
        RECT 45.170 80.185 46.750 80.515 ;
        RECT 80.015 80.185 81.595 80.515 ;
        RECT 114.860 80.185 116.440 80.515 ;
        RECT 149.705 80.185 151.285 80.515 ;
        RECT 27.750 77.465 29.330 77.795 ;
        RECT 62.595 77.465 64.175 77.795 ;
        RECT 97.440 77.465 99.020 77.795 ;
        RECT 132.285 77.465 133.865 77.795 ;
        RECT 45.170 74.745 46.750 75.075 ;
        RECT 80.015 74.745 81.595 75.075 ;
        RECT 114.860 74.745 116.440 75.075 ;
        RECT 149.705 74.745 151.285 75.075 ;
        RECT 27.700 74.270 29.260 74.280 ;
        RECT 27.630 72.680 29.350 74.270 ;
        RECT 62.530 72.680 64.210 74.400 ;
        RECT 97.390 74.300 98.950 74.340 ;
        RECT 27.700 63.130 29.260 72.680 ;
        RECT 27.700 60.870 53.830 63.130 ;
        RECT 62.640 63.080 64.200 72.680 ;
        RECT 97.340 72.580 99.000 74.300 ;
        RECT 132.320 74.030 133.880 74.060 ;
        RECT 62.550 61.130 64.230 63.080 ;
        RECT 97.390 63.040 98.950 72.580 ;
        RECT 132.320 72.560 133.930 74.030 ;
        RECT 62.640 61.110 64.200 61.130 ;
        RECT 97.320 61.090 99.000 63.040 ;
        RECT 132.320 62.770 133.880 72.560 ;
        RECT 97.390 61.050 98.950 61.090 ;
        RECT 132.170 60.770 134.390 62.770 ;
        RECT 54.930 54.700 77.070 59.620 ;
        RECT 95.020 50.660 105.690 60.270 ;
        RECT 117.160 54.670 134.820 58.500 ;
        RECT 62.020 49.675 62.960 49.850 ;
        RECT 64.680 49.725 65.580 50.260 ;
        RECT 61.950 49.265 62.990 49.675 ;
        RECT 64.630 49.275 65.640 49.725 ;
        RECT 78.760 49.665 79.770 49.670 ;
        RECT 62.020 45.035 62.960 49.265 ;
        RECT 64.680 45.055 65.580 49.275 ;
        RECT 78.710 49.135 79.800 49.665 ;
        RECT 124.250 49.275 125.190 49.450 ;
        RECT 126.910 49.325 127.810 49.860 ;
        RECT 78.760 48.085 79.770 49.135 ;
        RECT 124.180 48.865 125.220 49.275 ;
        RECT 126.860 48.875 127.870 49.325 ;
        RECT 140.990 49.265 142.000 49.270 ;
        RECT 78.700 47.555 79.790 48.085 ;
        RECT 78.760 46.515 79.770 47.555 ;
        RECT 78.690 45.985 79.780 46.515 ;
        RECT 61.950 44.625 62.990 45.035 ;
        RECT 62.020 40.465 62.960 44.625 ;
        RECT 64.630 44.605 65.640 45.055 ;
        RECT 78.760 44.925 79.770 45.985 ;
        RECT 64.680 40.485 65.580 44.605 ;
        RECT 78.720 44.395 79.810 44.925 ;
        RECT 124.250 44.635 125.190 48.865 ;
        RECT 126.910 44.655 127.810 48.875 ;
        RECT 140.940 48.735 142.030 49.265 ;
        RECT 140.990 47.685 142.000 48.735 ;
        RECT 140.930 47.155 142.020 47.685 ;
        RECT 140.990 46.115 142.000 47.155 ;
        RECT 140.920 45.585 142.010 46.115 ;
        RECT 78.760 43.345 79.770 44.395 ;
        RECT 124.180 44.225 125.220 44.635 ;
        RECT 78.720 42.815 79.810 43.345 ;
        RECT 78.760 41.765 79.770 42.815 ;
        RECT 78.720 41.235 79.810 41.765 ;
        RECT 61.960 40.055 63.000 40.465 ;
        RECT 62.020 35.865 62.960 40.055 ;
        RECT 64.620 40.035 65.630 40.485 ;
        RECT 64.680 35.865 65.580 40.035 ;
        RECT 61.980 35.515 62.990 35.865 ;
        RECT 64.640 35.465 65.640 35.865 ;
        RECT 64.680 35.440 65.580 35.465 ;
        RECT 73.500 25.770 74.620 40.290 ;
        RECT 78.760 40.185 79.770 41.235 ;
        RECT 78.700 39.655 79.790 40.185 ;
        RECT 124.250 40.065 125.190 44.225 ;
        RECT 126.860 44.205 127.870 44.655 ;
        RECT 140.990 44.525 142.000 45.585 ;
        RECT 126.910 40.085 127.810 44.205 ;
        RECT 140.950 43.995 142.040 44.525 ;
        RECT 140.990 42.945 142.000 43.995 ;
        RECT 140.950 42.415 142.040 42.945 ;
        RECT 140.990 41.365 142.000 42.415 ;
        RECT 140.950 40.835 142.040 41.365 ;
        RECT 124.190 39.655 125.230 40.065 ;
        RECT 78.760 38.605 79.770 39.655 ;
        RECT 78.710 38.075 79.800 38.605 ;
        RECT 78.760 37.025 79.770 38.075 ;
        RECT 78.720 36.495 79.810 37.025 ;
        RECT 78.760 35.455 79.770 36.495 ;
        RECT 124.250 35.465 125.190 39.655 ;
        RECT 126.850 39.635 127.860 40.085 ;
        RECT 126.910 35.465 127.810 39.635 ;
        RECT 78.720 34.925 79.810 35.455 ;
        RECT 124.210 35.115 125.220 35.465 ;
        RECT 126.870 35.065 127.870 35.465 ;
        RECT 126.910 35.040 127.810 35.065 ;
        RECT 78.760 33.825 79.770 34.925 ;
        RECT 78.710 33.320 79.770 33.825 ;
        RECT 78.710 33.205 79.750 33.320 ;
        RECT 87.245 25.565 108.095 26.435 ;
        RECT 59.990 21.815 60.910 21.840 ;
        RECT 87.245 21.815 88.115 25.565 ;
        RECT 135.730 25.370 136.850 39.890 ;
        RECT 140.990 39.785 142.000 40.835 ;
        RECT 140.930 39.255 142.020 39.785 ;
        RECT 140.990 38.205 142.000 39.255 ;
        RECT 140.940 37.675 142.030 38.205 ;
        RECT 140.990 36.625 142.000 37.675 ;
        RECT 140.950 36.095 142.040 36.625 ;
        RECT 140.990 35.055 142.000 36.095 ;
        RECT 140.950 34.525 142.040 35.055 ;
        RECT 140.990 33.425 142.000 34.525 ;
        RECT 140.940 32.920 142.000 33.425 ;
        RECT 140.940 32.805 141.980 32.920 ;
        RECT 59.990 20.945 88.115 21.815 ;
        RECT 59.990 20.920 60.910 20.945 ;
        RECT 55.150 10.850 64.860 18.920 ;
        RECT 73.660 10.790 84.410 18.850 ;
        RECT 68.240 7.400 70.050 8.000 ;
        RECT 46.165 5.380 46.755 5.405 ;
        RECT 46.160 4.780 57.010 5.380 ;
        RECT 46.165 4.755 46.755 4.780 ;
        RECT 68.240 2.835 68.840 7.400 ;
        RECT 90.320 2.925 90.920 23.730 ;
        RECT 94.350 11.450 105.980 18.660 ;
        RECT 117.190 13.030 127.820 18.860 ;
        RECT 112.400 6.590 129.570 7.190 ;
        RECT 112.400 3.135 113.000 6.590 ;
        RECT 134.480 3.365 135.080 20.610 ;
        RECT 135.840 13.390 146.360 18.670 ;
        RECT 150.530 4.705 151.130 20.760 ;
        RECT 150.505 4.115 151.155 4.705 ;
        RECT 150.530 4.110 151.130 4.115 ;
        RECT 68.215 2.245 68.865 2.835 ;
        RECT 90.295 2.335 90.945 2.925 ;
        RECT 112.375 2.545 113.025 3.135 ;
        RECT 134.455 2.775 135.105 3.365 ;
        RECT 150.530 3.065 151.130 3.100 ;
        RECT 134.480 2.770 135.080 2.775 ;
        RECT 112.400 2.540 113.000 2.545 ;
        RECT 150.505 2.475 151.155 3.065 ;
        RECT 150.530 2.440 151.130 2.475 ;
        RECT 90.320 2.330 90.920 2.335 ;
        RECT 68.240 2.240 68.840 2.245 ;
      LAYER via3 ;
        RECT 60.020 223.410 60.340 223.730 ;
        RECT 74.980 223.580 75.300 223.900 ;
        RECT 24.990 218.510 25.310 218.830 ;
        RECT 70.220 221.550 70.540 221.870 ;
        RECT 73.870 221.510 74.190 221.830 ;
        RECT 129.560 223.580 129.880 223.900 ;
        RECT 143.800 222.490 144.120 222.810 ;
        RECT 151.180 222.270 151.500 222.590 ;
        RECT 105.950 219.840 106.270 220.160 ;
        RECT 87.180 218.440 87.500 218.760 ;
        RECT 126.190 219.260 126.510 219.580 ;
        RECT 83.810 217.730 84.130 218.050 ;
        RECT 153.650 217.390 153.970 217.710 ;
        RECT 72.020 216.890 72.340 217.210 ;
        RECT 27.780 213.470 28.100 213.790 ;
        RECT 28.180 213.470 28.500 213.790 ;
        RECT 28.580 213.470 28.900 213.790 ;
        RECT 28.980 213.470 29.300 213.790 ;
        RECT 62.625 213.470 62.945 213.790 ;
        RECT 63.025 213.470 63.345 213.790 ;
        RECT 63.425 213.470 63.745 213.790 ;
        RECT 63.825 213.470 64.145 213.790 ;
        RECT 97.470 213.470 97.790 213.790 ;
        RECT 97.870 213.470 98.190 213.790 ;
        RECT 98.270 213.470 98.590 213.790 ;
        RECT 98.670 213.470 98.990 213.790 ;
        RECT 132.315 213.470 132.635 213.790 ;
        RECT 132.715 213.470 133.035 213.790 ;
        RECT 133.115 213.470 133.435 213.790 ;
        RECT 133.515 213.470 133.835 213.790 ;
        RECT 45.200 210.750 45.520 211.070 ;
        RECT 45.600 210.750 45.920 211.070 ;
        RECT 46.000 210.750 46.320 211.070 ;
        RECT 46.400 210.750 46.720 211.070 ;
        RECT 80.045 210.750 80.365 211.070 ;
        RECT 80.445 210.750 80.765 211.070 ;
        RECT 80.845 210.750 81.165 211.070 ;
        RECT 81.245 210.750 81.565 211.070 ;
        RECT 114.890 210.750 115.210 211.070 ;
        RECT 115.290 210.750 115.610 211.070 ;
        RECT 115.690 210.750 116.010 211.070 ;
        RECT 116.090 210.750 116.410 211.070 ;
        RECT 149.735 210.750 150.055 211.070 ;
        RECT 150.135 210.750 150.455 211.070 ;
        RECT 150.535 210.750 150.855 211.070 ;
        RECT 150.935 210.750 151.255 211.070 ;
        RECT 27.780 208.030 28.100 208.350 ;
        RECT 28.180 208.030 28.500 208.350 ;
        RECT 28.580 208.030 28.900 208.350 ;
        RECT 28.980 208.030 29.300 208.350 ;
        RECT 62.625 208.030 62.945 208.350 ;
        RECT 63.025 208.030 63.345 208.350 ;
        RECT 63.425 208.030 63.745 208.350 ;
        RECT 63.825 208.030 64.145 208.350 ;
        RECT 97.470 208.030 97.790 208.350 ;
        RECT 97.870 208.030 98.190 208.350 ;
        RECT 98.270 208.030 98.590 208.350 ;
        RECT 98.670 208.030 98.990 208.350 ;
        RECT 132.315 208.030 132.635 208.350 ;
        RECT 132.715 208.030 133.035 208.350 ;
        RECT 133.115 208.030 133.435 208.350 ;
        RECT 133.515 208.030 133.835 208.350 ;
        RECT 45.200 205.310 45.520 205.630 ;
        RECT 45.600 205.310 45.920 205.630 ;
        RECT 46.000 205.310 46.320 205.630 ;
        RECT 46.400 205.310 46.720 205.630 ;
        RECT 80.045 205.310 80.365 205.630 ;
        RECT 80.445 205.310 80.765 205.630 ;
        RECT 80.845 205.310 81.165 205.630 ;
        RECT 81.245 205.310 81.565 205.630 ;
        RECT 114.890 205.310 115.210 205.630 ;
        RECT 115.290 205.310 115.610 205.630 ;
        RECT 115.690 205.310 116.010 205.630 ;
        RECT 116.090 205.310 116.410 205.630 ;
        RECT 149.735 205.310 150.055 205.630 ;
        RECT 150.135 205.310 150.455 205.630 ;
        RECT 150.535 205.310 150.855 205.630 ;
        RECT 150.935 205.310 151.255 205.630 ;
        RECT 27.780 202.590 28.100 202.910 ;
        RECT 28.180 202.590 28.500 202.910 ;
        RECT 28.580 202.590 28.900 202.910 ;
        RECT 28.980 202.590 29.300 202.910 ;
        RECT 62.625 202.590 62.945 202.910 ;
        RECT 63.025 202.590 63.345 202.910 ;
        RECT 63.425 202.590 63.745 202.910 ;
        RECT 63.825 202.590 64.145 202.910 ;
        RECT 97.470 202.590 97.790 202.910 ;
        RECT 97.870 202.590 98.190 202.910 ;
        RECT 98.270 202.590 98.590 202.910 ;
        RECT 98.670 202.590 98.990 202.910 ;
        RECT 132.315 202.590 132.635 202.910 ;
        RECT 132.715 202.590 133.035 202.910 ;
        RECT 133.115 202.590 133.435 202.910 ;
        RECT 133.515 202.590 133.835 202.910 ;
        RECT 45.200 199.870 45.520 200.190 ;
        RECT 45.600 199.870 45.920 200.190 ;
        RECT 46.000 199.870 46.320 200.190 ;
        RECT 46.400 199.870 46.720 200.190 ;
        RECT 80.045 199.870 80.365 200.190 ;
        RECT 80.445 199.870 80.765 200.190 ;
        RECT 80.845 199.870 81.165 200.190 ;
        RECT 81.245 199.870 81.565 200.190 ;
        RECT 114.890 199.870 115.210 200.190 ;
        RECT 115.290 199.870 115.610 200.190 ;
        RECT 115.690 199.870 116.010 200.190 ;
        RECT 116.090 199.870 116.410 200.190 ;
        RECT 149.735 199.870 150.055 200.190 ;
        RECT 150.135 199.870 150.455 200.190 ;
        RECT 150.535 199.870 150.855 200.190 ;
        RECT 150.935 199.870 151.255 200.190 ;
        RECT 27.780 197.150 28.100 197.470 ;
        RECT 28.180 197.150 28.500 197.470 ;
        RECT 28.580 197.150 28.900 197.470 ;
        RECT 28.980 197.150 29.300 197.470 ;
        RECT 62.625 197.150 62.945 197.470 ;
        RECT 63.025 197.150 63.345 197.470 ;
        RECT 63.425 197.150 63.745 197.470 ;
        RECT 63.825 197.150 64.145 197.470 ;
        RECT 97.470 197.150 97.790 197.470 ;
        RECT 97.870 197.150 98.190 197.470 ;
        RECT 98.270 197.150 98.590 197.470 ;
        RECT 98.670 197.150 98.990 197.470 ;
        RECT 132.315 197.150 132.635 197.470 ;
        RECT 132.715 197.150 133.035 197.470 ;
        RECT 133.115 197.150 133.435 197.470 ;
        RECT 133.515 197.150 133.835 197.470 ;
        RECT 45.200 194.430 45.520 194.750 ;
        RECT 45.600 194.430 45.920 194.750 ;
        RECT 46.000 194.430 46.320 194.750 ;
        RECT 46.400 194.430 46.720 194.750 ;
        RECT 80.045 194.430 80.365 194.750 ;
        RECT 80.445 194.430 80.765 194.750 ;
        RECT 80.845 194.430 81.165 194.750 ;
        RECT 81.245 194.430 81.565 194.750 ;
        RECT 114.890 194.430 115.210 194.750 ;
        RECT 115.290 194.430 115.610 194.750 ;
        RECT 115.690 194.430 116.010 194.750 ;
        RECT 116.090 194.430 116.410 194.750 ;
        RECT 149.735 194.430 150.055 194.750 ;
        RECT 150.135 194.430 150.455 194.750 ;
        RECT 150.535 194.430 150.855 194.750 ;
        RECT 150.935 194.430 151.255 194.750 ;
        RECT 27.780 191.710 28.100 192.030 ;
        RECT 28.180 191.710 28.500 192.030 ;
        RECT 28.580 191.710 28.900 192.030 ;
        RECT 28.980 191.710 29.300 192.030 ;
        RECT 62.625 191.710 62.945 192.030 ;
        RECT 63.025 191.710 63.345 192.030 ;
        RECT 63.425 191.710 63.745 192.030 ;
        RECT 63.825 191.710 64.145 192.030 ;
        RECT 97.470 191.710 97.790 192.030 ;
        RECT 97.870 191.710 98.190 192.030 ;
        RECT 98.270 191.710 98.590 192.030 ;
        RECT 98.670 191.710 98.990 192.030 ;
        RECT 132.315 191.710 132.635 192.030 ;
        RECT 132.715 191.710 133.035 192.030 ;
        RECT 133.115 191.710 133.435 192.030 ;
        RECT 133.515 191.710 133.835 192.030 ;
        RECT 45.200 188.990 45.520 189.310 ;
        RECT 45.600 188.990 45.920 189.310 ;
        RECT 46.000 188.990 46.320 189.310 ;
        RECT 46.400 188.990 46.720 189.310 ;
        RECT 80.045 188.990 80.365 189.310 ;
        RECT 80.445 188.990 80.765 189.310 ;
        RECT 80.845 188.990 81.165 189.310 ;
        RECT 81.245 188.990 81.565 189.310 ;
        RECT 114.890 188.990 115.210 189.310 ;
        RECT 115.290 188.990 115.610 189.310 ;
        RECT 115.690 188.990 116.010 189.310 ;
        RECT 116.090 188.990 116.410 189.310 ;
        RECT 149.735 188.990 150.055 189.310 ;
        RECT 150.135 188.990 150.455 189.310 ;
        RECT 150.535 188.990 150.855 189.310 ;
        RECT 150.935 188.990 151.255 189.310 ;
        RECT 27.780 186.270 28.100 186.590 ;
        RECT 28.180 186.270 28.500 186.590 ;
        RECT 28.580 186.270 28.900 186.590 ;
        RECT 28.980 186.270 29.300 186.590 ;
        RECT 62.625 186.270 62.945 186.590 ;
        RECT 63.025 186.270 63.345 186.590 ;
        RECT 63.425 186.270 63.745 186.590 ;
        RECT 63.825 186.270 64.145 186.590 ;
        RECT 97.470 186.270 97.790 186.590 ;
        RECT 97.870 186.270 98.190 186.590 ;
        RECT 98.270 186.270 98.590 186.590 ;
        RECT 98.670 186.270 98.990 186.590 ;
        RECT 132.315 186.270 132.635 186.590 ;
        RECT 132.715 186.270 133.035 186.590 ;
        RECT 133.115 186.270 133.435 186.590 ;
        RECT 133.515 186.270 133.835 186.590 ;
        RECT 45.200 183.550 45.520 183.870 ;
        RECT 45.600 183.550 45.920 183.870 ;
        RECT 46.000 183.550 46.320 183.870 ;
        RECT 46.400 183.550 46.720 183.870 ;
        RECT 80.045 183.550 80.365 183.870 ;
        RECT 80.445 183.550 80.765 183.870 ;
        RECT 80.845 183.550 81.165 183.870 ;
        RECT 81.245 183.550 81.565 183.870 ;
        RECT 114.890 183.550 115.210 183.870 ;
        RECT 115.290 183.550 115.610 183.870 ;
        RECT 115.690 183.550 116.010 183.870 ;
        RECT 116.090 183.550 116.410 183.870 ;
        RECT 149.735 183.550 150.055 183.870 ;
        RECT 150.135 183.550 150.455 183.870 ;
        RECT 150.535 183.550 150.855 183.870 ;
        RECT 150.935 183.550 151.255 183.870 ;
        RECT 27.780 180.830 28.100 181.150 ;
        RECT 28.180 180.830 28.500 181.150 ;
        RECT 28.580 180.830 28.900 181.150 ;
        RECT 28.980 180.830 29.300 181.150 ;
        RECT 62.625 180.830 62.945 181.150 ;
        RECT 63.025 180.830 63.345 181.150 ;
        RECT 63.425 180.830 63.745 181.150 ;
        RECT 63.825 180.830 64.145 181.150 ;
        RECT 97.470 180.830 97.790 181.150 ;
        RECT 97.870 180.830 98.190 181.150 ;
        RECT 98.270 180.830 98.590 181.150 ;
        RECT 98.670 180.830 98.990 181.150 ;
        RECT 132.315 180.830 132.635 181.150 ;
        RECT 132.715 180.830 133.035 181.150 ;
        RECT 133.115 180.830 133.435 181.150 ;
        RECT 133.515 180.830 133.835 181.150 ;
        RECT 45.200 178.110 45.520 178.430 ;
        RECT 45.600 178.110 45.920 178.430 ;
        RECT 46.000 178.110 46.320 178.430 ;
        RECT 46.400 178.110 46.720 178.430 ;
        RECT 80.045 178.110 80.365 178.430 ;
        RECT 80.445 178.110 80.765 178.430 ;
        RECT 80.845 178.110 81.165 178.430 ;
        RECT 81.245 178.110 81.565 178.430 ;
        RECT 114.890 178.110 115.210 178.430 ;
        RECT 115.290 178.110 115.610 178.430 ;
        RECT 115.690 178.110 116.010 178.430 ;
        RECT 116.090 178.110 116.410 178.430 ;
        RECT 149.735 178.110 150.055 178.430 ;
        RECT 150.135 178.110 150.455 178.430 ;
        RECT 150.535 178.110 150.855 178.430 ;
        RECT 150.935 178.110 151.255 178.430 ;
        RECT 75.820 175.730 76.140 176.050 ;
        RECT 27.780 175.390 28.100 175.710 ;
        RECT 28.180 175.390 28.500 175.710 ;
        RECT 28.580 175.390 28.900 175.710 ;
        RECT 28.980 175.390 29.300 175.710 ;
        RECT 62.625 175.390 62.945 175.710 ;
        RECT 63.025 175.390 63.345 175.710 ;
        RECT 63.425 175.390 63.745 175.710 ;
        RECT 63.825 175.390 64.145 175.710 ;
        RECT 97.470 175.390 97.790 175.710 ;
        RECT 97.870 175.390 98.190 175.710 ;
        RECT 98.270 175.390 98.590 175.710 ;
        RECT 98.670 175.390 98.990 175.710 ;
        RECT 132.315 175.390 132.635 175.710 ;
        RECT 132.715 175.390 133.035 175.710 ;
        RECT 133.115 175.390 133.435 175.710 ;
        RECT 133.515 175.390 133.835 175.710 ;
        RECT 45.200 172.670 45.520 172.990 ;
        RECT 45.600 172.670 45.920 172.990 ;
        RECT 46.000 172.670 46.320 172.990 ;
        RECT 46.400 172.670 46.720 172.990 ;
        RECT 80.045 172.670 80.365 172.990 ;
        RECT 80.445 172.670 80.765 172.990 ;
        RECT 80.845 172.670 81.165 172.990 ;
        RECT 81.245 172.670 81.565 172.990 ;
        RECT 114.890 172.670 115.210 172.990 ;
        RECT 115.290 172.670 115.610 172.990 ;
        RECT 115.690 172.670 116.010 172.990 ;
        RECT 116.090 172.670 116.410 172.990 ;
        RECT 149.735 172.670 150.055 172.990 ;
        RECT 150.135 172.670 150.455 172.990 ;
        RECT 150.535 172.670 150.855 172.990 ;
        RECT 150.935 172.670 151.255 172.990 ;
        RECT 27.780 169.950 28.100 170.270 ;
        RECT 28.180 169.950 28.500 170.270 ;
        RECT 28.580 169.950 28.900 170.270 ;
        RECT 28.980 169.950 29.300 170.270 ;
        RECT 62.625 169.950 62.945 170.270 ;
        RECT 63.025 169.950 63.345 170.270 ;
        RECT 63.425 169.950 63.745 170.270 ;
        RECT 63.825 169.950 64.145 170.270 ;
        RECT 97.470 169.950 97.790 170.270 ;
        RECT 97.870 169.950 98.190 170.270 ;
        RECT 98.270 169.950 98.590 170.270 ;
        RECT 98.670 169.950 98.990 170.270 ;
        RECT 132.315 169.950 132.635 170.270 ;
        RECT 132.715 169.950 133.035 170.270 ;
        RECT 133.115 169.950 133.435 170.270 ;
        RECT 133.515 169.950 133.835 170.270 ;
        RECT 45.200 167.230 45.520 167.550 ;
        RECT 45.600 167.230 45.920 167.550 ;
        RECT 46.000 167.230 46.320 167.550 ;
        RECT 46.400 167.230 46.720 167.550 ;
        RECT 80.045 167.230 80.365 167.550 ;
        RECT 80.445 167.230 80.765 167.550 ;
        RECT 80.845 167.230 81.165 167.550 ;
        RECT 81.245 167.230 81.565 167.550 ;
        RECT 114.890 167.230 115.210 167.550 ;
        RECT 115.290 167.230 115.610 167.550 ;
        RECT 115.690 167.230 116.010 167.550 ;
        RECT 116.090 167.230 116.410 167.550 ;
        RECT 149.735 167.230 150.055 167.550 ;
        RECT 150.135 167.230 150.455 167.550 ;
        RECT 150.535 167.230 150.855 167.550 ;
        RECT 150.935 167.230 151.255 167.550 ;
        RECT 27.780 164.510 28.100 164.830 ;
        RECT 28.180 164.510 28.500 164.830 ;
        RECT 28.580 164.510 28.900 164.830 ;
        RECT 28.980 164.510 29.300 164.830 ;
        RECT 62.625 164.510 62.945 164.830 ;
        RECT 63.025 164.510 63.345 164.830 ;
        RECT 63.425 164.510 63.745 164.830 ;
        RECT 63.825 164.510 64.145 164.830 ;
        RECT 97.470 164.510 97.790 164.830 ;
        RECT 97.870 164.510 98.190 164.830 ;
        RECT 98.270 164.510 98.590 164.830 ;
        RECT 98.670 164.510 98.990 164.830 ;
        RECT 132.315 164.510 132.635 164.830 ;
        RECT 132.715 164.510 133.035 164.830 ;
        RECT 133.115 164.510 133.435 164.830 ;
        RECT 133.515 164.510 133.835 164.830 ;
        RECT 45.200 161.790 45.520 162.110 ;
        RECT 45.600 161.790 45.920 162.110 ;
        RECT 46.000 161.790 46.320 162.110 ;
        RECT 46.400 161.790 46.720 162.110 ;
        RECT 80.045 161.790 80.365 162.110 ;
        RECT 80.445 161.790 80.765 162.110 ;
        RECT 80.845 161.790 81.165 162.110 ;
        RECT 81.245 161.790 81.565 162.110 ;
        RECT 114.890 161.790 115.210 162.110 ;
        RECT 115.290 161.790 115.610 162.110 ;
        RECT 115.690 161.790 116.010 162.110 ;
        RECT 116.090 161.790 116.410 162.110 ;
        RECT 149.735 161.790 150.055 162.110 ;
        RECT 150.135 161.790 150.455 162.110 ;
        RECT 150.535 161.790 150.855 162.110 ;
        RECT 150.935 161.790 151.255 162.110 ;
        RECT 27.780 159.070 28.100 159.390 ;
        RECT 28.180 159.070 28.500 159.390 ;
        RECT 28.580 159.070 28.900 159.390 ;
        RECT 28.980 159.070 29.300 159.390 ;
        RECT 62.625 159.070 62.945 159.390 ;
        RECT 63.025 159.070 63.345 159.390 ;
        RECT 63.425 159.070 63.745 159.390 ;
        RECT 63.825 159.070 64.145 159.390 ;
        RECT 97.470 159.070 97.790 159.390 ;
        RECT 97.870 159.070 98.190 159.390 ;
        RECT 98.270 159.070 98.590 159.390 ;
        RECT 98.670 159.070 98.990 159.390 ;
        RECT 132.315 159.070 132.635 159.390 ;
        RECT 132.715 159.070 133.035 159.390 ;
        RECT 133.115 159.070 133.435 159.390 ;
        RECT 133.515 159.070 133.835 159.390 ;
        RECT 45.200 156.350 45.520 156.670 ;
        RECT 45.600 156.350 45.920 156.670 ;
        RECT 46.000 156.350 46.320 156.670 ;
        RECT 46.400 156.350 46.720 156.670 ;
        RECT 80.045 156.350 80.365 156.670 ;
        RECT 80.445 156.350 80.765 156.670 ;
        RECT 80.845 156.350 81.165 156.670 ;
        RECT 81.245 156.350 81.565 156.670 ;
        RECT 114.890 156.350 115.210 156.670 ;
        RECT 115.290 156.350 115.610 156.670 ;
        RECT 115.690 156.350 116.010 156.670 ;
        RECT 116.090 156.350 116.410 156.670 ;
        RECT 149.735 156.350 150.055 156.670 ;
        RECT 150.135 156.350 150.455 156.670 ;
        RECT 150.535 156.350 150.855 156.670 ;
        RECT 150.935 156.350 151.255 156.670 ;
        RECT 75.820 153.970 76.140 154.290 ;
        RECT 27.780 153.630 28.100 153.950 ;
        RECT 28.180 153.630 28.500 153.950 ;
        RECT 28.580 153.630 28.900 153.950 ;
        RECT 28.980 153.630 29.300 153.950 ;
        RECT 62.625 153.630 62.945 153.950 ;
        RECT 63.025 153.630 63.345 153.950 ;
        RECT 63.425 153.630 63.745 153.950 ;
        RECT 63.825 153.630 64.145 153.950 ;
        RECT 97.470 153.630 97.790 153.950 ;
        RECT 97.870 153.630 98.190 153.950 ;
        RECT 98.270 153.630 98.590 153.950 ;
        RECT 98.670 153.630 98.990 153.950 ;
        RECT 132.315 153.630 132.635 153.950 ;
        RECT 132.715 153.630 133.035 153.950 ;
        RECT 133.115 153.630 133.435 153.950 ;
        RECT 133.515 153.630 133.835 153.950 ;
        RECT 45.200 150.910 45.520 151.230 ;
        RECT 45.600 150.910 45.920 151.230 ;
        RECT 46.000 150.910 46.320 151.230 ;
        RECT 46.400 150.910 46.720 151.230 ;
        RECT 80.045 150.910 80.365 151.230 ;
        RECT 80.445 150.910 80.765 151.230 ;
        RECT 80.845 150.910 81.165 151.230 ;
        RECT 81.245 150.910 81.565 151.230 ;
        RECT 114.890 150.910 115.210 151.230 ;
        RECT 115.290 150.910 115.610 151.230 ;
        RECT 115.690 150.910 116.010 151.230 ;
        RECT 116.090 150.910 116.410 151.230 ;
        RECT 149.735 150.910 150.055 151.230 ;
        RECT 150.135 150.910 150.455 151.230 ;
        RECT 150.535 150.910 150.855 151.230 ;
        RECT 150.935 150.910 151.255 151.230 ;
        RECT 27.780 148.190 28.100 148.510 ;
        RECT 28.180 148.190 28.500 148.510 ;
        RECT 28.580 148.190 28.900 148.510 ;
        RECT 28.980 148.190 29.300 148.510 ;
        RECT 62.625 148.190 62.945 148.510 ;
        RECT 63.025 148.190 63.345 148.510 ;
        RECT 63.425 148.190 63.745 148.510 ;
        RECT 63.825 148.190 64.145 148.510 ;
        RECT 97.470 148.190 97.790 148.510 ;
        RECT 97.870 148.190 98.190 148.510 ;
        RECT 98.270 148.190 98.590 148.510 ;
        RECT 98.670 148.190 98.990 148.510 ;
        RECT 132.315 148.190 132.635 148.510 ;
        RECT 132.715 148.190 133.035 148.510 ;
        RECT 133.115 148.190 133.435 148.510 ;
        RECT 133.515 148.190 133.835 148.510 ;
        RECT 45.200 145.470 45.520 145.790 ;
        RECT 45.600 145.470 45.920 145.790 ;
        RECT 46.000 145.470 46.320 145.790 ;
        RECT 46.400 145.470 46.720 145.790 ;
        RECT 80.045 145.470 80.365 145.790 ;
        RECT 80.445 145.470 80.765 145.790 ;
        RECT 80.845 145.470 81.165 145.790 ;
        RECT 81.245 145.470 81.565 145.790 ;
        RECT 114.890 145.470 115.210 145.790 ;
        RECT 115.290 145.470 115.610 145.790 ;
        RECT 115.690 145.470 116.010 145.790 ;
        RECT 116.090 145.470 116.410 145.790 ;
        RECT 149.735 145.470 150.055 145.790 ;
        RECT 150.135 145.470 150.455 145.790 ;
        RECT 150.535 145.470 150.855 145.790 ;
        RECT 150.935 145.470 151.255 145.790 ;
        RECT 27.780 142.750 28.100 143.070 ;
        RECT 28.180 142.750 28.500 143.070 ;
        RECT 28.580 142.750 28.900 143.070 ;
        RECT 28.980 142.750 29.300 143.070 ;
        RECT 62.625 142.750 62.945 143.070 ;
        RECT 63.025 142.750 63.345 143.070 ;
        RECT 63.425 142.750 63.745 143.070 ;
        RECT 63.825 142.750 64.145 143.070 ;
        RECT 97.470 142.750 97.790 143.070 ;
        RECT 97.870 142.750 98.190 143.070 ;
        RECT 98.270 142.750 98.590 143.070 ;
        RECT 98.670 142.750 98.990 143.070 ;
        RECT 132.315 142.750 132.635 143.070 ;
        RECT 132.715 142.750 133.035 143.070 ;
        RECT 133.115 142.750 133.435 143.070 ;
        RECT 133.515 142.750 133.835 143.070 ;
        RECT 45.200 140.030 45.520 140.350 ;
        RECT 45.600 140.030 45.920 140.350 ;
        RECT 46.000 140.030 46.320 140.350 ;
        RECT 46.400 140.030 46.720 140.350 ;
        RECT 80.045 140.030 80.365 140.350 ;
        RECT 80.445 140.030 80.765 140.350 ;
        RECT 80.845 140.030 81.165 140.350 ;
        RECT 81.245 140.030 81.565 140.350 ;
        RECT 114.890 140.030 115.210 140.350 ;
        RECT 115.290 140.030 115.610 140.350 ;
        RECT 115.690 140.030 116.010 140.350 ;
        RECT 116.090 140.030 116.410 140.350 ;
        RECT 149.735 140.030 150.055 140.350 ;
        RECT 150.135 140.030 150.455 140.350 ;
        RECT 150.535 140.030 150.855 140.350 ;
        RECT 150.935 140.030 151.255 140.350 ;
        RECT 27.780 137.310 28.100 137.630 ;
        RECT 28.180 137.310 28.500 137.630 ;
        RECT 28.580 137.310 28.900 137.630 ;
        RECT 28.980 137.310 29.300 137.630 ;
        RECT 62.625 137.310 62.945 137.630 ;
        RECT 63.025 137.310 63.345 137.630 ;
        RECT 63.425 137.310 63.745 137.630 ;
        RECT 63.825 137.310 64.145 137.630 ;
        RECT 97.470 137.310 97.790 137.630 ;
        RECT 97.870 137.310 98.190 137.630 ;
        RECT 98.270 137.310 98.590 137.630 ;
        RECT 98.670 137.310 98.990 137.630 ;
        RECT 132.315 137.310 132.635 137.630 ;
        RECT 132.715 137.310 133.035 137.630 ;
        RECT 133.115 137.310 133.435 137.630 ;
        RECT 133.515 137.310 133.835 137.630 ;
        RECT 45.200 134.590 45.520 134.910 ;
        RECT 45.600 134.590 45.920 134.910 ;
        RECT 46.000 134.590 46.320 134.910 ;
        RECT 46.400 134.590 46.720 134.910 ;
        RECT 80.045 134.590 80.365 134.910 ;
        RECT 80.445 134.590 80.765 134.910 ;
        RECT 80.845 134.590 81.165 134.910 ;
        RECT 81.245 134.590 81.565 134.910 ;
        RECT 114.890 134.590 115.210 134.910 ;
        RECT 115.290 134.590 115.610 134.910 ;
        RECT 115.690 134.590 116.010 134.910 ;
        RECT 116.090 134.590 116.410 134.910 ;
        RECT 149.735 134.590 150.055 134.910 ;
        RECT 150.135 134.590 150.455 134.910 ;
        RECT 150.535 134.590 150.855 134.910 ;
        RECT 150.935 134.590 151.255 134.910 ;
        RECT 27.780 131.870 28.100 132.190 ;
        RECT 28.180 131.870 28.500 132.190 ;
        RECT 28.580 131.870 28.900 132.190 ;
        RECT 28.980 131.870 29.300 132.190 ;
        RECT 62.625 131.870 62.945 132.190 ;
        RECT 63.025 131.870 63.345 132.190 ;
        RECT 63.425 131.870 63.745 132.190 ;
        RECT 63.825 131.870 64.145 132.190 ;
        RECT 97.470 131.870 97.790 132.190 ;
        RECT 97.870 131.870 98.190 132.190 ;
        RECT 98.270 131.870 98.590 132.190 ;
        RECT 98.670 131.870 98.990 132.190 ;
        RECT 132.315 131.870 132.635 132.190 ;
        RECT 132.715 131.870 133.035 132.190 ;
        RECT 133.115 131.870 133.435 132.190 ;
        RECT 133.515 131.870 133.835 132.190 ;
        RECT 45.200 129.150 45.520 129.470 ;
        RECT 45.600 129.150 45.920 129.470 ;
        RECT 46.000 129.150 46.320 129.470 ;
        RECT 46.400 129.150 46.720 129.470 ;
        RECT 80.045 129.150 80.365 129.470 ;
        RECT 80.445 129.150 80.765 129.470 ;
        RECT 80.845 129.150 81.165 129.470 ;
        RECT 81.245 129.150 81.565 129.470 ;
        RECT 114.890 129.150 115.210 129.470 ;
        RECT 115.290 129.150 115.610 129.470 ;
        RECT 115.690 129.150 116.010 129.470 ;
        RECT 116.090 129.150 116.410 129.470 ;
        RECT 149.735 129.150 150.055 129.470 ;
        RECT 150.135 129.150 150.455 129.470 ;
        RECT 150.535 129.150 150.855 129.470 ;
        RECT 150.935 129.150 151.255 129.470 ;
        RECT 27.780 126.430 28.100 126.750 ;
        RECT 28.180 126.430 28.500 126.750 ;
        RECT 28.580 126.430 28.900 126.750 ;
        RECT 28.980 126.430 29.300 126.750 ;
        RECT 62.625 126.430 62.945 126.750 ;
        RECT 63.025 126.430 63.345 126.750 ;
        RECT 63.425 126.430 63.745 126.750 ;
        RECT 63.825 126.430 64.145 126.750 ;
        RECT 97.470 126.430 97.790 126.750 ;
        RECT 97.870 126.430 98.190 126.750 ;
        RECT 98.270 126.430 98.590 126.750 ;
        RECT 98.670 126.430 98.990 126.750 ;
        RECT 132.315 126.430 132.635 126.750 ;
        RECT 132.715 126.430 133.035 126.750 ;
        RECT 133.115 126.430 133.435 126.750 ;
        RECT 133.515 126.430 133.835 126.750 ;
        RECT 45.200 123.710 45.520 124.030 ;
        RECT 45.600 123.710 45.920 124.030 ;
        RECT 46.000 123.710 46.320 124.030 ;
        RECT 46.400 123.710 46.720 124.030 ;
        RECT 80.045 123.710 80.365 124.030 ;
        RECT 80.445 123.710 80.765 124.030 ;
        RECT 80.845 123.710 81.165 124.030 ;
        RECT 81.245 123.710 81.565 124.030 ;
        RECT 114.890 123.710 115.210 124.030 ;
        RECT 115.290 123.710 115.610 124.030 ;
        RECT 115.690 123.710 116.010 124.030 ;
        RECT 116.090 123.710 116.410 124.030 ;
        RECT 149.735 123.710 150.055 124.030 ;
        RECT 150.135 123.710 150.455 124.030 ;
        RECT 150.535 123.710 150.855 124.030 ;
        RECT 150.935 123.710 151.255 124.030 ;
        RECT 27.780 120.990 28.100 121.310 ;
        RECT 28.180 120.990 28.500 121.310 ;
        RECT 28.580 120.990 28.900 121.310 ;
        RECT 28.980 120.990 29.300 121.310 ;
        RECT 62.625 120.990 62.945 121.310 ;
        RECT 63.025 120.990 63.345 121.310 ;
        RECT 63.425 120.990 63.745 121.310 ;
        RECT 63.825 120.990 64.145 121.310 ;
        RECT 97.470 120.990 97.790 121.310 ;
        RECT 97.870 120.990 98.190 121.310 ;
        RECT 98.270 120.990 98.590 121.310 ;
        RECT 98.670 120.990 98.990 121.310 ;
        RECT 132.315 120.990 132.635 121.310 ;
        RECT 132.715 120.990 133.035 121.310 ;
        RECT 133.115 120.990 133.435 121.310 ;
        RECT 133.515 120.990 133.835 121.310 ;
        RECT 45.200 118.270 45.520 118.590 ;
        RECT 45.600 118.270 45.920 118.590 ;
        RECT 46.000 118.270 46.320 118.590 ;
        RECT 46.400 118.270 46.720 118.590 ;
        RECT 80.045 118.270 80.365 118.590 ;
        RECT 80.445 118.270 80.765 118.590 ;
        RECT 80.845 118.270 81.165 118.590 ;
        RECT 81.245 118.270 81.565 118.590 ;
        RECT 114.890 118.270 115.210 118.590 ;
        RECT 115.290 118.270 115.610 118.590 ;
        RECT 115.690 118.270 116.010 118.590 ;
        RECT 116.090 118.270 116.410 118.590 ;
        RECT 149.735 118.270 150.055 118.590 ;
        RECT 150.135 118.270 150.455 118.590 ;
        RECT 150.535 118.270 150.855 118.590 ;
        RECT 150.935 118.270 151.255 118.590 ;
        RECT 27.780 115.550 28.100 115.870 ;
        RECT 28.180 115.550 28.500 115.870 ;
        RECT 28.580 115.550 28.900 115.870 ;
        RECT 28.980 115.550 29.300 115.870 ;
        RECT 62.625 115.550 62.945 115.870 ;
        RECT 63.025 115.550 63.345 115.870 ;
        RECT 63.425 115.550 63.745 115.870 ;
        RECT 63.825 115.550 64.145 115.870 ;
        RECT 97.470 115.550 97.790 115.870 ;
        RECT 97.870 115.550 98.190 115.870 ;
        RECT 98.270 115.550 98.590 115.870 ;
        RECT 98.670 115.550 98.990 115.870 ;
        RECT 132.315 115.550 132.635 115.870 ;
        RECT 132.715 115.550 133.035 115.870 ;
        RECT 133.115 115.550 133.435 115.870 ;
        RECT 133.515 115.550 133.835 115.870 ;
        RECT 45.200 112.830 45.520 113.150 ;
        RECT 45.600 112.830 45.920 113.150 ;
        RECT 46.000 112.830 46.320 113.150 ;
        RECT 46.400 112.830 46.720 113.150 ;
        RECT 80.045 112.830 80.365 113.150 ;
        RECT 80.445 112.830 80.765 113.150 ;
        RECT 80.845 112.830 81.165 113.150 ;
        RECT 81.245 112.830 81.565 113.150 ;
        RECT 114.890 112.830 115.210 113.150 ;
        RECT 115.290 112.830 115.610 113.150 ;
        RECT 115.690 112.830 116.010 113.150 ;
        RECT 116.090 112.830 116.410 113.150 ;
        RECT 149.735 112.830 150.055 113.150 ;
        RECT 150.135 112.830 150.455 113.150 ;
        RECT 150.535 112.830 150.855 113.150 ;
        RECT 150.935 112.830 151.255 113.150 ;
        RECT 27.780 110.110 28.100 110.430 ;
        RECT 28.180 110.110 28.500 110.430 ;
        RECT 28.580 110.110 28.900 110.430 ;
        RECT 28.980 110.110 29.300 110.430 ;
        RECT 62.625 110.110 62.945 110.430 ;
        RECT 63.025 110.110 63.345 110.430 ;
        RECT 63.425 110.110 63.745 110.430 ;
        RECT 63.825 110.110 64.145 110.430 ;
        RECT 97.470 110.110 97.790 110.430 ;
        RECT 97.870 110.110 98.190 110.430 ;
        RECT 98.270 110.110 98.590 110.430 ;
        RECT 98.670 110.110 98.990 110.430 ;
        RECT 132.315 110.110 132.635 110.430 ;
        RECT 132.715 110.110 133.035 110.430 ;
        RECT 133.115 110.110 133.435 110.430 ;
        RECT 133.515 110.110 133.835 110.430 ;
        RECT 45.200 107.390 45.520 107.710 ;
        RECT 45.600 107.390 45.920 107.710 ;
        RECT 46.000 107.390 46.320 107.710 ;
        RECT 46.400 107.390 46.720 107.710 ;
        RECT 80.045 107.390 80.365 107.710 ;
        RECT 80.445 107.390 80.765 107.710 ;
        RECT 80.845 107.390 81.165 107.710 ;
        RECT 81.245 107.390 81.565 107.710 ;
        RECT 114.890 107.390 115.210 107.710 ;
        RECT 115.290 107.390 115.610 107.710 ;
        RECT 115.690 107.390 116.010 107.710 ;
        RECT 116.090 107.390 116.410 107.710 ;
        RECT 149.735 107.390 150.055 107.710 ;
        RECT 150.135 107.390 150.455 107.710 ;
        RECT 150.535 107.390 150.855 107.710 ;
        RECT 150.935 107.390 151.255 107.710 ;
        RECT 27.780 104.670 28.100 104.990 ;
        RECT 28.180 104.670 28.500 104.990 ;
        RECT 28.580 104.670 28.900 104.990 ;
        RECT 28.980 104.670 29.300 104.990 ;
        RECT 62.625 104.670 62.945 104.990 ;
        RECT 63.025 104.670 63.345 104.990 ;
        RECT 63.425 104.670 63.745 104.990 ;
        RECT 63.825 104.670 64.145 104.990 ;
        RECT 97.470 104.670 97.790 104.990 ;
        RECT 97.870 104.670 98.190 104.990 ;
        RECT 98.270 104.670 98.590 104.990 ;
        RECT 98.670 104.670 98.990 104.990 ;
        RECT 132.315 104.670 132.635 104.990 ;
        RECT 132.715 104.670 133.035 104.990 ;
        RECT 133.115 104.670 133.435 104.990 ;
        RECT 133.515 104.670 133.835 104.990 ;
        RECT 45.200 101.950 45.520 102.270 ;
        RECT 45.600 101.950 45.920 102.270 ;
        RECT 46.000 101.950 46.320 102.270 ;
        RECT 46.400 101.950 46.720 102.270 ;
        RECT 80.045 101.950 80.365 102.270 ;
        RECT 80.445 101.950 80.765 102.270 ;
        RECT 80.845 101.950 81.165 102.270 ;
        RECT 81.245 101.950 81.565 102.270 ;
        RECT 114.890 101.950 115.210 102.270 ;
        RECT 115.290 101.950 115.610 102.270 ;
        RECT 115.690 101.950 116.010 102.270 ;
        RECT 116.090 101.950 116.410 102.270 ;
        RECT 149.735 101.950 150.055 102.270 ;
        RECT 150.135 101.950 150.455 102.270 ;
        RECT 150.535 101.950 150.855 102.270 ;
        RECT 150.935 101.950 151.255 102.270 ;
        RECT 27.780 99.230 28.100 99.550 ;
        RECT 28.180 99.230 28.500 99.550 ;
        RECT 28.580 99.230 28.900 99.550 ;
        RECT 28.980 99.230 29.300 99.550 ;
        RECT 62.625 99.230 62.945 99.550 ;
        RECT 63.025 99.230 63.345 99.550 ;
        RECT 63.425 99.230 63.745 99.550 ;
        RECT 63.825 99.230 64.145 99.550 ;
        RECT 97.470 99.230 97.790 99.550 ;
        RECT 97.870 99.230 98.190 99.550 ;
        RECT 98.270 99.230 98.590 99.550 ;
        RECT 98.670 99.230 98.990 99.550 ;
        RECT 132.315 99.230 132.635 99.550 ;
        RECT 132.715 99.230 133.035 99.550 ;
        RECT 133.115 99.230 133.435 99.550 ;
        RECT 133.515 99.230 133.835 99.550 ;
        RECT 45.200 96.510 45.520 96.830 ;
        RECT 45.600 96.510 45.920 96.830 ;
        RECT 46.000 96.510 46.320 96.830 ;
        RECT 46.400 96.510 46.720 96.830 ;
        RECT 80.045 96.510 80.365 96.830 ;
        RECT 80.445 96.510 80.765 96.830 ;
        RECT 80.845 96.510 81.165 96.830 ;
        RECT 81.245 96.510 81.565 96.830 ;
        RECT 114.890 96.510 115.210 96.830 ;
        RECT 115.290 96.510 115.610 96.830 ;
        RECT 115.690 96.510 116.010 96.830 ;
        RECT 116.090 96.510 116.410 96.830 ;
        RECT 149.735 96.510 150.055 96.830 ;
        RECT 150.135 96.510 150.455 96.830 ;
        RECT 150.535 96.510 150.855 96.830 ;
        RECT 150.935 96.510 151.255 96.830 ;
        RECT 27.780 93.790 28.100 94.110 ;
        RECT 28.180 93.790 28.500 94.110 ;
        RECT 28.580 93.790 28.900 94.110 ;
        RECT 28.980 93.790 29.300 94.110 ;
        RECT 62.625 93.790 62.945 94.110 ;
        RECT 63.025 93.790 63.345 94.110 ;
        RECT 63.425 93.790 63.745 94.110 ;
        RECT 63.825 93.790 64.145 94.110 ;
        RECT 97.470 93.790 97.790 94.110 ;
        RECT 97.870 93.790 98.190 94.110 ;
        RECT 98.270 93.790 98.590 94.110 ;
        RECT 98.670 93.790 98.990 94.110 ;
        RECT 132.315 93.790 132.635 94.110 ;
        RECT 132.715 93.790 133.035 94.110 ;
        RECT 133.115 93.790 133.435 94.110 ;
        RECT 133.515 93.790 133.835 94.110 ;
        RECT 45.200 91.070 45.520 91.390 ;
        RECT 45.600 91.070 45.920 91.390 ;
        RECT 46.000 91.070 46.320 91.390 ;
        RECT 46.400 91.070 46.720 91.390 ;
        RECT 80.045 91.070 80.365 91.390 ;
        RECT 80.445 91.070 80.765 91.390 ;
        RECT 80.845 91.070 81.165 91.390 ;
        RECT 81.245 91.070 81.565 91.390 ;
        RECT 114.890 91.070 115.210 91.390 ;
        RECT 115.290 91.070 115.610 91.390 ;
        RECT 115.690 91.070 116.010 91.390 ;
        RECT 116.090 91.070 116.410 91.390 ;
        RECT 149.735 91.070 150.055 91.390 ;
        RECT 150.135 91.070 150.455 91.390 ;
        RECT 150.535 91.070 150.855 91.390 ;
        RECT 150.935 91.070 151.255 91.390 ;
        RECT 27.780 88.350 28.100 88.670 ;
        RECT 28.180 88.350 28.500 88.670 ;
        RECT 28.580 88.350 28.900 88.670 ;
        RECT 28.980 88.350 29.300 88.670 ;
        RECT 62.625 88.350 62.945 88.670 ;
        RECT 63.025 88.350 63.345 88.670 ;
        RECT 63.425 88.350 63.745 88.670 ;
        RECT 63.825 88.350 64.145 88.670 ;
        RECT 97.470 88.350 97.790 88.670 ;
        RECT 97.870 88.350 98.190 88.670 ;
        RECT 98.270 88.350 98.590 88.670 ;
        RECT 98.670 88.350 98.990 88.670 ;
        RECT 132.315 88.350 132.635 88.670 ;
        RECT 132.715 88.350 133.035 88.670 ;
        RECT 133.115 88.350 133.435 88.670 ;
        RECT 133.515 88.350 133.835 88.670 ;
        RECT 45.200 85.630 45.520 85.950 ;
        RECT 45.600 85.630 45.920 85.950 ;
        RECT 46.000 85.630 46.320 85.950 ;
        RECT 46.400 85.630 46.720 85.950 ;
        RECT 80.045 85.630 80.365 85.950 ;
        RECT 80.445 85.630 80.765 85.950 ;
        RECT 80.845 85.630 81.165 85.950 ;
        RECT 81.245 85.630 81.565 85.950 ;
        RECT 114.890 85.630 115.210 85.950 ;
        RECT 115.290 85.630 115.610 85.950 ;
        RECT 115.690 85.630 116.010 85.950 ;
        RECT 116.090 85.630 116.410 85.950 ;
        RECT 149.735 85.630 150.055 85.950 ;
        RECT 150.135 85.630 150.455 85.950 ;
        RECT 150.535 85.630 150.855 85.950 ;
        RECT 150.935 85.630 151.255 85.950 ;
        RECT 27.780 82.910 28.100 83.230 ;
        RECT 28.180 82.910 28.500 83.230 ;
        RECT 28.580 82.910 28.900 83.230 ;
        RECT 28.980 82.910 29.300 83.230 ;
        RECT 62.625 82.910 62.945 83.230 ;
        RECT 63.025 82.910 63.345 83.230 ;
        RECT 63.425 82.910 63.745 83.230 ;
        RECT 63.825 82.910 64.145 83.230 ;
        RECT 97.470 82.910 97.790 83.230 ;
        RECT 97.870 82.910 98.190 83.230 ;
        RECT 98.270 82.910 98.590 83.230 ;
        RECT 98.670 82.910 98.990 83.230 ;
        RECT 132.315 82.910 132.635 83.230 ;
        RECT 132.715 82.910 133.035 83.230 ;
        RECT 133.115 82.910 133.435 83.230 ;
        RECT 133.515 82.910 133.835 83.230 ;
        RECT 45.200 80.190 45.520 80.510 ;
        RECT 45.600 80.190 45.920 80.510 ;
        RECT 46.000 80.190 46.320 80.510 ;
        RECT 46.400 80.190 46.720 80.510 ;
        RECT 80.045 80.190 80.365 80.510 ;
        RECT 80.445 80.190 80.765 80.510 ;
        RECT 80.845 80.190 81.165 80.510 ;
        RECT 81.245 80.190 81.565 80.510 ;
        RECT 114.890 80.190 115.210 80.510 ;
        RECT 115.290 80.190 115.610 80.510 ;
        RECT 115.690 80.190 116.010 80.510 ;
        RECT 116.090 80.190 116.410 80.510 ;
        RECT 149.735 80.190 150.055 80.510 ;
        RECT 150.135 80.190 150.455 80.510 ;
        RECT 150.535 80.190 150.855 80.510 ;
        RECT 150.935 80.190 151.255 80.510 ;
        RECT 27.780 77.470 28.100 77.790 ;
        RECT 28.180 77.470 28.500 77.790 ;
        RECT 28.580 77.470 28.900 77.790 ;
        RECT 28.980 77.470 29.300 77.790 ;
        RECT 62.625 77.470 62.945 77.790 ;
        RECT 63.025 77.470 63.345 77.790 ;
        RECT 63.425 77.470 63.745 77.790 ;
        RECT 63.825 77.470 64.145 77.790 ;
        RECT 97.470 77.470 97.790 77.790 ;
        RECT 97.870 77.470 98.190 77.790 ;
        RECT 98.270 77.470 98.590 77.790 ;
        RECT 98.670 77.470 98.990 77.790 ;
        RECT 132.315 77.470 132.635 77.790 ;
        RECT 132.715 77.470 133.035 77.790 ;
        RECT 133.115 77.470 133.435 77.790 ;
        RECT 133.515 77.470 133.835 77.790 ;
        RECT 45.200 74.750 45.520 75.070 ;
        RECT 45.600 74.750 45.920 75.070 ;
        RECT 46.000 74.750 46.320 75.070 ;
        RECT 46.400 74.750 46.720 75.070 ;
        RECT 80.045 74.750 80.365 75.070 ;
        RECT 80.445 74.750 80.765 75.070 ;
        RECT 80.845 74.750 81.165 75.070 ;
        RECT 81.245 74.750 81.565 75.070 ;
        RECT 114.890 74.750 115.210 75.070 ;
        RECT 115.290 74.750 115.610 75.070 ;
        RECT 115.690 74.750 116.010 75.070 ;
        RECT 116.090 74.750 116.410 75.070 ;
        RECT 149.735 74.750 150.055 75.070 ;
        RECT 150.135 74.750 150.455 75.070 ;
        RECT 150.535 74.750 150.855 75.070 ;
        RECT 150.935 74.750 151.255 75.070 ;
        RECT 27.680 72.680 29.300 74.270 ;
        RECT 62.580 72.680 64.160 74.400 ;
        RECT 97.390 72.580 98.950 74.300 ;
        RECT 51.110 60.980 53.680 63.040 ;
        RECT 62.600 61.130 64.180 63.080 ;
        RECT 132.410 72.560 133.880 74.030 ;
        RECT 97.370 61.090 98.950 63.040 ;
        RECT 132.220 60.770 134.340 62.770 ;
        RECT 55.340 55.020 76.610 59.300 ;
        RECT 95.400 55.090 105.220 59.770 ;
        RECT 117.310 54.830 134.530 58.370 ;
        RECT 55.390 11.400 64.190 18.240 ;
        RECT 74.330 11.280 83.680 18.120 ;
        RECT 46.165 4.785 46.755 5.375 ;
        RECT 94.640 11.670 105.730 18.200 ;
        RECT 117.320 13.120 127.600 18.610 ;
        RECT 135.980 13.520 146.160 18.400 ;
        RECT 150.535 4.115 151.125 4.705 ;
        RECT 68.245 2.245 68.835 2.835 ;
        RECT 90.325 2.335 90.915 2.925 ;
        RECT 112.405 2.545 112.995 3.135 ;
        RECT 134.485 2.775 135.075 3.365 ;
        RECT 150.530 2.470 151.130 3.070 ;
      LAYER met4 ;
        RECT 63.170 224.760 63.180 225.250 ;
        RECT 140.130 224.760 140.150 225.480 ;
        RECT 143.810 224.760 143.830 225.350 ;
        RECT 147.480 224.760 147.510 225.140 ;
        RECT 3.990 224.390 4.290 224.760 ;
        RECT 7.670 224.390 7.970 224.760 ;
        RECT 11.350 224.390 11.650 224.760 ;
        RECT 15.030 224.390 15.330 224.760 ;
        RECT 18.710 224.390 19.010 224.760 ;
        RECT 22.390 224.390 22.690 224.760 ;
        RECT 26.070 224.390 26.370 224.760 ;
        RECT 29.750 224.390 30.050 224.760 ;
        RECT 33.430 224.390 33.730 224.760 ;
        RECT 37.110 224.390 37.410 224.760 ;
        RECT 40.790 224.390 41.090 224.760 ;
        RECT 44.470 224.390 44.770 224.760 ;
        RECT 48.150 224.390 48.450 224.760 ;
        RECT 51.830 224.390 52.130 224.760 ;
        RECT 55.510 224.390 55.810 224.760 ;
        RECT 59.190 224.390 59.490 224.760 ;
        RECT 2.050 224.090 59.490 224.390 ;
        RECT 62.870 224.155 63.180 224.760 ;
        RECT 2.050 220.760 2.350 224.090 ;
        RECT 62.865 223.750 63.180 224.155 ;
        RECT 66.540 224.210 66.850 224.760 ;
        RECT 70.230 224.250 70.530 224.760 ;
        RECT 66.540 223.770 66.860 224.210 ;
        RECT 60.015 223.720 60.345 223.735 ;
        RECT 62.865 223.725 63.175 223.750 ;
        RECT 61.335 223.720 63.175 223.725 ;
        RECT 60.015 223.420 63.175 223.720 ;
        RECT 60.015 223.405 60.345 223.420 ;
        RECT 61.335 223.415 63.175 223.420 ;
        RECT 66.560 222.670 66.860 223.770 ;
        RECT 25.000 222.370 66.860 222.670 ;
        RECT 70.230 223.770 70.540 224.250 ;
        RECT 73.910 223.800 74.210 224.760 ;
        RECT 25.000 218.835 25.300 222.370 ;
        RECT 70.230 221.875 70.530 223.770 ;
        RECT 73.880 223.510 74.210 223.800 ;
        RECT 74.975 223.890 75.305 223.905 ;
        RECT 77.590 223.890 77.890 224.760 ;
        RECT 74.975 223.590 77.900 223.890 ;
        RECT 74.975 223.575 75.305 223.590 ;
        RECT 70.215 221.545 70.545 221.875 ;
        RECT 73.880 221.835 74.180 223.510 ;
        RECT 73.865 221.505 74.195 221.835 ;
        RECT 81.270 220.510 81.570 224.760 ;
        RECT 84.950 224.030 85.250 224.760 ;
        RECT 88.630 224.490 88.930 224.760 ;
        RECT 84.950 223.370 85.260 224.030 ;
        RECT 84.960 221.580 85.260 223.370 ;
        RECT 81.260 220.020 81.570 220.510 ;
        RECT 83.820 221.280 85.260 221.580 ;
        RECT 88.620 223.370 88.930 224.490 ;
        RECT 129.555 223.890 129.885 223.905 ;
        RECT 136.470 223.890 136.770 224.760 ;
        RECT 129.555 223.590 136.770 223.890 ;
        RECT 129.555 223.575 129.885 223.590 ;
        RECT 81.260 219.330 81.560 220.020 ;
        RECT 72.800 219.030 81.560 219.330 ;
        RECT 24.985 218.505 25.315 218.835 ;
        RECT 72.015 217.200 72.345 217.215 ;
        RECT 72.800 217.200 73.100 219.030 ;
        RECT 83.820 218.055 84.120 221.280 ;
        RECT 87.175 218.750 87.505 218.765 ;
        RECT 88.620 218.750 88.920 223.370 ;
        RECT 140.130 222.970 140.430 224.760 ;
        RECT 105.960 222.670 140.430 222.970 ;
        RECT 143.810 222.815 144.110 224.760 ;
        RECT 105.960 220.165 106.260 222.670 ;
        RECT 143.795 222.485 144.125 222.815 ;
        RECT 147.480 220.460 147.780 224.760 ;
        RECT 151.190 222.595 151.490 224.760 ;
        RECT 151.175 222.265 151.505 222.595 ;
        RECT 105.945 219.835 106.275 220.165 ;
        RECT 126.200 220.160 147.780 220.460 ;
        RECT 126.200 219.585 126.500 220.160 ;
        RECT 126.185 219.255 126.515 219.585 ;
        RECT 87.175 218.450 88.920 218.750 ;
        RECT 87.175 218.435 87.505 218.450 ;
        RECT 83.805 217.725 84.135 218.055 ;
        RECT 153.645 217.700 153.975 217.715 ;
        RECT 154.870 217.700 155.170 224.760 ;
        RECT 153.645 217.400 155.170 217.700 ;
        RECT 153.645 217.385 153.975 217.400 ;
        RECT 72.015 216.900 73.100 217.200 ;
        RECT 72.015 216.885 72.345 216.900 ;
        RECT 27.740 76.710 29.340 213.870 ;
        RECT 27.680 74.275 29.380 76.710 ;
        RECT 45.160 74.670 46.760 213.870 ;
        RECT 62.585 76.840 64.185 213.870 ;
        RECT 75.815 175.725 76.145 176.055 ;
        RECT 75.830 154.295 76.130 175.725 ;
        RECT 75.815 153.965 76.145 154.295 ;
        RECT 27.675 72.680 29.380 74.275 ;
        RECT 27.675 72.675 29.305 72.680 ;
        RECT 45.200 70.780 46.700 74.670 ;
        RECT 62.580 74.405 64.190 76.840 ;
        RECT 80.005 74.670 81.605 213.870 ;
        RECT 97.430 76.840 99.030 213.870 ;
        RECT 62.575 72.680 64.190 74.405 ;
        RECT 62.575 72.675 64.165 72.680 ;
        RECT 80.050 70.780 81.550 74.670 ;
        RECT 97.390 74.305 99.080 76.840 ;
        RECT 114.850 74.670 116.450 213.870 ;
        RECT 132.275 76.840 133.875 213.870 ;
        RECT 97.385 72.580 99.080 74.305 ;
        RECT 97.385 72.575 98.955 72.580 ;
        RECT 114.950 70.780 116.450 74.670 ;
        RECT 132.250 72.580 133.940 76.840 ;
        RECT 149.695 74.670 151.295 213.870 ;
        RECT 132.250 72.560 133.885 72.580 ;
        RECT 132.405 72.555 133.885 72.560 ;
        RECT 149.760 70.780 151.260 74.670 ;
        RECT 2.500 69.280 151.260 70.780 ;
        RECT 149.910 63.120 157.210 63.150 ;
        RECT 50.990 54.710 158.080 63.120 ;
        RECT 50.990 54.590 93.820 54.710 ;
        RECT 107.870 54.590 158.080 54.710 ;
        RECT 149.910 54.570 157.210 54.590 ;
        RECT 99.610 19.000 100.800 19.040 ;
        RECT 51.320 18.980 152.970 19.000 ;
        RECT 2.500 10.470 152.970 18.980 ;
        RECT 46.160 1.000 46.760 5.380 ;
        RECT 68.240 1.000 68.840 2.840 ;
        RECT 90.320 1.000 90.920 2.930 ;
        RECT 112.400 1.000 113.000 3.140 ;
        RECT 134.480 1.000 135.080 3.370 ;
        RECT 150.530 3.075 151.130 4.710 ;
        RECT 150.525 3.070 151.135 3.075 ;
        RECT 150.525 2.470 157.160 3.070 ;
        RECT 150.525 2.465 151.135 2.470 ;
        RECT 156.560 1.000 157.160 2.470 ;
  END
END tt_um_argunda_tiny_opamp
END LIBRARY


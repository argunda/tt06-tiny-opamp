magic
tech sky130A
magscale 1 2
timestamp 1713541782
<< viali >>
rect 11345 28169 11379 28203
rect 11161 27965 11195 27999
rect 15669 27965 15703 27999
rect 17601 27965 17635 27999
rect 19257 27965 19291 27999
rect 20177 27965 20211 27999
rect 20453 27965 20487 27999
rect 21833 27965 21867 27999
rect 24041 27965 24075 27999
rect 25789 27965 25823 27999
rect 15853 27829 15887 27863
rect 17785 27829 17819 27863
rect 19901 27829 19935 27863
rect 20085 27829 20119 27863
rect 20269 27829 20303 27863
rect 21649 27829 21683 27863
rect 23857 27829 23891 27863
rect 25881 27829 25915 27863
rect 6745 27625 6779 27659
rect 14565 27625 14599 27659
rect 15209 27625 15243 27659
rect 19073 27625 19107 27659
rect 1409 27557 1443 27591
rect 3801 27557 3835 27591
rect 4629 27557 4663 27591
rect 5181 27557 5215 27591
rect 15025 27557 15059 27591
rect 15393 27557 15427 27591
rect 15761 27557 15795 27591
rect 19432 27557 19466 27591
rect 1777 27489 1811 27523
rect 2596 27489 2630 27523
rect 4169 27489 4203 27523
rect 4813 27489 4847 27523
rect 4905 27489 4939 27523
rect 5089 27489 5123 27523
rect 5549 27489 5583 27523
rect 6009 27489 6043 27523
rect 6377 27489 6411 27523
rect 7205 27489 7239 27523
rect 7573 27489 7607 27523
rect 8217 27489 8251 27523
rect 8953 27489 8987 27523
rect 9413 27489 9447 27523
rect 9680 27489 9714 27523
rect 11161 27489 11195 27523
rect 11417 27489 11451 27523
rect 12725 27489 12759 27523
rect 13185 27489 13219 27523
rect 13441 27489 13475 27523
rect 16385 27489 16419 27523
rect 17693 27489 17727 27523
rect 17960 27489 17994 27523
rect 20637 27489 20671 27523
rect 21097 27489 21131 27523
rect 22681 27489 22715 27523
rect 23296 27489 23330 27523
rect 2329 27421 2363 27455
rect 6285 27421 6319 27455
rect 7665 27421 7699 27455
rect 8125 27421 8159 27455
rect 8585 27421 8619 27455
rect 8861 27421 8895 27455
rect 16129 27421 16163 27455
rect 19165 27421 19199 27455
rect 22937 27421 22971 27455
rect 23029 27421 23063 27455
rect 7021 27353 7055 27387
rect 7941 27353 7975 27387
rect 12541 27353 12575 27387
rect 14657 27353 14691 27387
rect 20545 27353 20579 27387
rect 21557 27353 21591 27387
rect 3709 27285 3743 27319
rect 4445 27285 4479 27319
rect 4997 27285 5031 27319
rect 5825 27285 5859 27319
rect 9229 27285 9263 27319
rect 10793 27285 10827 27319
rect 13001 27285 13035 27319
rect 15025 27285 15059 27319
rect 17509 27285 17543 27319
rect 20729 27285 20763 27319
rect 21005 27285 21039 27319
rect 24409 27285 24443 27319
rect 2789 27081 2823 27115
rect 3433 27081 3467 27115
rect 7849 27081 7883 27115
rect 8953 27081 8987 27115
rect 11345 27081 11379 27115
rect 13093 27081 13127 27115
rect 15025 27081 15059 27115
rect 18337 27081 18371 27115
rect 23029 27081 23063 27115
rect 23213 27081 23247 27115
rect 3249 27013 3283 27047
rect 4905 27013 4939 27047
rect 7757 27013 7791 27047
rect 11805 27013 11839 27047
rect 16773 27013 16807 27047
rect 22017 27013 22051 27047
rect 11713 26945 11747 26979
rect 12357 26945 12391 26979
rect 15393 26945 15427 26979
rect 17509 26945 17543 26979
rect 22385 26945 22419 26979
rect 24869 26945 24903 26979
rect 2973 26877 3007 26911
rect 3801 26877 3835 26911
rect 4077 26877 4111 26911
rect 4353 26877 4387 26911
rect 6018 26877 6052 26911
rect 6285 26877 6319 26911
rect 8769 26877 8803 26911
rect 11253 26877 11287 26911
rect 12449 26877 12483 26911
rect 12633 26877 12667 26911
rect 12725 26877 12759 26911
rect 12817 26877 12851 26911
rect 14657 26877 14691 26911
rect 15117 26877 15151 26911
rect 15301 26877 15335 26911
rect 17877 26877 17911 26911
rect 18245 26877 18279 26911
rect 19073 26877 19107 26911
rect 20637 26877 20671 26911
rect 20904 26877 20938 26911
rect 23305 26877 23339 26911
rect 7389 26809 7423 26843
rect 12173 26809 12207 26843
rect 14841 26809 14875 26843
rect 15209 26809 15243 26843
rect 15638 26809 15672 26843
rect 19340 26809 19374 26843
rect 3433 26741 3467 26775
rect 3893 26741 3927 26775
rect 4261 26741 4295 26775
rect 11989 26741 12023 26775
rect 12081 26741 12115 26775
rect 16957 26741 16991 26775
rect 18061 26741 18095 26775
rect 20453 26741 20487 26775
rect 24317 26741 24351 26775
rect 4563 26537 4597 26571
rect 6101 26537 6135 26571
rect 7389 26537 7423 26571
rect 7757 26537 7791 26571
rect 8033 26537 8067 26571
rect 10425 26537 10459 26571
rect 14197 26537 14231 26571
rect 14749 26537 14783 26571
rect 14841 26537 14875 26571
rect 4353 26469 4387 26503
rect 13829 26469 13863 26503
rect 14059 26435 14093 26469
rect 7297 26401 7331 26435
rect 7481 26401 7515 26435
rect 7573 26401 7607 26435
rect 7849 26401 7883 26435
rect 7941 26401 7975 26435
rect 8125 26401 8159 26435
rect 9321 26401 9355 26435
rect 10057 26401 10091 26435
rect 12173 26401 12207 26435
rect 12265 26401 12299 26435
rect 12449 26401 12483 26435
rect 12541 26401 12575 26435
rect 12633 26401 12667 26435
rect 14565 26401 14599 26435
rect 15117 26401 15151 26435
rect 16497 26401 16531 26435
rect 16753 26401 16787 26435
rect 20830 26401 20864 26435
rect 6561 26333 6595 26367
rect 9229 26333 9263 26367
rect 9965 26333 9999 26367
rect 12725 26333 12759 26367
rect 14381 26333 14415 26367
rect 14841 26333 14875 26367
rect 15025 26333 15059 26367
rect 21097 26333 21131 26367
rect 4721 26265 4755 26299
rect 6285 26265 6319 26299
rect 7573 26265 7607 26299
rect 9689 26265 9723 26299
rect 17877 26265 17911 26299
rect 19717 26265 19751 26299
rect 4537 26197 4571 26231
rect 14013 26197 14047 26231
rect 6009 25993 6043 26027
rect 6377 25993 6411 26027
rect 8401 25993 8435 26027
rect 11897 25993 11931 26027
rect 12541 25993 12575 26027
rect 13093 25993 13127 26027
rect 15301 25993 15335 26027
rect 16313 25993 16347 26027
rect 20913 25993 20947 26027
rect 3065 25925 3099 25959
rect 6469 25925 6503 25959
rect 6929 25925 6963 25959
rect 10977 25925 11011 25959
rect 15485 25925 15519 25959
rect 3801 25857 3835 25891
rect 11069 25857 11103 25891
rect 21281 25857 21315 25891
rect 1685 25789 1719 25823
rect 4169 25789 4203 25823
rect 5825 25789 5859 25823
rect 6929 25789 6963 25823
rect 7205 25789 7239 25823
rect 8585 25789 8619 25823
rect 8861 25789 8895 25823
rect 11345 25789 11379 25823
rect 11621 25789 11655 25823
rect 12173 25789 12207 25823
rect 12909 25789 12943 25823
rect 13001 25789 13035 25823
rect 13185 25789 13219 25823
rect 14933 25789 14967 25823
rect 16129 25789 16163 25823
rect 18337 25789 18371 25823
rect 20085 25789 20119 25823
rect 20361 25789 20395 25823
rect 1952 25721 1986 25755
rect 4436 25721 4470 25755
rect 6837 25721 6871 25755
rect 10609 25721 10643 25755
rect 12725 25721 12759 25755
rect 19818 25721 19852 25755
rect 21548 25721 21582 25755
rect 3249 25653 3283 25687
rect 5549 25653 5583 25687
rect 6285 25653 6319 25687
rect 7113 25653 7147 25687
rect 8769 25653 8803 25687
rect 11161 25653 11195 25687
rect 11529 25653 11563 25687
rect 11713 25653 11747 25687
rect 15301 25653 15335 25687
rect 18521 25653 18555 25687
rect 18705 25653 18739 25687
rect 22661 25653 22695 25687
rect 3157 25449 3191 25483
rect 3709 25449 3743 25483
rect 3877 25449 3911 25483
rect 4721 25449 4755 25483
rect 7941 25449 7975 25483
rect 8309 25449 8343 25483
rect 9137 25449 9171 25483
rect 12265 25449 12299 25483
rect 14397 25449 14431 25483
rect 14565 25449 14599 25483
rect 15301 25449 15335 25483
rect 18429 25449 18463 25483
rect 21741 25449 21775 25483
rect 4077 25381 4111 25415
rect 13645 25381 13679 25415
rect 13861 25381 13895 25415
rect 14197 25381 14231 25415
rect 14933 25381 14967 25415
rect 15117 25381 15151 25415
rect 18061 25381 18095 25415
rect 18277 25381 18311 25415
rect 2973 25313 3007 25347
rect 3249 25313 3283 25347
rect 3341 25313 3375 25347
rect 3433 25313 3467 25347
rect 4905 25313 4939 25347
rect 7849 25313 7883 25347
rect 8033 25313 8067 25347
rect 8125 25313 8159 25347
rect 8309 25313 8343 25347
rect 8769 25313 8803 25347
rect 12725 25313 12759 25347
rect 16773 25313 16807 25347
rect 18521 25313 18555 25347
rect 19616 25313 19650 25347
rect 21281 25313 21315 25347
rect 21465 25313 21499 25347
rect 21649 25313 21683 25347
rect 21925 25313 21959 25347
rect 24061 25313 24095 25347
rect 24317 25313 24351 25347
rect 3617 25245 3651 25279
rect 8677 25245 8711 25279
rect 16865 25245 16899 25279
rect 19073 25245 19107 25279
rect 19349 25245 19383 25279
rect 2973 25177 3007 25211
rect 3525 25177 3559 25211
rect 14013 25177 14047 25211
rect 3893 25109 3927 25143
rect 12633 25109 12667 25143
rect 13829 25109 13863 25143
rect 14381 25109 14415 25143
rect 17141 25109 17175 25143
rect 18245 25109 18279 25143
rect 20729 25109 20763 25143
rect 22937 25109 22971 25143
rect 6653 24905 6687 24939
rect 7205 24905 7239 24939
rect 10241 24905 10275 24939
rect 12541 24905 12575 24939
rect 15209 24905 15243 24939
rect 18889 24905 18923 24939
rect 19625 24905 19659 24939
rect 21557 24905 21591 24939
rect 22477 24905 22511 24939
rect 6285 24837 6319 24871
rect 14841 24837 14875 24871
rect 6469 24769 6503 24803
rect 7021 24769 7055 24803
rect 7113 24769 7147 24803
rect 10517 24769 10551 24803
rect 12357 24769 12391 24803
rect 16221 24769 16255 24803
rect 20913 24769 20947 24803
rect 22661 24769 22695 24803
rect 6561 24701 6595 24735
rect 7297 24701 7331 24735
rect 7389 24701 7423 24735
rect 9873 24701 9907 24735
rect 12817 24701 12851 24735
rect 13921 24701 13955 24735
rect 14381 24701 14415 24735
rect 15945 24701 15979 24735
rect 19809 24701 19843 24735
rect 22385 24701 22419 24735
rect 6009 24633 6043 24667
rect 10241 24633 10275 24667
rect 10784 24633 10818 24667
rect 14105 24633 14139 24667
rect 14565 24633 14599 24667
rect 16466 24633 16500 24667
rect 18705 24633 18739 24667
rect 19349 24633 19383 24667
rect 19533 24633 19567 24667
rect 21189 24633 21223 24667
rect 10425 24565 10459 24599
rect 11897 24565 11931 24599
rect 14289 24565 14323 24599
rect 14749 24565 14783 24599
rect 15209 24565 15243 24599
rect 15393 24565 15427 24599
rect 16129 24565 16163 24599
rect 17601 24565 17635 24599
rect 18905 24565 18939 24599
rect 19073 24565 19107 24599
rect 19165 24565 19199 24599
rect 21097 24565 21131 24599
rect 22661 24565 22695 24599
rect 4353 24361 4387 24395
rect 4813 24361 4847 24395
rect 8309 24361 8343 24395
rect 9755 24361 9789 24395
rect 10701 24361 10735 24395
rect 10977 24361 11011 24395
rect 14105 24361 14139 24395
rect 14657 24361 14691 24395
rect 15393 24361 15427 24395
rect 18797 24361 18831 24395
rect 18981 24361 19015 24395
rect 19993 24361 20027 24395
rect 20453 24361 20487 24395
rect 6929 24293 6963 24327
rect 9965 24293 9999 24327
rect 16374 24293 16408 24327
rect 1317 24225 1351 24259
rect 1768 24225 1802 24259
rect 2973 24225 3007 24259
rect 3240 24225 3274 24259
rect 4629 24225 4663 24259
rect 4721 24225 4755 24259
rect 5181 24225 5215 24259
rect 6193 24225 6227 24259
rect 7297 24225 7331 24259
rect 7941 24225 7975 24259
rect 9505 24225 9539 24259
rect 10517 24225 10551 24259
rect 11254 24225 11288 24259
rect 11621 24225 11655 24259
rect 11805 24225 11839 24259
rect 12449 24225 12483 24259
rect 12541 24225 12575 24259
rect 13921 24225 13955 24259
rect 14289 24225 14323 24259
rect 15209 24225 15243 24259
rect 16129 24225 16163 24259
rect 17969 24225 18003 24259
rect 18153 24225 18187 24259
rect 18245 24225 18279 24259
rect 18521 24225 18555 24259
rect 18922 24225 18956 24259
rect 20361 24225 20395 24259
rect 22017 24225 22051 24259
rect 22109 24225 22143 24259
rect 22293 24225 22327 24259
rect 22569 24225 22603 24259
rect 23121 24225 23155 24259
rect 23305 24225 23339 24259
rect 23397 24225 23431 24259
rect 23581 24225 23615 24259
rect 24124 24225 24158 24259
rect 1501 24157 1535 24191
rect 6009 24157 6043 24191
rect 6101 24157 6135 24191
rect 6285 24157 6319 24191
rect 7205 24157 7239 24191
rect 7665 24157 7699 24191
rect 7849 24157 7883 24191
rect 11161 24157 11195 24191
rect 11345 24157 11379 24191
rect 11437 24157 11471 24191
rect 13737 24157 13771 24191
rect 19441 24157 19475 24191
rect 20545 24157 20579 24191
rect 22661 24157 22695 24191
rect 23857 24157 23891 24191
rect 4445 24089 4479 24123
rect 6653 24089 6687 24123
rect 9597 24089 9631 24123
rect 14841 24089 14875 24123
rect 19349 24089 19383 24123
rect 22937 24089 22971 24123
rect 1133 24021 1167 24055
rect 2881 24021 2915 24055
rect 4997 24021 5031 24055
rect 5365 24021 5399 24055
rect 5825 24021 5859 24055
rect 6469 24021 6503 24055
rect 9045 24021 9079 24055
rect 9413 24021 9447 24055
rect 9781 24021 9815 24055
rect 11805 24021 11839 24055
rect 14657 24021 14691 24055
rect 17509 24021 17543 24055
rect 18337 24021 18371 24055
rect 18429 24021 18463 24055
rect 22477 24021 22511 24055
rect 22569 24021 22603 24055
rect 23213 24021 23247 24055
rect 23765 24021 23799 24055
rect 25237 24021 25271 24055
rect 2697 23817 2731 23851
rect 4261 23817 4295 23851
rect 4813 23817 4847 23851
rect 4997 23817 5031 23851
rect 6469 23817 6503 23851
rect 16129 23817 16163 23851
rect 19993 23817 20027 23851
rect 20545 23817 20579 23851
rect 23857 23817 23891 23851
rect 24501 23817 24535 23851
rect 2237 23749 2271 23783
rect 20821 23681 20855 23715
rect 21649 23681 21683 23715
rect 857 23613 891 23647
rect 2605 23613 2639 23647
rect 2881 23613 2915 23647
rect 4077 23613 4111 23647
rect 4169 23613 4203 23647
rect 5365 23613 5399 23647
rect 6193 23613 6227 23647
rect 6469 23613 6503 23647
rect 9137 23613 9171 23647
rect 9321 23613 9355 23647
rect 9413 23613 9447 23647
rect 12357 23613 12391 23647
rect 12549 23615 12583 23649
rect 14013 23613 14047 23647
rect 17509 23613 17543 23647
rect 17602 23613 17636 23647
rect 17785 23613 17819 23647
rect 18015 23613 18049 23647
rect 20913 23613 20947 23647
rect 21833 23613 21867 23647
rect 22201 23613 22235 23647
rect 22385 23613 22419 23647
rect 22569 23613 22603 23647
rect 22937 23613 22971 23647
rect 24041 23613 24075 23647
rect 24133 23613 24167 23647
rect 24409 23613 24443 23647
rect 24685 23613 24719 23647
rect 1124 23545 1158 23579
rect 6285 23545 6319 23579
rect 17417 23545 17451 23579
rect 17877 23545 17911 23579
rect 18705 23545 18739 23579
rect 22753 23545 22787 23579
rect 22845 23545 22879 23579
rect 24225 23545 24259 23579
rect 2421 23477 2455 23511
rect 3893 23477 3927 23511
rect 4629 23477 4663 23511
rect 4997 23477 5031 23511
rect 8953 23477 8987 23511
rect 9597 23477 9631 23511
rect 12541 23477 12575 23511
rect 14197 23477 14231 23511
rect 18153 23477 18187 23511
rect 22477 23477 22511 23511
rect 23121 23477 23155 23511
rect 1133 23273 1167 23307
rect 3433 23273 3467 23307
rect 3525 23273 3559 23307
rect 8861 23273 8895 23307
rect 9153 23273 9187 23307
rect 9321 23273 9355 23307
rect 10793 23273 10827 23307
rect 13093 23273 13127 23307
rect 13829 23273 13863 23307
rect 17325 23273 17359 23307
rect 18429 23273 18463 23307
rect 21557 23273 21591 23307
rect 21649 23273 21683 23307
rect 1777 23205 1811 23239
rect 1993 23205 2027 23239
rect 3065 23205 3099 23239
rect 3265 23205 3299 23239
rect 8953 23205 8987 23239
rect 9680 23205 9714 23239
rect 11136 23205 11170 23239
rect 13921 23205 13955 23239
rect 14933 23205 14967 23239
rect 15117 23205 15151 23239
rect 18061 23205 18095 23239
rect 19533 23205 19567 23239
rect 3709 23137 3743 23171
rect 4445 23137 4479 23171
rect 4629 23137 4663 23171
rect 6653 23137 6687 23171
rect 8401 23137 8435 23171
rect 8677 23137 8711 23171
rect 8861 23137 8895 23171
rect 9413 23137 9447 23171
rect 11253 23137 11287 23171
rect 11897 23137 11931 23171
rect 12045 23137 12079 23171
rect 12173 23137 12207 23171
rect 12265 23137 12299 23171
rect 12401 23137 12435 23171
rect 12633 23137 12667 23171
rect 12902 23137 12936 23171
rect 13191 23137 13225 23171
rect 13369 23137 13403 23171
rect 13553 23137 13587 23171
rect 14381 23137 14415 23171
rect 14565 23137 14599 23171
rect 14841 23137 14875 23171
rect 15393 23137 15427 23171
rect 15945 23137 15979 23171
rect 16773 23137 16807 23171
rect 16866 23137 16900 23171
rect 17141 23137 17175 23171
rect 17233 23137 17267 23171
rect 17785 23137 17819 23171
rect 17877 23137 17911 23171
rect 18567 23137 18601 23171
rect 18705 23137 18739 23171
rect 18797 23137 18831 23171
rect 18925 23137 18959 23171
rect 19073 23137 19107 23171
rect 19625 23137 19659 23171
rect 21465 23137 21499 23171
rect 1593 23069 1627 23103
rect 6745 23069 6779 23103
rect 8309 23069 8343 23103
rect 11345 23069 11379 23103
rect 11621 23069 11655 23103
rect 12817 23069 12851 23103
rect 16589 23069 16623 23103
rect 1317 23001 1351 23035
rect 2145 23001 2179 23035
rect 7021 23001 7055 23035
rect 12541 23001 12575 23035
rect 13185 23001 13219 23035
rect 14197 23001 14231 23035
rect 17049 23001 17083 23035
rect 21281 23001 21315 23035
rect 1961 22933 1995 22967
rect 3249 22933 3283 22967
rect 4537 22933 4571 22967
rect 9137 22933 9171 22967
rect 10977 22933 11011 22967
rect 12909 22933 12943 22967
rect 13645 22933 13679 22967
rect 13737 22933 13771 22967
rect 14749 22933 14783 22967
rect 15117 22933 15151 22967
rect 15853 22933 15887 22967
rect 17601 22933 17635 22967
rect 18061 22933 18095 22967
rect 21833 22933 21867 22967
rect 2145 22729 2179 22763
rect 3249 22729 3283 22763
rect 3801 22729 3835 22763
rect 6377 22729 6411 22763
rect 7941 22729 7975 22763
rect 11253 22729 11287 22763
rect 12173 22729 12207 22763
rect 12541 22729 12575 22763
rect 12909 22729 12943 22763
rect 13829 22729 13863 22763
rect 16405 22729 16439 22763
rect 18705 22729 18739 22763
rect 20177 22729 20211 22763
rect 2329 22661 2363 22695
rect 5365 22661 5399 22695
rect 6837 22661 6871 22695
rect 7757 22661 7791 22695
rect 13921 22661 13955 22695
rect 16221 22661 16255 22695
rect 20085 22661 20119 22695
rect 20269 22661 20303 22695
rect 21189 22661 21223 22695
rect 4721 22593 4755 22627
rect 5549 22593 5583 22627
rect 6469 22593 6503 22627
rect 8677 22593 8711 22627
rect 8769 22593 8803 22627
rect 15577 22593 15611 22627
rect 15853 22593 15887 22627
rect 19165 22593 19199 22627
rect 20637 22593 20671 22627
rect 22385 22593 22419 22627
rect 22477 22593 22511 22627
rect 23305 22593 23339 22627
rect 23857 22593 23891 22627
rect 1777 22525 1811 22559
rect 1961 22525 1995 22559
rect 2237 22525 2271 22559
rect 2421 22525 2455 22559
rect 3433 22525 3467 22559
rect 3709 22525 3743 22559
rect 3801 22525 3835 22559
rect 3893 22525 3927 22559
rect 4813 22525 4847 22559
rect 4997 22525 5031 22559
rect 5089 22525 5123 22559
rect 5181 22525 5215 22559
rect 5457 22525 5491 22559
rect 5641 22525 5675 22559
rect 5825 22525 5859 22559
rect 6193 22525 6227 22559
rect 6653 22525 6687 22559
rect 7665 22525 7699 22559
rect 8493 22525 8527 22559
rect 8585 22525 8619 22559
rect 10977 22525 11011 22559
rect 11161 22525 11195 22559
rect 11253 22525 11287 22559
rect 11805 22525 11839 22559
rect 11989 22525 12023 22559
rect 12817 22525 12851 22559
rect 12909 22525 12943 22559
rect 14013 22525 14047 22559
rect 14105 22525 14139 22559
rect 15485 22525 15519 22559
rect 19073 22525 19107 22559
rect 19969 22525 20003 22559
rect 20386 22525 20420 22559
rect 21005 22525 21039 22559
rect 21373 22525 21407 22559
rect 21557 22525 21591 22559
rect 22293 22525 22327 22559
rect 22569 22525 22603 22559
rect 23489 22525 23523 22559
rect 3617 22457 3651 22491
rect 4077 22457 4111 22491
rect 4353 22457 4387 22491
rect 4537 22457 4571 22491
rect 6377 22457 6411 22491
rect 7573 22457 7607 22491
rect 7941 22457 7975 22491
rect 13737 22457 13771 22491
rect 16589 22457 16623 22491
rect 20729 22457 20763 22491
rect 24124 22457 24158 22491
rect 5917 22389 5951 22423
rect 6009 22389 6043 22423
rect 6193 22389 6227 22423
rect 8953 22389 8987 22423
rect 14289 22389 14323 22423
rect 16389 22389 16423 22423
rect 20821 22389 20855 22423
rect 21465 22389 21499 22423
rect 22109 22389 22143 22423
rect 23673 22389 23707 22423
rect 25237 22389 25271 22423
rect 4813 22185 4847 22219
rect 24317 22185 24351 22219
rect 4445 22117 4479 22151
rect 10609 22117 10643 22151
rect 10793 22117 10827 22151
rect 13369 22117 13403 22151
rect 13553 22117 13587 22151
rect 13737 22117 13771 22151
rect 19042 22117 19076 22151
rect 20637 22117 20671 22151
rect 21741 22117 21775 22151
rect 1501 22049 1535 22083
rect 1593 22049 1627 22083
rect 1777 22049 1811 22083
rect 4629 22049 4663 22083
rect 7113 22049 7147 22083
rect 8493 22049 8527 22083
rect 8677 22049 8711 22083
rect 9321 22049 9355 22083
rect 9413 22049 9447 22083
rect 9597 22049 9631 22083
rect 10517 22049 10551 22083
rect 10977 22049 11011 22083
rect 11161 22049 11195 22083
rect 11253 22049 11287 22083
rect 11345 22049 11379 22083
rect 16405 22049 16439 22083
rect 20361 22049 20395 22083
rect 20453 22049 20487 22083
rect 21649 22049 21683 22083
rect 22017 22049 22051 22083
rect 22385 22049 22419 22083
rect 22569 22049 22603 22083
rect 22661 22049 22695 22083
rect 22845 22049 22879 22083
rect 22937 22049 22971 22083
rect 23121 22049 23155 22083
rect 23305 22049 23339 22083
rect 23393 22049 23427 22083
rect 23489 22049 23523 22083
rect 24501 22049 24535 22083
rect 2605 21981 2639 22015
rect 11621 21981 11655 22015
rect 16497 21981 16531 22015
rect 18797 21981 18831 22015
rect 22109 21981 22143 22015
rect 9597 21913 9631 21947
rect 10793 21913 10827 21947
rect 20637 21913 20671 21947
rect 22293 21913 22327 21947
rect 23673 21913 23707 21947
rect 1777 21845 1811 21879
rect 2053 21845 2087 21879
rect 6929 21845 6963 21879
rect 8309 21845 8343 21879
rect 8493 21845 8527 21879
rect 16773 21845 16807 21879
rect 20177 21845 20211 21879
rect 2421 21641 2455 21675
rect 5457 21641 5491 21675
rect 8585 21641 8619 21675
rect 9413 21641 9447 21675
rect 14197 21641 14231 21675
rect 16221 21641 16255 21675
rect 19165 21641 19199 21675
rect 21281 21641 21315 21675
rect 22017 21641 22051 21675
rect 23213 21641 23247 21675
rect 3065 21573 3099 21607
rect 8401 21573 8435 21607
rect 11897 21573 11931 21607
rect 16405 21573 16439 21607
rect 17417 21573 17451 21607
rect 24041 21573 24075 21607
rect 5549 21505 5583 21539
rect 14381 21505 14415 21539
rect 17693 21505 17727 21539
rect 20913 21505 20947 21539
rect 22385 21505 22419 21539
rect 23305 21505 23339 21539
rect 23857 21505 23891 21539
rect 1041 21437 1075 21471
rect 1308 21437 1342 21471
rect 2789 21437 2823 21471
rect 3249 21437 3283 21471
rect 4997 21437 5031 21471
rect 5273 21437 5307 21471
rect 5457 21437 5491 21471
rect 7113 21437 7147 21471
rect 7205 21437 7239 21471
rect 7481 21437 7515 21471
rect 7757 21437 7791 21471
rect 7849 21437 7883 21471
rect 8585 21437 8619 21471
rect 8953 21437 8987 21471
rect 9551 21437 9585 21471
rect 9964 21437 9998 21471
rect 10057 21437 10091 21471
rect 10333 21437 10367 21471
rect 10517 21437 10551 21471
rect 11805 21437 11839 21471
rect 11989 21437 12023 21471
rect 14013 21437 14047 21471
rect 14197 21437 14231 21471
rect 16129 21437 16163 21471
rect 16313 21437 16347 21471
rect 16589 21437 16623 21471
rect 17233 21437 17267 21471
rect 17785 21437 17819 21471
rect 18061 21437 18095 21471
rect 18245 21437 18279 21471
rect 18981 21437 19015 21471
rect 20821 21437 20855 21471
rect 21097 21437 21131 21471
rect 21373 21437 21407 21471
rect 21557 21437 21591 21471
rect 22201 21437 22235 21471
rect 23397 21437 23431 21471
rect 24133 21437 24167 21471
rect 3065 21369 3099 21403
rect 3494 21369 3528 21403
rect 5816 21369 5850 21403
rect 9689 21369 9723 21403
rect 9781 21369 9815 21403
rect 10425 21369 10459 21403
rect 14648 21369 14682 21403
rect 16681 21369 16715 21403
rect 18153 21369 18187 21403
rect 2881 21301 2915 21335
rect 4629 21301 4663 21335
rect 4813 21301 4847 21335
rect 6929 21301 6963 21335
rect 15761 21301 15795 21335
rect 15853 21301 15887 21335
rect 21649 21301 21683 21335
rect 23029 21301 23063 21335
rect 23857 21301 23891 21335
rect 1777 21097 1811 21131
rect 3249 21097 3283 21131
rect 9137 21097 9171 21131
rect 14841 21097 14875 21131
rect 18797 21097 18831 21131
rect 19257 21097 19291 21131
rect 22753 21097 22787 21131
rect 9689 21029 9723 21063
rect 10425 21029 10459 21063
rect 11161 21029 11195 21063
rect 11989 21029 12023 21063
rect 16748 21029 16782 21063
rect 17417 21029 17451 21063
rect 19441 21029 19475 21063
rect 19901 21029 19935 21063
rect 19994 21029 20028 21063
rect 2053 20961 2087 20995
rect 3525 20961 3559 20995
rect 4997 20961 5031 20995
rect 5273 20961 5307 20995
rect 5365 20961 5399 20995
rect 5825 20961 5859 20995
rect 7573 20961 7607 20995
rect 7849 20961 7883 20995
rect 11805 20961 11839 20995
rect 12081 20961 12115 20995
rect 12541 20961 12575 20995
rect 12808 20961 12842 20995
rect 14197 20961 14231 20995
rect 14381 20961 14415 20995
rect 15025 20961 15059 20995
rect 15209 20961 15243 20995
rect 17325 20961 17359 20995
rect 17509 20961 17543 20995
rect 19165 20961 19199 20995
rect 19809 20961 19843 20995
rect 20111 20961 20145 20995
rect 20269 20961 20303 20995
rect 21833 20961 21867 20995
rect 22017 20961 22051 20995
rect 23121 20961 23155 20995
rect 23213 20961 23247 20995
rect 1777 20893 1811 20927
rect 3249 20893 3283 20927
rect 5181 20893 5215 20927
rect 5549 20893 5583 20927
rect 9873 20893 9907 20927
rect 9965 20893 9999 20927
rect 15301 20893 15335 20927
rect 16865 20893 16899 20927
rect 16957 20893 16991 20927
rect 17233 20893 17267 20927
rect 18337 20893 18371 20927
rect 18889 20893 18923 20927
rect 19073 20893 19107 20927
rect 19533 20893 19567 20927
rect 3433 20825 3467 20859
rect 4813 20825 4847 20859
rect 10425 20825 10459 20859
rect 10977 20825 11011 20859
rect 11529 20825 11563 20859
rect 13921 20825 13955 20859
rect 16589 20825 16623 20859
rect 18705 20825 18739 20859
rect 19625 20825 19659 20859
rect 1961 20757 1995 20791
rect 5457 20757 5491 20791
rect 11161 20757 11195 20791
rect 11621 20757 11655 20791
rect 14013 20757 14047 20791
rect 14381 20757 14415 20791
rect 21833 20757 21867 20791
rect 23397 20757 23431 20791
rect 5825 20553 5859 20587
rect 8769 20553 8803 20587
rect 9413 20553 9447 20587
rect 9505 20553 9539 20587
rect 11805 20553 11839 20587
rect 12817 20553 12851 20587
rect 16313 20553 16347 20587
rect 20177 20553 20211 20587
rect 20913 20553 20947 20587
rect 22201 20553 22235 20587
rect 6745 20485 6779 20519
rect 8401 20417 8435 20451
rect 9597 20417 9631 20451
rect 13829 20417 13863 20451
rect 15393 20417 15427 20451
rect 16773 20417 16807 20451
rect 16957 20417 16991 20451
rect 20453 20417 20487 20451
rect 20637 20417 20671 20451
rect 20821 20417 20855 20451
rect 22385 20417 22419 20451
rect 1777 20349 1811 20383
rect 5825 20349 5859 20383
rect 6009 20349 6043 20383
rect 6929 20349 6963 20383
rect 7113 20349 7147 20383
rect 8585 20349 8619 20383
rect 9045 20349 9079 20383
rect 9229 20349 9263 20383
rect 9321 20349 9355 20383
rect 11161 20349 11195 20383
rect 11989 20349 12023 20383
rect 12357 20349 12391 20383
rect 13093 20349 13127 20383
rect 13553 20349 13587 20383
rect 13645 20349 13679 20383
rect 18705 20349 18739 20383
rect 20361 20349 20395 20383
rect 20545 20349 20579 20383
rect 21005 20349 21039 20383
rect 21097 20349 21131 20383
rect 21649 20349 21683 20383
rect 21741 20349 21775 20383
rect 22109 20349 22143 20383
rect 22477 20349 22511 20383
rect 22845 20349 22879 20383
rect 7297 20281 7331 20315
rect 12081 20281 12115 20315
rect 12173 20281 12207 20315
rect 12817 20281 12851 20315
rect 13829 20281 13863 20315
rect 18337 20281 18371 20315
rect 18797 20281 18831 20315
rect 21465 20281 21499 20315
rect 22385 20281 22419 20315
rect 22661 20281 22695 20315
rect 22753 20281 22787 20315
rect 1593 20213 1627 20247
rect 7021 20213 7055 20247
rect 8953 20213 8987 20247
rect 11345 20213 11379 20247
rect 13001 20213 13035 20247
rect 14841 20213 14875 20247
rect 16681 20213 16715 20247
rect 18061 20213 18095 20247
rect 23029 20213 23063 20247
rect 4353 20009 4387 20043
rect 4813 20009 4847 20043
rect 6653 20009 6687 20043
rect 7113 20009 7147 20043
rect 7297 20009 7331 20043
rect 7573 20009 7607 20043
rect 8401 20009 8435 20043
rect 12357 20009 12391 20043
rect 13553 20009 13587 20043
rect 13645 20009 13679 20043
rect 13813 20009 13847 20043
rect 15485 20009 15519 20043
rect 16681 20009 16715 20043
rect 17233 20009 17267 20043
rect 20729 20009 20763 20043
rect 21465 20009 21499 20043
rect 22109 20009 22143 20043
rect 24317 20009 24351 20043
rect 1584 19941 1618 19975
rect 3141 19941 3175 19975
rect 3341 19941 3375 19975
rect 6469 19941 6503 19975
rect 7408 19941 7442 19975
rect 11244 19941 11278 19975
rect 14013 19941 14047 19975
rect 21925 19941 21959 19975
rect 1317 19873 1351 19907
rect 5181 19873 5215 19907
rect 6101 19873 6135 19907
rect 6745 19873 6779 19907
rect 7205 19873 7239 19907
rect 8033 19873 8067 19907
rect 8217 19873 8251 19907
rect 9965 19873 9999 19907
rect 10057 19873 10091 19907
rect 13093 19873 13127 19907
rect 13185 19873 13219 19907
rect 14105 19873 14139 19907
rect 14361 19873 14395 19907
rect 16221 19873 16255 19907
rect 16773 19873 16807 19907
rect 18889 19873 18923 19907
rect 19533 19873 19567 19907
rect 20913 19873 20947 19907
rect 21097 19873 21131 19907
rect 21281 19873 21315 19907
rect 21557 19873 21591 19907
rect 21741 19873 21775 19907
rect 23204 19873 23238 19907
rect 4997 19805 5031 19839
rect 5089 19805 5123 19839
rect 5273 19805 5307 19839
rect 6837 19805 6871 19839
rect 7573 19805 7607 19839
rect 10977 19805 11011 19839
rect 13277 19805 13311 19839
rect 20085 19805 20119 19839
rect 22937 19805 22971 19839
rect 2973 19737 3007 19771
rect 3985 19737 4019 19771
rect 2697 19669 2731 19703
rect 3157 19669 3191 19703
rect 4353 19669 4387 19703
rect 4537 19669 4571 19703
rect 6469 19669 6503 19703
rect 6837 19669 6871 19703
rect 10149 19669 10183 19703
rect 10333 19669 10367 19703
rect 13001 19669 13035 19703
rect 13277 19669 13311 19703
rect 13829 19669 13863 19703
rect 16313 19669 16347 19703
rect 16865 19669 16899 19703
rect 18797 19669 18831 19703
rect 21281 19669 21315 19703
rect 1777 19465 1811 19499
rect 1961 19465 1995 19499
rect 5549 19465 5583 19499
rect 6101 19465 6135 19499
rect 6929 19465 6963 19499
rect 16037 19465 16071 19499
rect 20085 19465 20119 19499
rect 20545 19465 20579 19499
rect 21833 19465 21867 19499
rect 23213 19465 23247 19499
rect 1409 19397 1443 19431
rect 9689 19397 9723 19431
rect 10057 19397 10091 19431
rect 13093 19397 13127 19431
rect 14013 19397 14047 19431
rect 20729 19397 20763 19431
rect 3617 19329 3651 19363
rect 3709 19329 3743 19363
rect 8677 19329 8711 19363
rect 9505 19329 9539 19363
rect 15761 19329 15795 19363
rect 20637 19329 20671 19363
rect 22201 19329 22235 19363
rect 2421 19261 2455 19295
rect 2605 19261 2639 19295
rect 3433 19261 3467 19295
rect 3893 19261 3927 19295
rect 3985 19261 4019 19295
rect 4169 19261 4203 19295
rect 6653 19261 6687 19295
rect 6929 19261 6963 19295
rect 8769 19261 8803 19295
rect 9413 19261 9447 19295
rect 9873 19261 9907 19295
rect 10149 19261 10183 19295
rect 10333 19261 10367 19295
rect 10425 19261 10459 19295
rect 11713 19261 11747 19295
rect 15669 19261 15703 19295
rect 17969 19261 18003 19295
rect 18061 19261 18095 19295
rect 18245 19261 18279 19295
rect 18337 19261 18371 19295
rect 18705 19261 18739 19295
rect 21005 19261 21039 19295
rect 22109 19261 22143 19295
rect 22293 19261 22327 19295
rect 22569 19261 22603 19295
rect 22753 19261 22787 19295
rect 22937 19261 22971 19295
rect 23397 19261 23431 19295
rect 1777 19193 1811 19227
rect 2697 19193 2731 19227
rect 2881 19193 2915 19227
rect 3065 19193 3099 19227
rect 3249 19193 3283 19227
rect 3709 19193 3743 19227
rect 4436 19193 4470 19227
rect 6285 19193 6319 19227
rect 6745 19193 6779 19227
rect 11980 19193 12014 19227
rect 15301 19193 15335 19227
rect 18972 19193 19006 19227
rect 21817 19193 21851 19227
rect 22017 19193 22051 19227
rect 2513 19125 2547 19159
rect 5917 19125 5951 19159
rect 6085 19125 6119 19159
rect 8401 19125 8435 19159
rect 9045 19125 9079 19159
rect 18521 19125 18555 19159
rect 20269 19125 20303 19159
rect 20913 19125 20947 19159
rect 21649 19125 21683 19159
rect 4169 18921 4203 18955
rect 4905 18921 4939 18955
rect 11805 18921 11839 18955
rect 11989 18921 12023 18955
rect 14289 18921 14323 18955
rect 18711 18921 18745 18955
rect 18797 18921 18831 18955
rect 8861 18853 8895 18887
rect 9045 18853 9079 18887
rect 13185 18853 13219 18887
rect 18613 18853 18647 18887
rect 20361 18853 20395 18887
rect 20729 18853 20763 18887
rect 23581 18853 23615 18887
rect 3617 18785 3651 18819
rect 4445 18785 4479 18819
rect 5089 18785 5123 18819
rect 6745 18785 6779 18819
rect 8769 18785 8803 18819
rect 10977 18785 11011 18819
rect 11621 18785 11655 18819
rect 11713 18785 11747 18819
rect 11897 18785 11931 18819
rect 12173 18785 12207 18819
rect 13645 18785 13679 18819
rect 13829 18785 13863 18819
rect 13921 18785 13955 18819
rect 14013 18785 14047 18819
rect 16865 18785 16899 18819
rect 17325 18785 17359 18819
rect 17509 18785 17543 18819
rect 17601 18785 17635 18819
rect 18889 18785 18923 18819
rect 20269 18785 20303 18819
rect 20913 18785 20947 18819
rect 21005 18785 21039 18819
rect 22017 18785 22051 18819
rect 23857 18785 23891 18819
rect 6837 18717 6871 18751
rect 16957 18717 16991 18751
rect 17233 18717 17267 18751
rect 20453 18717 20487 18751
rect 20729 18717 20763 18751
rect 4537 18581 4571 18615
rect 7021 18581 7055 18615
rect 9045 18581 9079 18615
rect 13277 18581 13311 18615
rect 17325 18581 17359 18615
rect 19901 18581 19935 18615
rect 22201 18581 22235 18615
rect 2973 18377 3007 18411
rect 12081 18377 12115 18411
rect 12265 18377 12299 18411
rect 13207 18377 13241 18411
rect 13369 18377 13403 18411
rect 14841 18377 14875 18411
rect 17417 18377 17451 18411
rect 5365 18309 5399 18343
rect 7297 18309 7331 18343
rect 16865 18309 16899 18343
rect 4445 18241 4479 18275
rect 4905 18241 4939 18275
rect 5917 18241 5951 18275
rect 7138 18241 7172 18275
rect 7941 18241 7975 18275
rect 8769 18241 8803 18275
rect 8953 18241 8987 18275
rect 16773 18241 16807 18275
rect 1593 18173 1627 18207
rect 1860 18173 1894 18207
rect 4353 18173 4387 18207
rect 4997 18173 5031 18207
rect 6285 18173 6319 18207
rect 6653 18173 6687 18207
rect 6929 18173 6963 18207
rect 7849 18173 7883 18207
rect 8861 18173 8895 18207
rect 9045 18173 9079 18207
rect 9321 18173 9355 18207
rect 9597 18173 9631 18207
rect 9689 18173 9723 18207
rect 11713 18173 11747 18207
rect 13553 18173 13587 18207
rect 17049 18173 17083 18207
rect 17233 18173 17267 18207
rect 17325 18173 17359 18207
rect 17509 18173 17543 18207
rect 19533 18173 19567 18207
rect 19717 18173 19751 18207
rect 6193 18105 6227 18139
rect 6469 18105 6503 18139
rect 9505 18105 9539 18139
rect 12541 18105 12575 18139
rect 12725 18105 12759 18139
rect 13001 18105 13035 18139
rect 13201 18105 13235 18139
rect 16506 18105 16540 18139
rect 4721 18037 4755 18071
rect 6101 18037 6135 18071
rect 7021 18037 7055 18071
rect 8217 18037 8251 18071
rect 9229 18037 9263 18071
rect 9873 18037 9907 18071
rect 12081 18037 12115 18071
rect 12357 18037 12391 18071
rect 15393 18037 15427 18071
rect 19625 18037 19659 18071
rect 7205 17833 7239 17867
rect 8953 17833 8987 17867
rect 10977 17833 11011 17867
rect 14105 17833 14139 17867
rect 14381 17833 14415 17867
rect 19073 17833 19107 17867
rect 21005 17833 21039 17867
rect 10548 17765 10582 17799
rect 19870 17765 19904 17799
rect 3240 17697 3274 17731
rect 5917 17697 5951 17731
rect 6009 17697 6043 17731
rect 6377 17697 6411 17731
rect 7297 17697 7331 17731
rect 8309 17697 8343 17731
rect 8769 17697 8803 17731
rect 11161 17697 11195 17731
rect 11713 17697 11747 17731
rect 11989 17697 12023 17731
rect 12173 17697 12207 17731
rect 12357 17697 12391 17731
rect 13369 17697 13403 17731
rect 13461 17697 13495 17731
rect 13737 17697 13771 17731
rect 14749 17697 14783 17731
rect 14841 17697 14875 17731
rect 15025 17697 15059 17731
rect 16129 17697 16163 17731
rect 16681 17697 16715 17731
rect 17693 17697 17727 17731
rect 17949 17697 17983 17731
rect 19625 17697 19659 17731
rect 2973 17629 3007 17663
rect 8585 17629 8619 17663
rect 10793 17629 10827 17663
rect 13001 17629 13035 17663
rect 13277 17629 13311 17663
rect 13553 17629 13587 17663
rect 14565 17629 14599 17663
rect 14657 17629 14691 17663
rect 6561 17561 6595 17595
rect 9413 17561 9447 17595
rect 13093 17561 13127 17595
rect 14289 17561 14323 17595
rect 15209 17561 15243 17595
rect 4353 17493 4387 17527
rect 6285 17493 6319 17527
rect 8769 17493 8803 17527
rect 11529 17493 11563 17527
rect 14105 17493 14139 17527
rect 3709 17289 3743 17323
rect 8953 17289 8987 17323
rect 9873 17289 9907 17323
rect 10057 17289 10091 17323
rect 12541 17289 12575 17323
rect 13185 17289 13219 17323
rect 13369 17289 13403 17323
rect 16129 17289 16163 17323
rect 17049 17289 17083 17323
rect 12909 17153 12943 17187
rect 14105 17153 14139 17187
rect 14381 17153 14415 17187
rect 15301 17153 15335 17187
rect 16589 17153 16623 17187
rect 17785 17153 17819 17187
rect 18153 17153 18187 17187
rect 18245 17153 18279 17187
rect 18981 17153 19015 17187
rect 3341 17085 3375 17119
rect 3433 17085 3467 17119
rect 3617 17085 3651 17119
rect 3893 17085 3927 17119
rect 12725 17085 12759 17119
rect 14013 17085 14047 17119
rect 15209 17085 15243 17119
rect 15393 17085 15427 17119
rect 15485 17085 15519 17119
rect 15578 17085 15612 17119
rect 15761 17085 15795 17119
rect 15950 17085 15984 17119
rect 17325 17085 17359 17119
rect 17417 17085 17451 17119
rect 17509 17085 17543 17119
rect 17693 17085 17727 17119
rect 17969 17085 18003 17119
rect 18061 17085 18095 17119
rect 19073 17085 19107 17119
rect 20361 17085 20395 17119
rect 8401 17017 8435 17051
rect 9689 17017 9723 17051
rect 13001 17017 13035 17051
rect 15853 17017 15887 17051
rect 16221 17017 16255 17051
rect 16405 17017 16439 17051
rect 8585 16949 8619 16983
rect 8677 16949 8711 16983
rect 8769 16949 8803 16983
rect 9889 16949 9923 16983
rect 13211 16949 13245 16983
rect 18705 16949 18739 16983
rect 20453 16949 20487 16983
rect 4169 16745 4203 16779
rect 7941 16745 7975 16779
rect 9781 16745 9815 16779
rect 12541 16745 12575 16779
rect 15393 16745 15427 16779
rect 17509 16745 17543 16779
rect 17601 16745 17635 16779
rect 4445 16677 4479 16711
rect 6285 16677 6319 16711
rect 6377 16677 6411 16711
rect 11428 16677 11462 16711
rect 15025 16677 15059 16711
rect 15241 16677 15275 16711
rect 17785 16677 17819 16711
rect 18597 16677 18631 16711
rect 18797 16677 18831 16711
rect 2145 16609 2179 16643
rect 4353 16609 4387 16643
rect 4537 16609 4571 16643
rect 4721 16609 4755 16643
rect 5273 16609 5307 16643
rect 6101 16609 6135 16643
rect 6489 16631 6523 16665
rect 6653 16609 6687 16643
rect 6745 16609 6779 16643
rect 6929 16609 6963 16643
rect 7113 16609 7147 16643
rect 7205 16609 7239 16643
rect 7389 16609 7423 16643
rect 7757 16609 7791 16643
rect 9045 16609 9079 16643
rect 9597 16609 9631 16643
rect 9781 16609 9815 16643
rect 10149 16609 10183 16643
rect 11161 16609 11195 16643
rect 12817 16609 12851 16643
rect 15761 16609 15795 16643
rect 15945 16609 15979 16643
rect 16865 16609 16899 16643
rect 17350 16609 17384 16643
rect 18153 16609 18187 16643
rect 19993 16609 20027 16643
rect 20177 16609 20211 16643
rect 5365 16541 5399 16575
rect 7481 16541 7515 16575
rect 7573 16541 7607 16575
rect 8033 16541 8067 16575
rect 13093 16541 13127 16575
rect 17141 16541 17175 16575
rect 17233 16541 17267 16575
rect 5641 16473 5675 16507
rect 6101 16473 6135 16507
rect 12909 16473 12943 16507
rect 1961 16405 1995 16439
rect 10333 16405 10367 16439
rect 13001 16405 13035 16439
rect 15209 16405 15243 16439
rect 15945 16405 15979 16439
rect 17785 16405 17819 16439
rect 18429 16405 18463 16439
rect 18613 16405 18647 16439
rect 20085 16405 20119 16439
rect 3709 16201 3743 16235
rect 6837 16201 6871 16235
rect 7297 16201 7331 16235
rect 9413 16201 9447 16235
rect 15301 16201 15335 16235
rect 16773 16201 16807 16235
rect 17509 16201 17543 16235
rect 17969 16201 18003 16235
rect 19993 16201 20027 16235
rect 2881 16133 2915 16167
rect 14381 16133 14415 16167
rect 15761 16133 15795 16167
rect 20545 16133 20579 16167
rect 3341 16065 3375 16099
rect 11805 16065 11839 16099
rect 14105 16065 14139 16099
rect 21925 16065 21959 16099
rect 1501 15997 1535 16031
rect 1768 15997 1802 16031
rect 3433 15997 3467 16031
rect 4445 15997 4479 16031
rect 4537 15997 4571 16031
rect 4813 15997 4847 16031
rect 6653 15997 6687 16031
rect 7205 15997 7239 16031
rect 7389 15997 7423 16031
rect 8861 15997 8895 16031
rect 8953 15997 8987 16031
rect 9137 15997 9171 16031
rect 9229 15997 9263 16031
rect 10986 15997 11020 16031
rect 11253 15997 11287 16031
rect 11621 15997 11655 16031
rect 12909 15997 12943 16031
rect 13093 15997 13127 16031
rect 13185 15997 13219 16031
rect 13737 15997 13771 16031
rect 14013 15997 14047 16031
rect 15117 15997 15151 16031
rect 15209 15997 15243 16031
rect 15485 15997 15519 16031
rect 15761 15997 15795 16031
rect 17049 15997 17083 16031
rect 17141 15997 17175 16031
rect 17233 15997 17267 16031
rect 17393 15997 17427 16031
rect 17675 15997 17709 16031
rect 17877 15997 17911 16031
rect 18705 15997 18739 16031
rect 4629 15929 4663 15963
rect 6745 15929 6779 15963
rect 6929 15929 6963 15963
rect 15393 15929 15427 15963
rect 18153 15929 18187 15963
rect 21658 15929 21692 15963
rect 4261 15861 4295 15895
rect 9873 15861 9907 15895
rect 11437 15861 11471 15895
rect 12725 15861 12759 15895
rect 13645 15861 13679 15895
rect 15577 15861 15611 15895
rect 2145 15657 2179 15691
rect 6653 15657 6687 15691
rect 13277 15657 13311 15691
rect 17601 15657 17635 15691
rect 20177 15657 20211 15691
rect 6193 15589 6227 15623
rect 2329 15521 2363 15555
rect 5089 15521 5123 15555
rect 6091 15521 6125 15555
rect 6285 15521 6319 15555
rect 6561 15521 6595 15555
rect 6745 15521 6779 15555
rect 9045 15521 9079 15555
rect 13461 15521 13495 15555
rect 13553 15521 13587 15555
rect 16957 15521 16991 15555
rect 17050 15521 17084 15555
rect 17233 15521 17267 15555
rect 17325 15521 17359 15555
rect 17422 15521 17456 15555
rect 17969 15521 18003 15555
rect 19073 15521 19107 15555
rect 19533 15521 19567 15555
rect 19717 15521 19751 15555
rect 19809 15521 19843 15555
rect 19901 15521 19935 15555
rect 20269 15521 20303 15555
rect 20637 15521 20671 15555
rect 20913 15521 20947 15555
rect 21281 15521 21315 15555
rect 22762 15521 22796 15555
rect 23029 15521 23063 15555
rect 2513 15453 2547 15487
rect 5181 15453 5215 15487
rect 8585 15453 8619 15487
rect 8953 15453 8987 15487
rect 13277 15453 13311 15487
rect 17693 15453 17727 15487
rect 18705 15453 18739 15487
rect 18981 15453 19015 15487
rect 20453 15453 20487 15487
rect 21005 15453 21039 15487
rect 4721 15385 4755 15419
rect 17785 15385 17819 15419
rect 21465 15385 21499 15419
rect 9229 15317 9263 15351
rect 17877 15317 17911 15351
rect 20361 15317 20395 15351
rect 21649 15317 21683 15351
rect 7481 15113 7515 15147
rect 8677 15113 8711 15147
rect 8861 15113 8895 15147
rect 12081 15113 12115 15147
rect 19993 15113 20027 15147
rect 21649 15113 21683 15147
rect 2421 15045 2455 15079
rect 2973 15045 3007 15079
rect 3065 15045 3099 15079
rect 7297 15045 7331 15079
rect 9229 15045 9263 15079
rect 10517 15045 10551 15079
rect 16037 15045 16071 15079
rect 21557 15045 21591 15079
rect 2053 14977 2087 15011
rect 2513 14977 2547 15011
rect 3617 14977 3651 15011
rect 4169 14977 4203 15011
rect 9781 14977 9815 15011
rect 10057 14977 10091 15011
rect 10793 14977 10827 15011
rect 11253 14977 11287 15011
rect 11621 14977 11655 15011
rect 11805 14977 11839 15011
rect 14289 14977 14323 15011
rect 15577 14977 15611 15011
rect 18889 14977 18923 15011
rect 19809 14977 19843 15011
rect 20545 14977 20579 15011
rect 2605 14909 2639 14943
rect 3249 14909 3283 14943
rect 3433 14909 3467 14943
rect 3709 14909 3743 14943
rect 3801 14909 3835 14943
rect 3893 14909 3927 14943
rect 4353 14909 4387 14943
rect 4629 14909 4663 14943
rect 4813 14909 4847 14943
rect 5917 14909 5951 14943
rect 7849 14909 7883 14943
rect 7941 14909 7975 14943
rect 8493 14909 8527 14943
rect 8677 14909 8711 14943
rect 8769 14909 8803 14943
rect 9045 14909 9079 14943
rect 9689 14909 9723 14943
rect 10241 14909 10275 14943
rect 10885 14909 10919 14943
rect 11161 14909 11195 14943
rect 11530 14909 11564 14943
rect 11713 14909 11747 14943
rect 12257 14919 12291 14953
rect 12357 14909 12391 14943
rect 12541 14909 12575 14943
rect 12633 14909 12667 14943
rect 14565 14909 14599 14943
rect 14657 14909 14691 14943
rect 14749 14909 14783 14943
rect 14933 14909 14967 14943
rect 15669 14909 15703 14943
rect 18245 14909 18279 14943
rect 18981 14909 19015 14943
rect 19901 14909 19935 14943
rect 20085 14909 20119 14943
rect 20453 14909 20487 14943
rect 21005 14909 21039 14943
rect 21189 14909 21223 14943
rect 21373 14909 21407 14943
rect 21833 14909 21867 14943
rect 21925 14909 21959 14943
rect 3341 14841 3375 14875
rect 6184 14841 6218 14875
rect 7665 14841 7699 14875
rect 10517 14841 10551 14875
rect 13829 14841 13863 14875
rect 21281 14841 21315 14875
rect 4077 14773 4111 14807
rect 8125 14773 8159 14807
rect 10333 14773 10367 14807
rect 10609 14773 10643 14807
rect 11345 14773 11379 14807
rect 13921 14773 13955 14807
rect 18337 14773 18371 14807
rect 20821 14773 20855 14807
rect 6285 14569 6319 14603
rect 12449 14569 12483 14603
rect 13921 14569 13955 14603
rect 14289 14569 14323 14603
rect 15577 14569 15611 14603
rect 16129 14569 16163 14603
rect 17325 14569 17359 14603
rect 12808 14501 12842 14535
rect 15117 14501 15151 14535
rect 15729 14501 15763 14535
rect 15945 14501 15979 14535
rect 18889 14501 18923 14535
rect 3157 14433 3191 14467
rect 3341 14433 3375 14467
rect 3433 14433 3467 14467
rect 3801 14433 3835 14467
rect 6009 14433 6043 14467
rect 6193 14433 6227 14467
rect 6469 14433 6503 14467
rect 8493 14433 8527 14467
rect 8677 14433 8711 14467
rect 10612 14433 10646 14467
rect 11336 14433 11370 14467
rect 14289 14433 14323 14467
rect 14749 14433 14783 14467
rect 14933 14433 14967 14467
rect 16313 14433 16347 14467
rect 16497 14433 16531 14467
rect 16957 14433 16991 14467
rect 21465 14433 21499 14467
rect 3709 14365 3743 14399
rect 4169 14365 4203 14399
rect 5825 14365 5859 14399
rect 8953 14365 8987 14399
rect 10425 14365 10459 14399
rect 11069 14365 11103 14399
rect 12541 14365 12575 14399
rect 14013 14365 14047 14399
rect 16865 14365 16899 14399
rect 3157 14297 3191 14331
rect 8677 14297 8711 14331
rect 14197 14297 14231 14331
rect 19165 14297 19199 14331
rect 10793 14229 10827 14263
rect 15761 14229 15795 14263
rect 19349 14229 19383 14263
rect 21649 14229 21683 14263
rect 6009 14025 6043 14059
rect 8953 14025 8987 14059
rect 11437 14025 11471 14059
rect 7113 13957 7147 13991
rect 7481 13957 7515 13991
rect 21189 13957 21223 13991
rect 6837 13889 6871 13923
rect 19165 13889 19199 13923
rect 19809 13889 19843 13923
rect 20269 13889 20303 13923
rect 2053 13821 2087 13855
rect 3985 13821 4019 13855
rect 4169 13821 4203 13855
rect 5457 13821 5491 13855
rect 5733 13821 5767 13855
rect 5825 13821 5859 13855
rect 7849 13821 7883 13855
rect 8861 13821 8895 13855
rect 11621 13821 11655 13855
rect 13645 13821 13679 13855
rect 13829 13821 13863 13855
rect 18889 13821 18923 13855
rect 19073 13821 19107 13855
rect 19349 13821 19383 13855
rect 19533 13821 19567 13855
rect 19901 13821 19935 13855
rect 20545 13821 20579 13855
rect 20729 13821 20763 13855
rect 20821 13821 20855 13855
rect 20913 13821 20947 13855
rect 22569 13821 22603 13855
rect 5641 13753 5675 13787
rect 22302 13753 22336 13787
rect 1869 13685 1903 13719
rect 4169 13685 4203 13719
rect 7297 13685 7331 13719
rect 7389 13685 7423 13719
rect 13737 13685 13771 13719
rect 18705 13685 18739 13719
rect 19441 13685 19475 13719
rect 21097 13685 21131 13719
rect 6101 13481 6135 13515
rect 10057 13481 10091 13515
rect 10609 13481 10643 13515
rect 13461 13481 13495 13515
rect 15761 13481 15795 13515
rect 19533 13481 19567 13515
rect 19809 13481 19843 13515
rect 21649 13481 21683 13515
rect 4261 13413 4295 13447
rect 4629 13413 4663 13447
rect 7573 13413 7607 13447
rect 7849 13413 7883 13447
rect 9597 13413 9631 13447
rect 11437 13413 11471 13447
rect 13737 13413 13771 13447
rect 13921 13413 13955 13447
rect 14105 13413 14139 13447
rect 14611 13413 14645 13447
rect 17794 13413 17828 13447
rect 19073 13413 19107 13447
rect 19625 13413 19659 13447
rect 1501 13345 1535 13379
rect 1768 13345 1802 13379
rect 3157 13345 3191 13379
rect 3893 13345 3927 13379
rect 4537 13345 4571 13379
rect 4721 13345 4755 13379
rect 4905 13345 4939 13379
rect 9873 13345 9907 13379
rect 10149 13345 10183 13379
rect 10241 13345 10275 13379
rect 13093 13345 13127 13379
rect 14289 13345 14323 13379
rect 14381 13345 14415 13379
rect 14473 13345 14507 13379
rect 15209 13345 15243 13379
rect 15393 13345 15427 13379
rect 15669 13345 15703 13379
rect 15853 13345 15887 13379
rect 16129 13345 16163 13379
rect 16313 13345 16347 13379
rect 18705 13345 18739 13379
rect 19901 13345 19935 13379
rect 21465 13345 21499 13379
rect 3249 13277 3283 13311
rect 4077 13277 4111 13311
rect 10333 13277 10367 13311
rect 13001 13277 13035 13311
rect 14749 13277 14783 13311
rect 18061 13277 18095 13311
rect 18613 13277 18647 13311
rect 18797 13277 18831 13311
rect 18889 13277 18923 13311
rect 21281 13277 21315 13311
rect 2881 13209 2915 13243
rect 3525 13209 3559 13243
rect 3893 13209 3927 13243
rect 19349 13209 19383 13243
rect 4353 13141 4387 13175
rect 9689 13141 9723 13175
rect 10425 13141 10459 13175
rect 11713 13141 11747 13175
rect 13553 13141 13587 13175
rect 15577 13141 15611 13175
rect 16129 13141 16163 13175
rect 16681 13141 16715 13175
rect 18429 13141 18463 13175
rect 19625 13141 19659 13175
rect 2053 12937 2087 12971
rect 5825 12937 5859 12971
rect 7665 12937 7699 12971
rect 7849 12937 7883 12971
rect 9045 12937 9079 12971
rect 10333 12937 10367 12971
rect 10793 12937 10827 12971
rect 12633 12937 12667 12971
rect 13001 12937 13035 12971
rect 13737 12937 13771 12971
rect 15025 12937 15059 12971
rect 17877 12937 17911 12971
rect 4169 12869 4203 12903
rect 7941 12869 7975 12903
rect 17325 12869 17359 12903
rect 3709 12801 3743 12835
rect 6285 12801 6319 12835
rect 7481 12801 7515 12835
rect 8769 12801 8803 12835
rect 10057 12801 10091 12835
rect 11253 12801 11287 12835
rect 16129 12801 16163 12835
rect 16405 12801 16439 12835
rect 2237 12733 2271 12767
rect 2421 12733 2455 12767
rect 3801 12733 3835 12767
rect 6193 12733 6227 12767
rect 6653 12733 6687 12767
rect 6929 12733 6963 12767
rect 7665 12733 7699 12767
rect 7941 12733 7975 12767
rect 8125 12733 8159 12767
rect 8677 12733 8711 12767
rect 9781 12733 9815 12767
rect 9965 12733 9999 12767
rect 10517 12733 10551 12767
rect 14749 12733 14783 12767
rect 15025 12733 15059 12767
rect 15117 12733 15151 12767
rect 15301 12733 15335 12767
rect 16037 12733 16071 12767
rect 16773 12733 16807 12767
rect 16957 12733 16991 12767
rect 17049 12733 17083 12767
rect 17141 12733 17175 12767
rect 17417 12733 17451 12767
rect 17601 12733 17635 12767
rect 17785 12733 17819 12767
rect 18061 12733 18095 12767
rect 6745 12665 6779 12699
rect 7205 12665 7239 12699
rect 9873 12665 9907 12699
rect 10977 12665 11011 12699
rect 11520 12665 11554 12699
rect 13185 12665 13219 12699
rect 13721 12665 13755 12699
rect 13921 12665 13955 12699
rect 14841 12665 14875 12699
rect 7113 12597 7147 12631
rect 10609 12597 10643 12631
rect 10777 12597 10811 12631
rect 12817 12597 12851 12631
rect 12985 12597 13019 12631
rect 13553 12597 13587 12631
rect 15209 12597 15243 12631
rect 4721 12393 4755 12427
rect 9229 12393 9263 12427
rect 19165 12393 19199 12427
rect 7665 12325 7699 12359
rect 19349 12325 19383 12359
rect 19809 12325 19843 12359
rect 4813 12257 4847 12291
rect 5457 12257 5491 12291
rect 5641 12267 5675 12301
rect 6101 12257 6135 12291
rect 6193 12257 6227 12291
rect 6285 12257 6319 12291
rect 6469 12257 6503 12291
rect 6653 12257 6687 12291
rect 6837 12257 6871 12291
rect 7297 12257 7331 12291
rect 7573 12257 7607 12291
rect 7849 12257 7883 12291
rect 8769 12257 8803 12291
rect 11437 12257 11471 12291
rect 11621 12257 11655 12291
rect 12081 12257 12115 12291
rect 12357 12257 12391 12291
rect 18797 12257 18831 12291
rect 19257 12257 19291 12291
rect 19625 12257 19659 12291
rect 19901 12257 19935 12291
rect 19993 12257 20027 12291
rect 20361 12257 20395 12291
rect 20453 12257 20487 12291
rect 20637 12257 20671 12291
rect 20729 12257 20763 12291
rect 6929 12189 6963 12223
rect 7205 12189 7239 12223
rect 12265 12189 12299 12223
rect 18889 12189 18923 12223
rect 5549 12121 5583 12155
rect 20177 12121 20211 12155
rect 5825 12053 5859 12087
rect 6837 12053 6871 12087
rect 8033 12053 8067 12087
rect 8953 12053 8987 12087
rect 11529 12053 11563 12087
rect 11897 12053 11931 12087
rect 20913 12053 20947 12087
rect 3801 11849 3835 11883
rect 8861 11849 8895 11883
rect 10425 11849 10459 11883
rect 7205 11781 7239 11815
rect 13093 11781 13127 11815
rect 14105 11781 14139 11815
rect 15025 11781 15059 11815
rect 18429 11781 18463 11815
rect 19809 11781 19843 11815
rect 9413 11713 9447 11747
rect 9505 11713 9539 11747
rect 10333 11713 10367 11747
rect 14197 11713 14231 11747
rect 18153 11713 18187 11747
rect 21189 11713 21223 11747
rect 4925 11645 4959 11679
rect 5181 11645 5215 11679
rect 6929 11645 6963 11679
rect 7021 11645 7055 11679
rect 7297 11645 7331 11679
rect 8861 11645 8895 11679
rect 9137 11645 9171 11679
rect 9597 11645 9631 11679
rect 9689 11645 9723 11679
rect 10057 11645 10091 11679
rect 12173 11645 12207 11679
rect 13277 11645 13311 11679
rect 13369 11645 13403 11679
rect 13678 11645 13712 11679
rect 14473 11645 14507 11679
rect 15209 11645 15243 11679
rect 15669 11645 15703 11679
rect 15945 11645 15979 11679
rect 16037 11645 16071 11679
rect 18061 11645 18095 11679
rect 20922 11645 20956 11679
rect 9045 11577 9079 11611
rect 11989 11577 12023 11611
rect 13093 11577 13127 11611
rect 14289 11577 14323 11611
rect 15301 11577 15335 11611
rect 15853 11577 15887 11611
rect 6745 11509 6779 11543
rect 9229 11509 9263 11543
rect 10609 11509 10643 11543
rect 11805 11509 11839 11543
rect 13553 11509 13587 11543
rect 13737 11509 13771 11543
rect 14657 11509 14691 11543
rect 15393 11509 15427 11543
rect 15577 11509 15611 11543
rect 16221 11509 16255 11543
rect 8677 11305 8711 11339
rect 10333 11305 10367 11339
rect 10609 11305 10643 11339
rect 13093 11305 13127 11339
rect 13461 11305 13495 11339
rect 15209 11305 15243 11339
rect 10149 11237 10183 11271
rect 14657 11237 14691 11271
rect 16405 11237 16439 11271
rect 6745 11169 6779 11203
rect 6929 11169 6963 11203
rect 7113 11169 7147 11203
rect 7205 11169 7239 11203
rect 8125 11169 8159 11203
rect 8309 11169 8343 11203
rect 8674 11169 8708 11203
rect 10425 11169 10459 11203
rect 10517 11169 10551 11203
rect 10701 11169 10735 11203
rect 10977 11169 11011 11203
rect 11713 11169 11747 11203
rect 11969 11169 12003 11203
rect 13829 11169 13863 11203
rect 14565 11169 14599 11203
rect 14749 11169 14783 11203
rect 14841 11169 14875 11203
rect 15025 11169 15059 11203
rect 15577 11169 15611 11203
rect 15945 11169 15979 11203
rect 16129 11169 16163 11203
rect 16221 11169 16255 11203
rect 17702 11169 17736 11203
rect 17969 11169 18003 11203
rect 8217 11101 8251 11135
rect 9045 11101 9079 11135
rect 9137 11101 9171 11135
rect 11529 11101 11563 11135
rect 13737 11101 13771 11135
rect 8493 11033 8527 11067
rect 15393 11033 15427 11067
rect 16405 11033 16439 11067
rect 7389 10965 7423 10999
rect 10149 10965 10183 10999
rect 15853 10965 15887 10999
rect 16589 10965 16623 10999
rect 6285 10761 6319 10795
rect 11253 10761 11287 10795
rect 11621 10761 11655 10795
rect 17509 10761 17543 10795
rect 16681 10625 16715 10659
rect 7665 10557 7699 10591
rect 9873 10557 9907 10591
rect 11437 10557 11471 10591
rect 17325 10557 17359 10591
rect 17417 10557 17451 10591
rect 17601 10557 17635 10591
rect 7398 10489 7432 10523
rect 10140 10489 10174 10523
rect 9229 10217 9263 10251
rect 8116 10149 8150 10183
rect 7849 10081 7883 10115
<< metal1 >>
rect 552 28314 28428 28336
rect 552 28262 3882 28314
rect 3934 28262 3946 28314
rect 3998 28262 4010 28314
rect 4062 28262 4074 28314
rect 4126 28262 4138 28314
rect 4190 28262 10851 28314
rect 10903 28262 10915 28314
rect 10967 28262 10979 28314
rect 11031 28262 11043 28314
rect 11095 28262 11107 28314
rect 11159 28262 17820 28314
rect 17872 28262 17884 28314
rect 17936 28262 17948 28314
rect 18000 28262 18012 28314
rect 18064 28262 18076 28314
rect 18128 28262 24789 28314
rect 24841 28262 24853 28314
rect 24905 28262 24917 28314
rect 24969 28262 24981 28314
rect 25033 28262 25045 28314
rect 25097 28262 28428 28314
rect 552 28240 28428 28262
rect 11333 28203 11391 28209
rect 11333 28169 11345 28203
rect 11379 28200 11391 28203
rect 11422 28200 11428 28212
rect 11379 28172 11428 28200
rect 11379 28169 11391 28172
rect 11333 28163 11391 28169
rect 11422 28160 11428 28172
rect 11480 28160 11486 28212
rect 19518 28160 19524 28212
rect 19576 28160 19582 28212
rect 19536 28064 19564 28160
rect 19536 28036 20484 28064
rect 11146 27956 11152 28008
rect 11204 27956 11210 28008
rect 15654 27956 15660 28008
rect 15712 27956 15718 28008
rect 17494 27956 17500 28008
rect 17552 27996 17558 28008
rect 17589 27999 17647 28005
rect 17589 27996 17601 27999
rect 17552 27968 17601 27996
rect 17552 27956 17558 27968
rect 17589 27965 17601 27968
rect 17635 27965 17647 27999
rect 17589 27959 17647 27965
rect 19242 27956 19248 28008
rect 19300 27956 19306 28008
rect 20456 28005 20484 28036
rect 20165 27999 20223 28005
rect 20165 27965 20177 27999
rect 20211 27996 20223 27999
rect 20441 27999 20499 28005
rect 20211 27968 20300 27996
rect 20211 27965 20223 27968
rect 20165 27959 20223 27965
rect 15841 27863 15899 27869
rect 15841 27829 15853 27863
rect 15887 27860 15899 27863
rect 16206 27860 16212 27872
rect 15887 27832 16212 27860
rect 15887 27829 15899 27832
rect 15841 27823 15899 27829
rect 16206 27820 16212 27832
rect 16264 27820 16270 27872
rect 17773 27863 17831 27869
rect 17773 27829 17785 27863
rect 17819 27860 17831 27863
rect 18138 27860 18144 27872
rect 17819 27832 18144 27860
rect 17819 27829 17831 27832
rect 17773 27823 17831 27829
rect 18138 27820 18144 27832
rect 18196 27820 18202 27872
rect 19886 27820 19892 27872
rect 19944 27820 19950 27872
rect 20070 27820 20076 27872
rect 20128 27820 20134 27872
rect 20272 27869 20300 27968
rect 20441 27965 20453 27999
rect 20487 27965 20499 27999
rect 20441 27959 20499 27965
rect 21542 27956 21548 28008
rect 21600 27996 21606 28008
rect 21821 27999 21879 28005
rect 21821 27996 21833 27999
rect 21600 27968 21833 27996
rect 21600 27956 21606 27968
rect 21821 27965 21833 27968
rect 21867 27965 21879 27999
rect 21821 27959 21879 27965
rect 23566 27956 23572 28008
rect 23624 27996 23630 28008
rect 24029 27999 24087 28005
rect 24029 27996 24041 27999
rect 23624 27968 24041 27996
rect 23624 27956 23630 27968
rect 24029 27965 24041 27968
rect 24075 27965 24087 27999
rect 24029 27959 24087 27965
rect 25590 27956 25596 28008
rect 25648 27996 25654 28008
rect 25777 27999 25835 28005
rect 25777 27996 25789 27999
rect 25648 27968 25789 27996
rect 25648 27956 25654 27968
rect 25777 27965 25789 27968
rect 25823 27965 25835 27999
rect 25777 27959 25835 27965
rect 20257 27863 20315 27869
rect 20257 27829 20269 27863
rect 20303 27829 20315 27863
rect 20257 27823 20315 27829
rect 21634 27820 21640 27872
rect 21692 27820 21698 27872
rect 23842 27820 23848 27872
rect 23900 27820 23906 27872
rect 25866 27820 25872 27872
rect 25924 27820 25930 27872
rect 552 27770 28587 27792
rect 552 27718 7366 27770
rect 7418 27718 7430 27770
rect 7482 27718 7494 27770
rect 7546 27718 7558 27770
rect 7610 27718 7622 27770
rect 7674 27718 14335 27770
rect 14387 27718 14399 27770
rect 14451 27718 14463 27770
rect 14515 27718 14527 27770
rect 14579 27718 14591 27770
rect 14643 27718 21304 27770
rect 21356 27718 21368 27770
rect 21420 27718 21432 27770
rect 21484 27718 21496 27770
rect 21548 27718 21560 27770
rect 21612 27718 28273 27770
rect 28325 27718 28337 27770
rect 28389 27718 28401 27770
rect 28453 27718 28465 27770
rect 28517 27718 28529 27770
rect 28581 27718 28587 27770
rect 552 27696 28587 27718
rect 6733 27659 6791 27665
rect 6733 27625 6745 27659
rect 6779 27625 6791 27659
rect 6733 27619 6791 27625
rect 14553 27659 14611 27665
rect 14553 27625 14565 27659
rect 14599 27656 14611 27659
rect 15197 27659 15255 27665
rect 14599 27628 15148 27656
rect 14599 27625 14611 27628
rect 14553 27619 14611 27625
rect 1302 27548 1308 27600
rect 1360 27588 1366 27600
rect 1397 27591 1455 27597
rect 1397 27588 1409 27591
rect 1360 27560 1409 27588
rect 1360 27548 1366 27560
rect 1397 27557 1409 27560
rect 1443 27557 1455 27591
rect 1397 27551 1455 27557
rect 3326 27548 3332 27600
rect 3384 27588 3390 27600
rect 3789 27591 3847 27597
rect 3789 27588 3801 27591
rect 3384 27560 3801 27588
rect 3384 27548 3390 27560
rect 3789 27557 3801 27560
rect 3835 27557 3847 27591
rect 3789 27551 3847 27557
rect 4617 27591 4675 27597
rect 4617 27557 4629 27591
rect 4663 27588 4675 27591
rect 5169 27591 5227 27597
rect 4663 27560 4936 27588
rect 4663 27557 4675 27560
rect 4617 27551 4675 27557
rect 4908 27532 4936 27560
rect 5169 27557 5181 27591
rect 5215 27588 5227 27591
rect 5350 27588 5356 27600
rect 5215 27560 5356 27588
rect 5215 27557 5227 27560
rect 5169 27551 5227 27557
rect 5350 27548 5356 27560
rect 5408 27548 5414 27600
rect 6748 27588 6776 27619
rect 6748 27560 8248 27588
rect 1765 27523 1823 27529
rect 1765 27489 1777 27523
rect 1811 27520 1823 27523
rect 2222 27520 2228 27532
rect 1811 27492 2228 27520
rect 1811 27489 1823 27492
rect 1765 27483 1823 27489
rect 2222 27480 2228 27492
rect 2280 27480 2286 27532
rect 2590 27529 2596 27532
rect 2584 27483 2596 27529
rect 2590 27480 2596 27483
rect 2648 27480 2654 27532
rect 4157 27523 4215 27529
rect 4157 27489 4169 27523
rect 4203 27489 4215 27523
rect 4157 27483 4215 27489
rect 4801 27523 4859 27529
rect 4801 27489 4813 27523
rect 4847 27489 4859 27523
rect 4801 27483 4859 27489
rect 2314 27412 2320 27464
rect 2372 27412 2378 27464
rect 4172 27384 4200 27483
rect 4338 27412 4344 27464
rect 4396 27452 4402 27464
rect 4816 27452 4844 27483
rect 4890 27480 4896 27532
rect 4948 27480 4954 27532
rect 5077 27523 5135 27529
rect 5077 27489 5089 27523
rect 5123 27489 5135 27523
rect 5077 27483 5135 27489
rect 5092 27452 5120 27483
rect 5534 27480 5540 27532
rect 5592 27480 5598 27532
rect 5902 27480 5908 27532
rect 5960 27520 5966 27532
rect 5997 27523 6055 27529
rect 5997 27520 6009 27523
rect 5960 27492 6009 27520
rect 5960 27480 5966 27492
rect 5997 27489 6009 27492
rect 6043 27489 6055 27523
rect 5997 27483 6055 27489
rect 6365 27523 6423 27529
rect 6365 27489 6377 27523
rect 6411 27520 6423 27523
rect 7006 27520 7012 27532
rect 6411 27492 7012 27520
rect 6411 27489 6423 27492
rect 6365 27483 6423 27489
rect 7006 27480 7012 27492
rect 7064 27480 7070 27532
rect 7193 27523 7251 27529
rect 7193 27489 7205 27523
rect 7239 27520 7251 27523
rect 7561 27523 7619 27529
rect 7239 27492 7512 27520
rect 7239 27489 7251 27492
rect 7193 27483 7251 27489
rect 4396 27424 5120 27452
rect 4396 27412 4402 27424
rect 6086 27412 6092 27464
rect 6144 27452 6150 27464
rect 6273 27455 6331 27461
rect 6273 27452 6285 27455
rect 6144 27424 6285 27452
rect 6144 27412 6150 27424
rect 6273 27421 6285 27424
rect 6319 27421 6331 27455
rect 6273 27415 6331 27421
rect 6914 27384 6920 27396
rect 4172 27356 6920 27384
rect 6914 27344 6920 27356
rect 6972 27344 6978 27396
rect 7009 27387 7067 27393
rect 7009 27353 7021 27387
rect 7055 27384 7067 27387
rect 7282 27384 7288 27396
rect 7055 27356 7288 27384
rect 7055 27353 7067 27356
rect 7009 27347 7067 27353
rect 7282 27344 7288 27356
rect 7340 27344 7346 27396
rect 7484 27328 7512 27492
rect 7561 27489 7573 27523
rect 7607 27520 7619 27523
rect 7926 27520 7932 27532
rect 7607 27492 7932 27520
rect 7607 27489 7619 27492
rect 7561 27483 7619 27489
rect 7926 27480 7932 27492
rect 7984 27480 7990 27532
rect 8220 27529 8248 27560
rect 9508 27560 11192 27588
rect 9508 27532 9536 27560
rect 8205 27523 8263 27529
rect 8205 27489 8217 27523
rect 8251 27489 8263 27523
rect 8205 27483 8263 27489
rect 8938 27480 8944 27532
rect 8996 27480 9002 27532
rect 9401 27523 9459 27529
rect 9401 27489 9413 27523
rect 9447 27520 9459 27523
rect 9490 27520 9496 27532
rect 9447 27492 9496 27520
rect 9447 27489 9459 27492
rect 9401 27483 9459 27489
rect 9490 27480 9496 27492
rect 9548 27480 9554 27532
rect 9668 27523 9726 27529
rect 9668 27489 9680 27523
rect 9714 27520 9726 27523
rect 9950 27520 9956 27532
rect 9714 27492 9956 27520
rect 9714 27489 9726 27492
rect 9668 27483 9726 27489
rect 9950 27480 9956 27492
rect 10008 27480 10014 27532
rect 11164 27529 11192 27560
rect 13188 27560 14964 27588
rect 11149 27523 11207 27529
rect 11149 27489 11161 27523
rect 11195 27489 11207 27523
rect 11149 27483 11207 27489
rect 11238 27480 11244 27532
rect 11296 27520 11302 27532
rect 13188 27529 13216 27560
rect 11405 27523 11463 27529
rect 11405 27520 11417 27523
rect 11296 27492 11417 27520
rect 11296 27480 11302 27492
rect 11405 27489 11417 27492
rect 11451 27489 11463 27523
rect 12713 27523 12771 27529
rect 12713 27520 12725 27523
rect 11405 27483 11463 27489
rect 12544 27492 12725 27520
rect 7653 27455 7711 27461
rect 7653 27421 7665 27455
rect 7699 27452 7711 27455
rect 7834 27452 7840 27464
rect 7699 27424 7840 27452
rect 7699 27421 7711 27424
rect 7653 27415 7711 27421
rect 7834 27412 7840 27424
rect 7892 27412 7898 27464
rect 8113 27455 8171 27461
rect 8113 27421 8125 27455
rect 8159 27421 8171 27455
rect 8113 27415 8171 27421
rect 8573 27455 8631 27461
rect 8573 27421 8585 27455
rect 8619 27452 8631 27455
rect 8849 27455 8907 27461
rect 8849 27452 8861 27455
rect 8619 27424 8861 27452
rect 8619 27421 8631 27424
rect 8573 27415 8631 27421
rect 8849 27421 8861 27424
rect 8895 27421 8907 27455
rect 8849 27415 8907 27421
rect 7929 27387 7987 27393
rect 7929 27353 7941 27387
rect 7975 27384 7987 27387
rect 8128 27384 8156 27415
rect 7975 27356 8156 27384
rect 7975 27353 7987 27356
rect 7929 27347 7987 27353
rect 11146 27344 11152 27396
rect 11204 27344 11210 27396
rect 12544 27393 12572 27492
rect 12713 27489 12725 27492
rect 12759 27489 12771 27523
rect 12713 27483 12771 27489
rect 13173 27523 13231 27529
rect 13173 27489 13185 27523
rect 13219 27489 13231 27523
rect 13173 27483 13231 27489
rect 13262 27480 13268 27532
rect 13320 27520 13326 27532
rect 13429 27523 13487 27529
rect 13429 27520 13441 27523
rect 13320 27492 13441 27520
rect 13320 27480 13326 27492
rect 13429 27489 13441 27492
rect 13475 27489 13487 27523
rect 14936 27520 14964 27560
rect 15010 27548 15016 27600
rect 15068 27548 15074 27600
rect 15120 27588 15148 27628
rect 15197 27625 15209 27659
rect 15243 27656 15255 27659
rect 15654 27656 15660 27668
rect 15243 27628 15660 27656
rect 15243 27625 15255 27628
rect 15197 27619 15255 27625
rect 15654 27616 15660 27628
rect 15712 27616 15718 27668
rect 19061 27659 19119 27665
rect 19061 27625 19073 27659
rect 19107 27656 19119 27659
rect 19242 27656 19248 27668
rect 19107 27628 19248 27656
rect 19107 27625 19119 27628
rect 19061 27619 19119 27625
rect 19242 27616 19248 27628
rect 19300 27616 19306 27668
rect 21634 27616 21640 27668
rect 21692 27616 21698 27668
rect 15381 27591 15439 27597
rect 15381 27588 15393 27591
rect 15120 27560 15393 27588
rect 15381 27557 15393 27560
rect 15427 27557 15439 27591
rect 15381 27551 15439 27557
rect 15470 27548 15476 27600
rect 15528 27588 15534 27600
rect 15749 27591 15807 27597
rect 15749 27588 15761 27591
rect 15528 27560 15761 27588
rect 15528 27548 15534 27560
rect 15749 27557 15761 27560
rect 15795 27557 15807 27591
rect 19420 27591 19478 27597
rect 15749 27551 15807 27557
rect 16132 27560 17724 27588
rect 15194 27520 15200 27532
rect 14936 27492 15200 27520
rect 13429 27483 13487 27489
rect 15194 27480 15200 27492
rect 15252 27480 15258 27532
rect 15212 27452 15240 27480
rect 16132 27464 16160 27560
rect 16206 27480 16212 27532
rect 16264 27520 16270 27532
rect 17696 27529 17724 27560
rect 19420 27557 19432 27591
rect 19466 27588 19478 27591
rect 19886 27588 19892 27600
rect 19466 27560 19892 27588
rect 19466 27557 19478 27560
rect 19420 27551 19478 27557
rect 19886 27548 19892 27560
rect 19944 27548 19950 27600
rect 16373 27523 16431 27529
rect 16373 27520 16385 27523
rect 16264 27492 16385 27520
rect 16264 27480 16270 27492
rect 16373 27489 16385 27492
rect 16419 27489 16431 27523
rect 16373 27483 16431 27489
rect 17681 27523 17739 27529
rect 17681 27489 17693 27523
rect 17727 27489 17739 27523
rect 17681 27483 17739 27489
rect 17948 27523 18006 27529
rect 17948 27489 17960 27523
rect 17994 27520 18006 27523
rect 18322 27520 18328 27532
rect 17994 27492 18328 27520
rect 17994 27489 18006 27492
rect 17948 27483 18006 27489
rect 18322 27480 18328 27492
rect 18380 27480 18386 27532
rect 20625 27523 20683 27529
rect 20625 27520 20637 27523
rect 20548 27492 20637 27520
rect 16114 27452 16120 27464
rect 15212 27424 16120 27452
rect 16114 27412 16120 27424
rect 16172 27412 16178 27464
rect 19153 27455 19211 27461
rect 19153 27421 19165 27455
rect 19199 27421 19211 27455
rect 19153 27415 19211 27421
rect 12529 27387 12587 27393
rect 12529 27353 12541 27387
rect 12575 27353 12587 27387
rect 12529 27347 12587 27353
rect 14182 27344 14188 27396
rect 14240 27384 14246 27396
rect 14645 27387 14703 27393
rect 14645 27384 14657 27387
rect 14240 27356 14657 27384
rect 14240 27344 14246 27356
rect 14645 27353 14657 27356
rect 14691 27353 14703 27387
rect 14645 27347 14703 27353
rect 3694 27276 3700 27328
rect 3752 27276 3758 27328
rect 4430 27276 4436 27328
rect 4488 27276 4494 27328
rect 4982 27276 4988 27328
rect 5040 27276 5046 27328
rect 5813 27319 5871 27325
rect 5813 27285 5825 27319
rect 5859 27316 5871 27319
rect 5994 27316 6000 27328
rect 5859 27288 6000 27316
rect 5859 27285 5871 27288
rect 5813 27279 5871 27285
rect 5994 27276 6000 27288
rect 6052 27276 6058 27328
rect 7466 27276 7472 27328
rect 7524 27276 7530 27328
rect 9217 27319 9275 27325
rect 9217 27285 9229 27319
rect 9263 27316 9275 27319
rect 10686 27316 10692 27328
rect 9263 27288 10692 27316
rect 9263 27285 9275 27288
rect 9217 27279 9275 27285
rect 10686 27276 10692 27288
rect 10744 27276 10750 27328
rect 10781 27319 10839 27325
rect 10781 27285 10793 27319
rect 10827 27316 10839 27319
rect 11164 27316 11192 27344
rect 10827 27288 11192 27316
rect 12989 27319 13047 27325
rect 10827 27285 10839 27288
rect 10781 27279 10839 27285
rect 12989 27285 13001 27319
rect 13035 27316 13047 27319
rect 13446 27316 13452 27328
rect 13035 27288 13452 27316
rect 13035 27285 13047 27288
rect 12989 27279 13047 27285
rect 13446 27276 13452 27288
rect 13504 27276 13510 27328
rect 14826 27276 14832 27328
rect 14884 27316 14890 27328
rect 15013 27319 15071 27325
rect 15013 27316 15025 27319
rect 14884 27288 15025 27316
rect 14884 27276 14890 27288
rect 15013 27285 15025 27288
rect 15059 27285 15071 27319
rect 15013 27279 15071 27285
rect 15102 27276 15108 27328
rect 15160 27316 15166 27328
rect 17497 27319 17555 27325
rect 17497 27316 17509 27319
rect 15160 27288 17509 27316
rect 15160 27276 15166 27288
rect 17497 27285 17509 27288
rect 17543 27285 17555 27319
rect 19168 27316 19196 27415
rect 20548 27393 20576 27492
rect 20625 27489 20637 27492
rect 20671 27489 20683 27523
rect 20625 27483 20683 27489
rect 21085 27523 21143 27529
rect 21085 27489 21097 27523
rect 21131 27520 21143 27523
rect 21652 27520 21680 27616
rect 21131 27492 21680 27520
rect 22669 27523 22727 27529
rect 21131 27489 21143 27492
rect 21085 27483 21143 27489
rect 22669 27489 22681 27523
rect 22715 27520 22727 27523
rect 22830 27520 22836 27532
rect 22715 27492 22836 27520
rect 22715 27489 22727 27492
rect 22669 27483 22727 27489
rect 22830 27480 22836 27492
rect 22888 27480 22894 27532
rect 23290 27529 23296 27532
rect 23284 27483 23296 27529
rect 23290 27480 23296 27483
rect 23348 27480 23354 27532
rect 22925 27455 22983 27461
rect 22925 27421 22937 27455
rect 22971 27452 22983 27455
rect 23017 27455 23075 27461
rect 23017 27452 23029 27455
rect 22971 27424 23029 27452
rect 22971 27421 22983 27424
rect 22925 27415 22983 27421
rect 23017 27421 23029 27424
rect 23063 27421 23075 27455
rect 23017 27415 23075 27421
rect 20533 27387 20591 27393
rect 20533 27353 20545 27387
rect 20579 27353 20591 27387
rect 20533 27347 20591 27353
rect 20622 27344 20628 27396
rect 20680 27384 20686 27396
rect 21545 27387 21603 27393
rect 21545 27384 21557 27387
rect 20680 27356 21557 27384
rect 20680 27344 20686 27356
rect 21545 27353 21557 27356
rect 21591 27353 21603 27387
rect 21545 27347 21603 27353
rect 22940 27328 22968 27415
rect 19426 27316 19432 27328
rect 19168 27288 19432 27316
rect 17497 27279 17555 27285
rect 19426 27276 19432 27288
rect 19484 27276 19490 27328
rect 20714 27276 20720 27328
rect 20772 27276 20778 27328
rect 20898 27276 20904 27328
rect 20956 27316 20962 27328
rect 20993 27319 21051 27325
rect 20993 27316 21005 27319
rect 20956 27288 21005 27316
rect 20956 27276 20962 27288
rect 20993 27285 21005 27288
rect 21039 27285 21051 27319
rect 20993 27279 21051 27285
rect 22922 27276 22928 27328
rect 22980 27276 22986 27328
rect 24394 27276 24400 27328
rect 24452 27276 24458 27328
rect 552 27226 28428 27248
rect 552 27174 3882 27226
rect 3934 27174 3946 27226
rect 3998 27174 4010 27226
rect 4062 27174 4074 27226
rect 4126 27174 4138 27226
rect 4190 27174 10851 27226
rect 10903 27174 10915 27226
rect 10967 27174 10979 27226
rect 11031 27174 11043 27226
rect 11095 27174 11107 27226
rect 11159 27174 17820 27226
rect 17872 27174 17884 27226
rect 17936 27174 17948 27226
rect 18000 27174 18012 27226
rect 18064 27174 18076 27226
rect 18128 27174 24789 27226
rect 24841 27174 24853 27226
rect 24905 27174 24917 27226
rect 24969 27174 24981 27226
rect 25033 27174 25045 27226
rect 25097 27174 28428 27226
rect 552 27152 28428 27174
rect 2590 27072 2596 27124
rect 2648 27112 2654 27124
rect 2777 27115 2835 27121
rect 2777 27112 2789 27115
rect 2648 27084 2789 27112
rect 2648 27072 2654 27084
rect 2777 27081 2789 27084
rect 2823 27081 2835 27115
rect 2777 27075 2835 27081
rect 3421 27115 3479 27121
rect 3421 27081 3433 27115
rect 3467 27112 3479 27115
rect 4522 27112 4528 27124
rect 3467 27084 4528 27112
rect 3467 27081 3479 27084
rect 3421 27075 3479 27081
rect 4522 27072 4528 27084
rect 4580 27072 4586 27124
rect 7834 27072 7840 27124
rect 7892 27072 7898 27124
rect 8941 27115 8999 27121
rect 8941 27081 8953 27115
rect 8987 27112 8999 27115
rect 9398 27112 9404 27124
rect 8987 27084 9404 27112
rect 8987 27081 8999 27084
rect 8941 27075 8999 27081
rect 9398 27072 9404 27084
rect 9456 27072 9462 27124
rect 10686 27072 10692 27124
rect 10744 27072 10750 27124
rect 11333 27115 11391 27121
rect 11333 27112 11345 27115
rect 11164 27084 11345 27112
rect 3237 27047 3295 27053
rect 3237 27013 3249 27047
rect 3283 27013 3295 27047
rect 3237 27007 3295 27013
rect 2961 26911 3019 26917
rect 2961 26877 2973 26911
rect 3007 26908 3019 26911
rect 3252 26908 3280 27007
rect 3694 27004 3700 27056
rect 3752 27004 3758 27056
rect 4890 27044 4896 27056
rect 4264 27016 4896 27044
rect 3712 26976 3740 27004
rect 3712 26948 4108 26976
rect 3007 26880 3280 26908
rect 3007 26877 3019 26880
rect 2961 26871 3019 26877
rect 3694 26868 3700 26920
rect 3752 26908 3758 26920
rect 4080 26917 4108 26948
rect 3789 26911 3847 26917
rect 3789 26908 3801 26911
rect 3752 26880 3801 26908
rect 3752 26868 3758 26880
rect 3789 26877 3801 26880
rect 3835 26877 3847 26911
rect 3789 26871 3847 26877
rect 4065 26911 4123 26917
rect 4065 26877 4077 26911
rect 4111 26877 4123 26911
rect 4065 26871 4123 26877
rect 4264 26784 4292 27016
rect 4890 27004 4896 27016
rect 4948 27004 4954 27056
rect 7742 27004 7748 27056
rect 7800 27004 7806 27056
rect 4341 26911 4399 26917
rect 4341 26877 4353 26911
rect 4387 26877 4399 26911
rect 4341 26871 4399 26877
rect 4356 26784 4384 26871
rect 5994 26868 6000 26920
rect 6052 26917 6058 26920
rect 6052 26908 6064 26917
rect 6052 26880 6097 26908
rect 6052 26871 6064 26880
rect 6052 26868 6058 26871
rect 6270 26868 6276 26920
rect 6328 26868 6334 26920
rect 8754 26868 8760 26920
rect 8812 26868 8818 26920
rect 10704 26908 10732 27072
rect 11164 27044 11192 27084
rect 11333 27081 11345 27084
rect 11379 27081 11391 27115
rect 11333 27075 11391 27081
rect 13081 27115 13139 27121
rect 13081 27081 13093 27115
rect 13127 27112 13139 27115
rect 13262 27112 13268 27124
rect 13127 27084 13268 27112
rect 13127 27081 13139 27084
rect 13081 27075 13139 27081
rect 13262 27072 13268 27084
rect 13320 27072 13326 27124
rect 15010 27072 15016 27124
rect 15068 27072 15074 27124
rect 18322 27072 18328 27124
rect 18380 27072 18386 27124
rect 19076 27084 21680 27112
rect 11793 27047 11851 27053
rect 11793 27044 11805 27047
rect 11164 27016 11805 27044
rect 11164 26988 11192 27016
rect 11793 27013 11805 27016
rect 11839 27013 11851 27047
rect 11793 27007 11851 27013
rect 16758 27004 16764 27056
rect 16816 27044 16822 27056
rect 19076 27044 19104 27084
rect 16816 27016 17540 27044
rect 16816 27004 16822 27016
rect 11146 26936 11152 26988
rect 11204 26936 11210 26988
rect 11701 26979 11759 26985
rect 11701 26945 11713 26979
rect 11747 26945 11759 26979
rect 11701 26939 11759 26945
rect 12345 26979 12403 26985
rect 12345 26945 12357 26979
rect 12391 26976 12403 26979
rect 12391 26948 12756 26976
rect 12391 26945 12403 26948
rect 12345 26939 12403 26945
rect 11241 26911 11299 26917
rect 11241 26908 11253 26911
rect 10704 26880 11253 26908
rect 11241 26877 11253 26880
rect 11287 26908 11299 26911
rect 11716 26908 11744 26939
rect 11287 26880 11560 26908
rect 11716 26880 12388 26908
rect 11287 26877 11299 26880
rect 11241 26871 11299 26877
rect 7282 26800 7288 26852
rect 7340 26840 7346 26852
rect 7377 26843 7435 26849
rect 7377 26840 7389 26843
rect 7340 26812 7389 26840
rect 7340 26800 7346 26812
rect 7377 26809 7389 26812
rect 7423 26809 7435 26843
rect 11532 26840 11560 26880
rect 12161 26843 12219 26849
rect 12161 26840 12173 26843
rect 11532 26812 12173 26840
rect 7377 26803 7435 26809
rect 12161 26809 12173 26812
rect 12207 26809 12219 26843
rect 12360 26840 12388 26880
rect 12434 26868 12440 26920
rect 12492 26868 12498 26920
rect 12728 26917 12756 26948
rect 15194 26936 15200 26988
rect 15252 26976 15258 26988
rect 17512 26985 17540 27016
rect 17880 27016 19104 27044
rect 15381 26979 15439 26985
rect 15381 26976 15393 26979
rect 15252 26948 15393 26976
rect 15252 26936 15258 26948
rect 15381 26945 15393 26948
rect 15427 26945 15439 26979
rect 15381 26939 15439 26945
rect 17497 26979 17555 26985
rect 17497 26945 17509 26979
rect 17543 26945 17555 26979
rect 17497 26939 17555 26945
rect 12621 26911 12679 26917
rect 12621 26877 12633 26911
rect 12667 26877 12679 26911
rect 12621 26871 12679 26877
rect 12713 26911 12771 26917
rect 12713 26877 12725 26911
rect 12759 26877 12771 26911
rect 12713 26871 12771 26877
rect 12636 26840 12664 26871
rect 12802 26868 12808 26920
rect 12860 26868 12866 26920
rect 14645 26911 14703 26917
rect 14645 26877 14657 26911
rect 14691 26908 14703 26911
rect 14734 26908 14740 26920
rect 14691 26880 14740 26908
rect 14691 26877 14703 26880
rect 14645 26871 14703 26877
rect 14734 26868 14740 26880
rect 14792 26908 14798 26920
rect 15105 26911 15163 26917
rect 15105 26908 15117 26911
rect 14792 26880 15117 26908
rect 14792 26868 14798 26880
rect 15105 26877 15117 26880
rect 15151 26877 15163 26911
rect 15105 26871 15163 26877
rect 15286 26868 15292 26920
rect 15344 26868 15350 26920
rect 16666 26868 16672 26920
rect 16724 26908 16730 26920
rect 17880 26917 17908 27016
rect 17865 26911 17923 26917
rect 17865 26908 17877 26911
rect 16724 26880 17877 26908
rect 16724 26868 16730 26880
rect 17865 26877 17877 26880
rect 17911 26877 17923 26911
rect 17865 26871 17923 26877
rect 18138 26868 18144 26920
rect 18196 26908 18202 26920
rect 18233 26911 18291 26917
rect 18233 26908 18245 26911
rect 18196 26880 18245 26908
rect 18196 26868 18202 26880
rect 18233 26877 18245 26880
rect 18279 26877 18291 26911
rect 18233 26871 18291 26877
rect 19061 26911 19119 26917
rect 19061 26877 19073 26911
rect 19107 26908 19119 26911
rect 20438 26908 20444 26920
rect 19107 26880 20444 26908
rect 19107 26877 19119 26880
rect 19061 26871 19119 26877
rect 19444 26852 19472 26880
rect 20438 26868 20444 26880
rect 20496 26908 20502 26920
rect 20898 26917 20904 26920
rect 20625 26911 20683 26917
rect 20625 26908 20637 26911
rect 20496 26880 20637 26908
rect 20496 26868 20502 26880
rect 20625 26877 20637 26880
rect 20671 26877 20683 26911
rect 20892 26908 20904 26917
rect 20859 26880 20904 26908
rect 20625 26871 20683 26877
rect 20892 26871 20904 26880
rect 20898 26868 20904 26871
rect 20956 26868 20962 26920
rect 12360 26812 12664 26840
rect 14829 26843 14887 26849
rect 12161 26803 12219 26809
rect 14829 26809 14841 26843
rect 14875 26809 14887 26843
rect 14829 26803 14887 26809
rect 15197 26843 15255 26849
rect 15197 26809 15209 26843
rect 15243 26840 15255 26843
rect 15626 26843 15684 26849
rect 15626 26840 15638 26843
rect 15243 26812 15638 26840
rect 15243 26809 15255 26812
rect 15197 26803 15255 26809
rect 15626 26809 15638 26812
rect 15672 26809 15684 26843
rect 15626 26803 15684 26809
rect 19328 26843 19386 26849
rect 19328 26809 19340 26843
rect 19374 26809 19386 26843
rect 19328 26803 19386 26809
rect 3421 26775 3479 26781
rect 3421 26741 3433 26775
rect 3467 26772 3479 26775
rect 3881 26775 3939 26781
rect 3881 26772 3893 26775
rect 3467 26744 3893 26772
rect 3467 26741 3479 26744
rect 3421 26735 3479 26741
rect 3881 26741 3893 26744
rect 3927 26741 3939 26775
rect 3881 26735 3939 26741
rect 4246 26732 4252 26784
rect 4304 26732 4310 26784
rect 4338 26732 4344 26784
rect 4396 26732 4402 26784
rect 7466 26732 7472 26784
rect 7524 26772 7530 26784
rect 11422 26772 11428 26784
rect 7524 26744 11428 26772
rect 7524 26732 7530 26744
rect 11422 26732 11428 26744
rect 11480 26732 11486 26784
rect 11974 26732 11980 26784
rect 12032 26732 12038 26784
rect 12069 26775 12127 26781
rect 12069 26741 12081 26775
rect 12115 26772 12127 26775
rect 12618 26772 12624 26784
rect 12115 26744 12624 26772
rect 12115 26741 12127 26744
rect 12069 26735 12127 26741
rect 12618 26732 12624 26744
rect 12676 26732 12682 26784
rect 13906 26732 13912 26784
rect 13964 26772 13970 26784
rect 14844 26772 14872 26803
rect 15102 26772 15108 26784
rect 13964 26744 15108 26772
rect 13964 26732 13970 26744
rect 15102 26732 15108 26744
rect 15160 26732 15166 26784
rect 16942 26732 16948 26784
rect 17000 26732 17006 26784
rect 18049 26775 18107 26781
rect 18049 26741 18061 26775
rect 18095 26772 18107 26775
rect 18138 26772 18144 26784
rect 18095 26744 18144 26772
rect 18095 26741 18107 26744
rect 18049 26735 18107 26741
rect 18138 26732 18144 26744
rect 18196 26732 18202 26784
rect 19352 26772 19380 26803
rect 19426 26800 19432 26852
rect 19484 26800 19490 26852
rect 20070 26800 20076 26852
rect 20128 26800 20134 26852
rect 21652 26840 21680 27084
rect 22830 27072 22836 27124
rect 22888 27112 22894 27124
rect 23017 27115 23075 27121
rect 23017 27112 23029 27115
rect 22888 27084 23029 27112
rect 22888 27072 22894 27084
rect 23017 27081 23029 27084
rect 23063 27081 23075 27115
rect 23017 27075 23075 27081
rect 23201 27115 23259 27121
rect 23201 27081 23213 27115
rect 23247 27112 23259 27115
rect 23290 27112 23296 27124
rect 23247 27084 23296 27112
rect 23247 27081 23259 27084
rect 23201 27075 23259 27081
rect 23290 27072 23296 27084
rect 23348 27072 23354 27124
rect 24394 27072 24400 27124
rect 24452 27072 24458 27124
rect 22005 27047 22063 27053
rect 22005 27013 22017 27047
rect 22051 27044 22063 27047
rect 22051 27016 22416 27044
rect 22051 27013 22063 27016
rect 22005 27007 22063 27013
rect 22388 26985 22416 27016
rect 22373 26979 22431 26985
rect 22373 26945 22385 26979
rect 22419 26945 22431 26979
rect 24412 26976 24440 27072
rect 24857 26979 24915 26985
rect 24857 26976 24869 26979
rect 24412 26948 24869 26976
rect 22373 26939 22431 26945
rect 24857 26945 24869 26948
rect 24903 26945 24915 26979
rect 24857 26939 24915 26945
rect 23293 26911 23351 26917
rect 23293 26877 23305 26911
rect 23339 26908 23351 26911
rect 23842 26908 23848 26920
rect 23339 26880 23848 26908
rect 23339 26877 23351 26880
rect 23293 26871 23351 26877
rect 23842 26868 23848 26880
rect 23900 26868 23906 26920
rect 23750 26840 23756 26852
rect 21652 26812 23756 26840
rect 23750 26800 23756 26812
rect 23808 26840 23814 26852
rect 25866 26840 25872 26852
rect 23808 26812 25872 26840
rect 23808 26800 23814 26812
rect 25866 26800 25872 26812
rect 25924 26800 25930 26852
rect 20088 26772 20116 26800
rect 19352 26744 20116 26772
rect 20346 26732 20352 26784
rect 20404 26772 20410 26784
rect 20441 26775 20499 26781
rect 20441 26772 20453 26775
rect 20404 26744 20453 26772
rect 20404 26732 20410 26744
rect 20441 26741 20453 26744
rect 20487 26741 20499 26775
rect 20441 26735 20499 26741
rect 24210 26732 24216 26784
rect 24268 26772 24274 26784
rect 24305 26775 24363 26781
rect 24305 26772 24317 26775
rect 24268 26744 24317 26772
rect 24268 26732 24274 26744
rect 24305 26741 24317 26744
rect 24351 26741 24363 26775
rect 24305 26735 24363 26741
rect 552 26682 28587 26704
rect 552 26630 7366 26682
rect 7418 26630 7430 26682
rect 7482 26630 7494 26682
rect 7546 26630 7558 26682
rect 7610 26630 7622 26682
rect 7674 26630 14335 26682
rect 14387 26630 14399 26682
rect 14451 26630 14463 26682
rect 14515 26630 14527 26682
rect 14579 26630 14591 26682
rect 14643 26630 21304 26682
rect 21356 26630 21368 26682
rect 21420 26630 21432 26682
rect 21484 26630 21496 26682
rect 21548 26630 21560 26682
rect 21612 26630 28273 26682
rect 28325 26630 28337 26682
rect 28389 26630 28401 26682
rect 28453 26630 28465 26682
rect 28517 26630 28529 26682
rect 28581 26630 28587 26682
rect 552 26608 28587 26630
rect 4551 26571 4609 26577
rect 4551 26537 4563 26571
rect 4597 26568 4609 26571
rect 4982 26568 4988 26580
rect 4597 26540 4988 26568
rect 4597 26537 4609 26540
rect 4551 26531 4609 26537
rect 4982 26528 4988 26540
rect 5040 26528 5046 26580
rect 6086 26528 6092 26580
rect 6144 26528 6150 26580
rect 7282 26528 7288 26580
rect 7340 26568 7346 26580
rect 7377 26571 7435 26577
rect 7377 26568 7389 26571
rect 7340 26540 7389 26568
rect 7340 26528 7346 26540
rect 7377 26537 7389 26540
rect 7423 26568 7435 26571
rect 7558 26568 7564 26580
rect 7423 26540 7564 26568
rect 7423 26537 7435 26540
rect 7377 26531 7435 26537
rect 7558 26528 7564 26540
rect 7616 26528 7622 26580
rect 7742 26528 7748 26580
rect 7800 26568 7806 26580
rect 8021 26571 8079 26577
rect 8021 26568 8033 26571
rect 7800 26540 8033 26568
rect 7800 26528 7806 26540
rect 8021 26537 8033 26540
rect 8067 26537 8079 26571
rect 10413 26571 10471 26577
rect 8021 26531 8079 26537
rect 9646 26540 10180 26568
rect 4341 26503 4399 26509
rect 4341 26469 4353 26503
rect 4387 26500 4399 26503
rect 9646 26500 9674 26540
rect 4387 26472 4568 26500
rect 4387 26469 4399 26472
rect 4341 26463 4399 26469
rect 4540 26376 4568 26472
rect 7300 26472 8064 26500
rect 6822 26392 6828 26444
rect 6880 26432 6886 26444
rect 7300 26441 7328 26472
rect 7392 26441 7512 26442
rect 7285 26435 7343 26441
rect 7285 26432 7297 26435
rect 6880 26404 7297 26432
rect 6880 26392 6886 26404
rect 7285 26401 7297 26404
rect 7331 26401 7343 26435
rect 7285 26395 7343 26401
rect 7392 26435 7527 26441
rect 7392 26414 7481 26435
rect 4522 26324 4528 26376
rect 4580 26324 4586 26376
rect 5902 26324 5908 26376
rect 5960 26324 5966 26376
rect 6546 26324 6552 26376
rect 6604 26324 6610 26376
rect 7392 26364 7420 26414
rect 7469 26401 7481 26414
rect 7515 26401 7527 26435
rect 7469 26395 7527 26401
rect 7558 26392 7564 26444
rect 7616 26392 7622 26444
rect 7834 26392 7840 26444
rect 7892 26392 7898 26444
rect 7929 26435 7987 26441
rect 7929 26401 7941 26435
rect 7975 26432 7987 26435
rect 8036 26432 8064 26472
rect 8128 26472 9674 26500
rect 8128 26441 8156 26472
rect 7975 26404 8064 26432
rect 8113 26435 8171 26441
rect 7975 26401 7987 26404
rect 7929 26395 7987 26401
rect 8113 26401 8125 26435
rect 8159 26401 8171 26435
rect 8113 26395 8171 26401
rect 9309 26435 9367 26441
rect 9309 26401 9321 26435
rect 9355 26401 9367 26435
rect 9309 26395 9367 26401
rect 8128 26364 8156 26395
rect 7392 26336 8156 26364
rect 9217 26367 9275 26373
rect 9217 26333 9229 26367
rect 9263 26333 9275 26367
rect 9324 26364 9352 26395
rect 10042 26392 10048 26444
rect 10100 26392 10106 26444
rect 9953 26367 10011 26373
rect 9324 26336 9628 26364
rect 9217 26327 9275 26333
rect 4709 26299 4767 26305
rect 4709 26265 4721 26299
rect 4755 26296 4767 26299
rect 5920 26296 5948 26324
rect 4755 26268 5948 26296
rect 6273 26299 6331 26305
rect 4755 26265 4767 26268
rect 4709 26259 4767 26265
rect 6273 26265 6285 26299
rect 6319 26296 6331 26299
rect 6362 26296 6368 26308
rect 6319 26268 6368 26296
rect 6319 26265 6331 26268
rect 6273 26259 6331 26265
rect 6362 26256 6368 26268
rect 6420 26256 6426 26308
rect 7561 26299 7619 26305
rect 7561 26265 7573 26299
rect 7607 26265 7619 26299
rect 7561 26259 7619 26265
rect 4430 26188 4436 26240
rect 4488 26228 4494 26240
rect 4525 26231 4583 26237
rect 4525 26228 4537 26231
rect 4488 26200 4537 26228
rect 4488 26188 4494 26200
rect 4525 26197 4537 26200
rect 4571 26197 4583 26231
rect 7576 26228 7604 26259
rect 9232 26228 9260 26327
rect 7576 26200 9260 26228
rect 9600 26228 9628 26336
rect 9953 26333 9965 26367
rect 9999 26333 10011 26367
rect 10152 26364 10180 26540
rect 10413 26537 10425 26571
rect 10459 26568 10471 26571
rect 11146 26568 11152 26580
rect 10459 26540 11152 26568
rect 10459 26537 10471 26540
rect 10413 26531 10471 26537
rect 11146 26528 11152 26540
rect 11204 26528 11210 26580
rect 11974 26528 11980 26580
rect 12032 26568 12038 26580
rect 12032 26540 12572 26568
rect 12032 26528 12038 26540
rect 11164 26432 11192 26528
rect 12544 26444 12572 26540
rect 12802 26528 12808 26580
rect 12860 26528 12866 26580
rect 14182 26528 14188 26580
rect 14240 26528 14246 26580
rect 14734 26528 14740 26580
rect 14792 26528 14798 26580
rect 14829 26571 14887 26577
rect 14829 26537 14841 26571
rect 14875 26568 14887 26571
rect 15286 26568 15292 26580
rect 14875 26540 15292 26568
rect 14875 26537 14887 26540
rect 14829 26531 14887 26537
rect 15286 26528 15292 26540
rect 15344 26528 15350 26580
rect 16942 26528 16948 26580
rect 17000 26528 17006 26580
rect 12161 26435 12219 26441
rect 12161 26432 12173 26435
rect 11164 26404 12173 26432
rect 12161 26401 12173 26404
rect 12207 26401 12219 26435
rect 12161 26395 12219 26401
rect 12250 26392 12256 26444
rect 12308 26392 12314 26444
rect 12342 26392 12348 26444
rect 12400 26432 12406 26444
rect 12437 26435 12495 26441
rect 12437 26432 12449 26435
rect 12400 26404 12449 26432
rect 12400 26392 12406 26404
rect 12437 26401 12449 26404
rect 12483 26401 12495 26435
rect 12437 26395 12495 26401
rect 12526 26392 12532 26444
rect 12584 26392 12590 26444
rect 12618 26392 12624 26444
rect 12676 26392 12682 26444
rect 10152 26336 11836 26364
rect 9953 26327 10011 26333
rect 9677 26299 9735 26305
rect 9677 26265 9689 26299
rect 9723 26296 9735 26299
rect 9968 26296 9996 26327
rect 11808 26308 11836 26336
rect 11606 26296 11612 26308
rect 9723 26268 9996 26296
rect 10060 26268 11612 26296
rect 9723 26265 9735 26268
rect 9677 26259 9735 26265
rect 10060 26228 10088 26268
rect 11606 26256 11612 26268
rect 11664 26256 11670 26308
rect 11790 26256 11796 26308
rect 11848 26256 11854 26308
rect 12636 26296 12664 26392
rect 12713 26367 12771 26373
rect 12713 26333 12725 26367
rect 12759 26364 12771 26367
rect 12820 26364 12848 26528
rect 13817 26503 13875 26509
rect 13817 26469 13829 26503
rect 13863 26500 13875 26503
rect 13906 26500 13912 26512
rect 13863 26472 13912 26500
rect 13863 26469 13875 26472
rect 13817 26463 13875 26469
rect 13906 26460 13912 26472
rect 13964 26460 13970 26512
rect 16960 26500 16988 26528
rect 14047 26469 14105 26475
rect 14047 26435 14059 26469
rect 14093 26435 14105 26469
rect 15120 26472 16988 26500
rect 15120 26441 15148 26472
rect 14047 26432 14105 26435
rect 14553 26435 14611 26441
rect 14553 26432 14565 26435
rect 14047 26429 14565 26432
rect 14048 26404 14565 26429
rect 14553 26401 14565 26404
rect 14599 26432 14611 26435
rect 15105 26435 15163 26441
rect 14599 26404 15056 26432
rect 14599 26401 14611 26404
rect 14553 26395 14611 26401
rect 12759 26336 12848 26364
rect 14369 26367 14427 26373
rect 12759 26333 12771 26336
rect 12713 26327 12771 26333
rect 14369 26333 14381 26367
rect 14415 26333 14427 26367
rect 14369 26327 14427 26333
rect 13078 26296 13084 26308
rect 12636 26268 13084 26296
rect 13078 26256 13084 26268
rect 13136 26256 13142 26308
rect 9600 26200 10088 26228
rect 4525 26191 4583 26197
rect 13998 26188 14004 26240
rect 14056 26228 14062 26240
rect 14384 26228 14412 26327
rect 14734 26324 14740 26376
rect 14792 26364 14798 26376
rect 15028 26373 15056 26404
rect 15105 26401 15117 26435
rect 15151 26401 15163 26435
rect 15105 26395 15163 26401
rect 16114 26392 16120 26444
rect 16172 26432 16178 26444
rect 16485 26435 16543 26441
rect 16485 26432 16497 26435
rect 16172 26404 16497 26432
rect 16172 26392 16178 26404
rect 16485 26401 16497 26404
rect 16531 26401 16543 26435
rect 16485 26395 16543 26401
rect 16574 26392 16580 26444
rect 16632 26432 16638 26444
rect 16741 26435 16799 26441
rect 16741 26432 16753 26435
rect 16632 26404 16753 26432
rect 16632 26392 16638 26404
rect 16741 26401 16753 26404
rect 16787 26401 16799 26435
rect 16741 26395 16799 26401
rect 20806 26392 20812 26444
rect 20864 26441 20870 26444
rect 20864 26395 20876 26441
rect 20864 26392 20870 26395
rect 14829 26367 14887 26373
rect 14829 26364 14841 26367
rect 14792 26336 14841 26364
rect 14792 26324 14798 26336
rect 14829 26333 14841 26336
rect 14875 26333 14887 26367
rect 14829 26327 14887 26333
rect 15013 26367 15071 26373
rect 15013 26333 15025 26367
rect 15059 26364 15071 26367
rect 15194 26364 15200 26376
rect 15059 26336 15200 26364
rect 15059 26333 15071 26336
rect 15013 26327 15071 26333
rect 15194 26324 15200 26336
rect 15252 26324 15258 26376
rect 21085 26367 21143 26373
rect 21085 26333 21097 26367
rect 21131 26333 21143 26367
rect 21085 26327 21143 26333
rect 17865 26299 17923 26305
rect 17865 26265 17877 26299
rect 17911 26265 17923 26299
rect 17865 26259 17923 26265
rect 16758 26228 16764 26240
rect 14056 26200 16764 26228
rect 14056 26188 14062 26200
rect 16758 26188 16764 26200
rect 16816 26188 16822 26240
rect 16850 26188 16856 26240
rect 16908 26228 16914 26240
rect 17880 26228 17908 26259
rect 19702 26256 19708 26308
rect 19760 26256 19766 26308
rect 18230 26228 18236 26240
rect 16908 26200 18236 26228
rect 16908 26188 16914 26200
rect 18230 26188 18236 26200
rect 18288 26188 18294 26240
rect 20438 26188 20444 26240
rect 20496 26228 20502 26240
rect 21100 26228 21128 26327
rect 20496 26200 21128 26228
rect 20496 26188 20502 26200
rect 552 26138 28428 26160
rect 552 26086 3882 26138
rect 3934 26086 3946 26138
rect 3998 26086 4010 26138
rect 4062 26086 4074 26138
rect 4126 26086 4138 26138
rect 4190 26086 10851 26138
rect 10903 26086 10915 26138
rect 10967 26086 10979 26138
rect 11031 26086 11043 26138
rect 11095 26086 11107 26138
rect 11159 26086 17820 26138
rect 17872 26086 17884 26138
rect 17936 26086 17948 26138
rect 18000 26086 18012 26138
rect 18064 26086 18076 26138
rect 18128 26086 24789 26138
rect 24841 26086 24853 26138
rect 24905 26086 24917 26138
rect 24969 26086 24981 26138
rect 25033 26086 25045 26138
rect 25097 26086 28428 26138
rect 552 26064 28428 26086
rect 3804 25996 5764 26024
rect 3053 25959 3111 25965
rect 3053 25925 3065 25959
rect 3099 25956 3111 25959
rect 3804 25956 3832 25996
rect 3099 25928 3832 25956
rect 3099 25925 3111 25928
rect 3053 25919 3111 25925
rect 3804 25897 3832 25928
rect 3789 25891 3847 25897
rect 2746 25860 3188 25888
rect 1394 25780 1400 25832
rect 1452 25820 1458 25832
rect 1673 25823 1731 25829
rect 1673 25820 1685 25823
rect 1452 25792 1685 25820
rect 1452 25780 1458 25792
rect 1673 25789 1685 25792
rect 1719 25820 1731 25823
rect 2314 25820 2320 25832
rect 1719 25792 2320 25820
rect 1719 25789 1731 25792
rect 1673 25783 1731 25789
rect 2314 25780 2320 25792
rect 2372 25820 2378 25832
rect 2746 25820 2774 25860
rect 2372 25792 2774 25820
rect 2372 25780 2378 25792
rect 1940 25755 1998 25761
rect 1940 25721 1952 25755
rect 1986 25752 1998 25755
rect 2406 25752 2412 25764
rect 1986 25724 2412 25752
rect 1986 25721 1998 25724
rect 1940 25715 1998 25721
rect 2406 25712 2412 25724
rect 2464 25712 2470 25764
rect 3160 25752 3188 25860
rect 3789 25857 3801 25891
rect 3835 25857 3847 25891
rect 3789 25851 3847 25857
rect 5736 25888 5764 25996
rect 5994 25984 6000 26036
rect 6052 25984 6058 26036
rect 6365 26027 6423 26033
rect 6365 25993 6377 26027
rect 6411 26024 6423 26027
rect 6546 26024 6552 26036
rect 6411 25996 6552 26024
rect 6411 25993 6423 25996
rect 6365 25987 6423 25993
rect 6546 25984 6552 25996
rect 6604 25984 6610 26036
rect 7926 25984 7932 26036
rect 7984 26024 7990 26036
rect 8389 26027 8447 26033
rect 8389 26024 8401 26027
rect 7984 25996 8401 26024
rect 7984 25984 7990 25996
rect 8389 25993 8401 25996
rect 8435 25993 8447 26027
rect 8389 25987 8447 25993
rect 11885 26027 11943 26033
rect 11885 25993 11897 26027
rect 11931 25993 11943 26027
rect 11885 25987 11943 25993
rect 6012 25956 6040 25984
rect 6457 25959 6515 25965
rect 6457 25956 6469 25959
rect 6012 25928 6469 25956
rect 6457 25925 6469 25928
rect 6503 25925 6515 25959
rect 6457 25919 6515 25925
rect 5736 25860 6408 25888
rect 4157 25823 4215 25829
rect 4157 25789 4169 25823
rect 4203 25820 4215 25823
rect 5736 25820 5764 25860
rect 5813 25823 5871 25829
rect 5813 25820 5825 25823
rect 4203 25792 4936 25820
rect 5736 25792 5825 25820
rect 4203 25789 4215 25792
rect 4157 25783 4215 25789
rect 4172 25752 4200 25783
rect 3160 25724 4200 25752
rect 4424 25755 4482 25761
rect 4424 25721 4436 25755
rect 4470 25752 4482 25755
rect 4706 25752 4712 25764
rect 4470 25724 4712 25752
rect 4470 25721 4482 25724
rect 4424 25715 4482 25721
rect 4706 25712 4712 25724
rect 4764 25712 4770 25764
rect 4908 25752 4936 25792
rect 5813 25789 5825 25792
rect 5859 25789 5871 25823
rect 5813 25783 5871 25789
rect 6270 25780 6276 25832
rect 6328 25780 6334 25832
rect 6288 25752 6316 25780
rect 4908 25724 6316 25752
rect 6380 25752 6408 25860
rect 6564 25820 6592 25984
rect 6730 25916 6736 25968
rect 6788 25956 6794 25968
rect 6917 25959 6975 25965
rect 6917 25956 6929 25959
rect 6788 25928 6929 25956
rect 6788 25916 6794 25928
rect 6917 25925 6929 25928
rect 6963 25925 6975 25959
rect 6917 25919 6975 25925
rect 7006 25916 7012 25968
rect 7064 25916 7070 25968
rect 10965 25959 11023 25965
rect 10965 25925 10977 25959
rect 11011 25956 11023 25959
rect 11330 25956 11336 25968
rect 11011 25928 11336 25956
rect 11011 25925 11023 25928
rect 10965 25919 11023 25925
rect 11330 25916 11336 25928
rect 11388 25956 11394 25968
rect 11900 25956 11928 25987
rect 12526 25984 12532 26036
rect 12584 25984 12590 26036
rect 13078 25984 13084 26036
rect 13136 25984 13142 26036
rect 15289 26027 15347 26033
rect 15289 25993 15301 26027
rect 15335 26024 15347 26027
rect 16301 26027 16359 26033
rect 15335 25996 16252 26024
rect 15335 25993 15347 25996
rect 15289 25987 15347 25993
rect 13906 25956 13912 25968
rect 11388 25928 13912 25956
rect 11388 25916 11394 25928
rect 13906 25916 13912 25928
rect 13964 25916 13970 25968
rect 6917 25823 6975 25829
rect 6917 25820 6929 25823
rect 6564 25792 6929 25820
rect 6917 25789 6929 25792
rect 6963 25789 6975 25823
rect 7024 25820 7052 25916
rect 11057 25891 11115 25897
rect 11057 25857 11069 25891
rect 11103 25857 11115 25891
rect 14826 25888 14832 25900
rect 11057 25851 11115 25857
rect 11440 25860 12204 25888
rect 7193 25823 7251 25829
rect 7193 25820 7205 25823
rect 7024 25792 7205 25820
rect 6917 25783 6975 25789
rect 7193 25789 7205 25792
rect 7239 25789 7251 25823
rect 7193 25783 7251 25789
rect 7926 25780 7932 25832
rect 7984 25820 7990 25832
rect 8573 25823 8631 25829
rect 8573 25820 8585 25823
rect 7984 25792 8585 25820
rect 7984 25780 7990 25792
rect 8573 25789 8585 25792
rect 8619 25789 8631 25823
rect 8573 25783 8631 25789
rect 8662 25780 8668 25832
rect 8720 25820 8726 25832
rect 8849 25823 8907 25829
rect 8849 25820 8861 25823
rect 8720 25792 8861 25820
rect 8720 25780 8726 25792
rect 8849 25789 8861 25792
rect 8895 25789 8907 25823
rect 11072 25820 11100 25851
rect 11333 25823 11391 25829
rect 11333 25820 11345 25823
rect 11072 25792 11345 25820
rect 8849 25783 8907 25789
rect 11333 25789 11345 25792
rect 11379 25789 11391 25823
rect 11333 25783 11391 25789
rect 6822 25752 6828 25764
rect 6380 25724 6828 25752
rect 6822 25712 6828 25724
rect 6880 25712 6886 25764
rect 7742 25712 7748 25764
rect 7800 25752 7806 25764
rect 10597 25755 10655 25761
rect 10597 25752 10609 25755
rect 7800 25724 10609 25752
rect 7800 25712 7806 25724
rect 10597 25721 10609 25724
rect 10643 25752 10655 25755
rect 11440 25752 11468 25860
rect 12176 25829 12204 25860
rect 12406 25860 14832 25888
rect 11609 25823 11667 25829
rect 11609 25789 11621 25823
rect 11655 25789 11667 25823
rect 11609 25783 11667 25789
rect 12161 25823 12219 25829
rect 12161 25789 12173 25823
rect 12207 25789 12219 25823
rect 12161 25783 12219 25789
rect 10643 25724 11468 25752
rect 11624 25752 11652 25783
rect 12250 25780 12256 25832
rect 12308 25780 12314 25832
rect 12268 25752 12296 25780
rect 11624 25724 12296 25752
rect 10643 25721 10655 25724
rect 10597 25715 10655 25721
rect 3142 25644 3148 25696
rect 3200 25684 3206 25696
rect 3237 25687 3295 25693
rect 3237 25684 3249 25687
rect 3200 25656 3249 25684
rect 3200 25644 3206 25656
rect 3237 25653 3249 25656
rect 3283 25653 3295 25687
rect 3237 25647 3295 25653
rect 5537 25687 5595 25693
rect 5537 25653 5549 25687
rect 5583 25684 5595 25687
rect 5994 25684 6000 25696
rect 5583 25656 6000 25684
rect 5583 25653 5595 25656
rect 5537 25647 5595 25653
rect 5994 25644 6000 25656
rect 6052 25644 6058 25696
rect 6273 25687 6331 25693
rect 6273 25653 6285 25687
rect 6319 25684 6331 25687
rect 6362 25684 6368 25696
rect 6319 25656 6368 25684
rect 6319 25653 6331 25656
rect 6273 25647 6331 25653
rect 6362 25644 6368 25656
rect 6420 25684 6426 25696
rect 7101 25687 7159 25693
rect 7101 25684 7113 25687
rect 6420 25656 7113 25684
rect 6420 25644 6426 25656
rect 7101 25653 7113 25656
rect 7147 25653 7159 25687
rect 7101 25647 7159 25653
rect 8754 25644 8760 25696
rect 8812 25684 8818 25696
rect 11149 25687 11207 25693
rect 11149 25684 11161 25687
rect 8812 25656 11161 25684
rect 8812 25644 8818 25656
rect 11149 25653 11161 25656
rect 11195 25653 11207 25687
rect 11149 25647 11207 25653
rect 11517 25687 11575 25693
rect 11517 25653 11529 25687
rect 11563 25684 11575 25687
rect 11701 25687 11759 25693
rect 11701 25684 11713 25687
rect 11563 25656 11713 25684
rect 11563 25653 11575 25656
rect 11517 25647 11575 25653
rect 11701 25653 11713 25656
rect 11747 25653 11759 25687
rect 11701 25647 11759 25653
rect 11882 25644 11888 25696
rect 11940 25684 11946 25696
rect 12406 25684 12434 25860
rect 14826 25848 14832 25860
rect 14884 25888 14890 25900
rect 15304 25888 15332 25987
rect 15473 25959 15531 25965
rect 15473 25925 15485 25959
rect 15519 25925 15531 25959
rect 16224 25956 16252 25996
rect 16301 25993 16313 26027
rect 16347 26024 16359 26027
rect 16574 26024 16580 26036
rect 16347 25996 16580 26024
rect 16347 25993 16359 25996
rect 16301 25987 16359 25993
rect 16574 25984 16580 25996
rect 16632 25984 16638 26036
rect 20806 25984 20812 26036
rect 20864 26024 20870 26036
rect 20901 26027 20959 26033
rect 20901 26024 20913 26027
rect 20864 25996 20913 26024
rect 20864 25984 20870 25996
rect 20901 25993 20913 25996
rect 20947 25993 20959 26027
rect 20901 25987 20959 25993
rect 18138 25956 18144 25968
rect 16224 25928 18144 25956
rect 15473 25919 15531 25925
rect 14884 25860 15332 25888
rect 14884 25848 14890 25860
rect 12897 25823 12955 25829
rect 12897 25820 12909 25823
rect 12636 25792 12909 25820
rect 12636 25764 12664 25792
rect 12897 25789 12909 25792
rect 12943 25820 12955 25823
rect 12989 25823 13047 25829
rect 12989 25820 13001 25823
rect 12943 25792 13001 25820
rect 12943 25789 12955 25792
rect 12897 25783 12955 25789
rect 12989 25789 13001 25792
rect 13035 25789 13047 25823
rect 12989 25783 13047 25789
rect 13173 25823 13231 25829
rect 13173 25789 13185 25823
rect 13219 25820 13231 25823
rect 13998 25820 14004 25832
rect 13219 25792 14004 25820
rect 13219 25789 13231 25792
rect 13173 25783 13231 25789
rect 12618 25712 12624 25764
rect 12676 25712 12682 25764
rect 12710 25712 12716 25764
rect 12768 25752 12774 25764
rect 13188 25752 13216 25783
rect 13998 25780 14004 25792
rect 14056 25780 14062 25832
rect 14918 25780 14924 25832
rect 14976 25780 14982 25832
rect 15488 25820 15516 25919
rect 18138 25916 18144 25928
rect 18196 25916 18202 25968
rect 20438 25888 20444 25900
rect 20088 25860 20444 25888
rect 16117 25823 16175 25829
rect 16117 25820 16129 25823
rect 15488 25792 16129 25820
rect 16117 25789 16129 25792
rect 16163 25789 16175 25823
rect 16117 25783 16175 25789
rect 18325 25823 18383 25829
rect 18325 25789 18337 25823
rect 18371 25820 18383 25823
rect 18414 25820 18420 25832
rect 18371 25792 18420 25820
rect 18371 25789 18383 25792
rect 18325 25783 18383 25789
rect 18414 25780 18420 25792
rect 18472 25780 18478 25832
rect 19978 25780 19984 25832
rect 20036 25820 20042 25832
rect 20088 25829 20116 25860
rect 20438 25848 20444 25860
rect 20496 25888 20502 25900
rect 21269 25891 21327 25897
rect 21269 25888 21281 25891
rect 20496 25860 21281 25888
rect 20496 25848 20502 25860
rect 21269 25857 21281 25860
rect 21315 25857 21327 25891
rect 21269 25851 21327 25857
rect 20073 25823 20131 25829
rect 20073 25820 20085 25823
rect 20036 25792 20085 25820
rect 20036 25780 20042 25792
rect 20073 25789 20085 25792
rect 20119 25789 20131 25823
rect 20073 25783 20131 25789
rect 20346 25780 20352 25832
rect 20404 25780 20410 25832
rect 21284 25820 21312 25851
rect 22922 25820 22928 25832
rect 21284 25792 22928 25820
rect 22922 25780 22928 25792
rect 22980 25820 22986 25832
rect 23842 25820 23848 25832
rect 22980 25792 23848 25820
rect 22980 25780 22986 25792
rect 23842 25780 23848 25792
rect 23900 25780 23906 25832
rect 19806 25755 19864 25761
rect 19806 25752 19818 25755
rect 12768 25724 13216 25752
rect 18524 25724 19818 25752
rect 12768 25712 12774 25724
rect 11940 25656 12434 25684
rect 11940 25644 11946 25656
rect 15286 25644 15292 25696
rect 15344 25644 15350 25696
rect 18524 25693 18552 25724
rect 19806 25721 19818 25724
rect 19852 25721 19864 25755
rect 19806 25715 19864 25721
rect 21536 25755 21594 25761
rect 21536 25721 21548 25755
rect 21582 25752 21594 25755
rect 21726 25752 21732 25764
rect 21582 25724 21732 25752
rect 21582 25721 21594 25724
rect 21536 25715 21594 25721
rect 21726 25712 21732 25724
rect 21784 25712 21790 25764
rect 18509 25687 18567 25693
rect 18509 25653 18521 25687
rect 18555 25653 18567 25687
rect 18509 25647 18567 25653
rect 18690 25644 18696 25696
rect 18748 25644 18754 25696
rect 22646 25644 22652 25696
rect 22704 25644 22710 25696
rect 552 25594 28587 25616
rect 552 25542 7366 25594
rect 7418 25542 7430 25594
rect 7482 25542 7494 25594
rect 7546 25542 7558 25594
rect 7610 25542 7622 25594
rect 7674 25542 14335 25594
rect 14387 25542 14399 25594
rect 14451 25542 14463 25594
rect 14515 25542 14527 25594
rect 14579 25542 14591 25594
rect 14643 25542 21304 25594
rect 21356 25542 21368 25594
rect 21420 25542 21432 25594
rect 21484 25542 21496 25594
rect 21548 25542 21560 25594
rect 21612 25542 28273 25594
rect 28325 25542 28337 25594
rect 28389 25542 28401 25594
rect 28453 25542 28465 25594
rect 28517 25542 28529 25594
rect 28581 25542 28587 25594
rect 552 25520 28587 25542
rect 2406 25440 2412 25492
rect 2464 25480 2470 25492
rect 2464 25452 2774 25480
rect 2464 25440 2470 25452
rect 2746 25208 2774 25452
rect 3142 25440 3148 25492
rect 3200 25440 3206 25492
rect 3694 25480 3700 25492
rect 3344 25452 3700 25480
rect 3344 25412 3372 25452
rect 3694 25440 3700 25452
rect 3752 25440 3758 25492
rect 3865 25483 3923 25489
rect 3865 25449 3877 25483
rect 3911 25480 3923 25483
rect 4338 25480 4344 25492
rect 3911 25452 4344 25480
rect 3911 25449 3923 25452
rect 3865 25443 3923 25449
rect 4338 25440 4344 25452
rect 4396 25480 4402 25492
rect 4396 25452 4660 25480
rect 4396 25440 4402 25452
rect 3252 25384 3372 25412
rect 3252 25353 3280 25384
rect 2961 25347 3019 25353
rect 2961 25313 2973 25347
rect 3007 25313 3019 25347
rect 2961 25307 3019 25313
rect 3237 25347 3295 25353
rect 3237 25313 3249 25347
rect 3283 25313 3295 25347
rect 3237 25307 3295 25313
rect 2976 25276 3004 25307
rect 3326 25304 3332 25356
rect 3384 25304 3390 25356
rect 3421 25347 3479 25353
rect 3421 25313 3433 25347
rect 3467 25344 3479 25347
rect 3712 25344 3740 25440
rect 4065 25415 4123 25421
rect 4065 25381 4077 25415
rect 4111 25381 4123 25415
rect 4632 25412 4660 25452
rect 4706 25440 4712 25492
rect 4764 25440 4770 25492
rect 7926 25440 7932 25492
rect 7984 25440 7990 25492
rect 8297 25483 8355 25489
rect 8297 25449 8309 25483
rect 8343 25480 8355 25483
rect 8662 25480 8668 25492
rect 8343 25452 8668 25480
rect 8343 25449 8355 25452
rect 8297 25443 8355 25449
rect 8662 25440 8668 25452
rect 8720 25440 8726 25492
rect 8754 25440 8760 25492
rect 8812 25440 8818 25492
rect 8938 25440 8944 25492
rect 8996 25480 9002 25492
rect 9125 25483 9183 25489
rect 9125 25480 9137 25483
rect 8996 25452 9137 25480
rect 8996 25440 9002 25452
rect 9125 25449 9137 25452
rect 9171 25449 9183 25483
rect 9125 25443 9183 25449
rect 12250 25440 12256 25492
rect 12308 25440 12314 25492
rect 13648 25452 14320 25480
rect 4632 25384 5488 25412
rect 4065 25375 4123 25381
rect 4080 25344 4108 25375
rect 5460 25356 5488 25384
rect 8036 25384 8340 25412
rect 3467 25316 3740 25344
rect 3804 25316 4108 25344
rect 3467 25313 3479 25316
rect 3421 25307 3479 25313
rect 3804 25288 3832 25316
rect 4890 25304 4896 25356
rect 4948 25304 4954 25356
rect 5442 25304 5448 25356
rect 5500 25304 5506 25356
rect 8036 25353 8064 25384
rect 8312 25356 8340 25384
rect 7837 25347 7895 25353
rect 7837 25313 7849 25347
rect 7883 25313 7895 25347
rect 7837 25307 7895 25313
rect 8021 25347 8079 25353
rect 8021 25313 8033 25347
rect 8067 25313 8079 25347
rect 8021 25307 8079 25313
rect 8113 25347 8171 25353
rect 8113 25313 8125 25347
rect 8159 25313 8171 25347
rect 8113 25307 8171 25313
rect 3605 25279 3663 25285
rect 2976 25248 3556 25276
rect 3528 25217 3556 25248
rect 3605 25245 3617 25279
rect 3651 25245 3663 25279
rect 3605 25239 3663 25245
rect 2961 25211 3019 25217
rect 2961 25208 2973 25211
rect 2746 25180 2973 25208
rect 2961 25177 2973 25180
rect 3007 25177 3019 25211
rect 2961 25171 3019 25177
rect 3513 25211 3571 25217
rect 3513 25177 3525 25211
rect 3559 25177 3571 25211
rect 3620 25208 3648 25239
rect 3786 25236 3792 25288
rect 3844 25236 3850 25288
rect 6638 25236 6644 25288
rect 6696 25276 6702 25288
rect 7852 25276 7880 25307
rect 8128 25276 8156 25307
rect 8294 25304 8300 25356
rect 8352 25304 8358 25356
rect 8772 25353 8800 25440
rect 11606 25372 11612 25424
rect 11664 25412 11670 25424
rect 13648 25421 13676 25452
rect 13633 25415 13691 25421
rect 13633 25412 13645 25415
rect 11664 25384 13645 25412
rect 11664 25372 11670 25384
rect 13633 25381 13645 25384
rect 13679 25381 13691 25415
rect 13633 25375 13691 25381
rect 13849 25415 13907 25421
rect 13849 25381 13861 25415
rect 13895 25412 13907 25415
rect 13998 25412 14004 25424
rect 13895 25384 14004 25412
rect 13895 25381 13907 25384
rect 13849 25375 13907 25381
rect 13998 25372 14004 25384
rect 14056 25372 14062 25424
rect 14185 25415 14243 25421
rect 14185 25381 14197 25415
rect 14231 25381 14243 25415
rect 14292 25412 14320 25452
rect 14366 25440 14372 25492
rect 14424 25489 14430 25492
rect 14424 25483 14443 25489
rect 14431 25449 14443 25483
rect 14424 25443 14443 25449
rect 14553 25483 14611 25489
rect 14553 25449 14565 25483
rect 14599 25480 14611 25483
rect 14826 25480 14832 25492
rect 14599 25452 14832 25480
rect 14599 25449 14611 25452
rect 14553 25443 14611 25449
rect 14424 25440 14430 25443
rect 14826 25440 14832 25452
rect 14884 25480 14890 25492
rect 14884 25452 14964 25480
rect 14884 25440 14890 25452
rect 14936 25421 14964 25452
rect 15286 25440 15292 25492
rect 15344 25440 15350 25492
rect 18414 25440 18420 25492
rect 18472 25440 18478 25492
rect 21726 25440 21732 25492
rect 21784 25440 21790 25492
rect 14921 25415 14979 25421
rect 14292 25384 14872 25412
rect 14185 25375 14243 25381
rect 8757 25347 8815 25353
rect 8757 25313 8769 25347
rect 8803 25313 8815 25347
rect 12713 25347 12771 25353
rect 12713 25344 12725 25347
rect 8757 25307 8815 25313
rect 12544 25316 12725 25344
rect 12544 25288 12572 25316
rect 12713 25313 12725 25316
rect 12759 25313 12771 25347
rect 12713 25307 12771 25313
rect 13722 25304 13728 25356
rect 13780 25304 13786 25356
rect 6696 25248 8156 25276
rect 6696 25236 6702 25248
rect 8662 25236 8668 25288
rect 8720 25236 8726 25288
rect 12526 25236 12532 25288
rect 12584 25236 12590 25288
rect 13740 25208 13768 25304
rect 14200 25276 14228 25375
rect 14844 25344 14872 25384
rect 14921 25381 14933 25415
rect 14967 25381 14979 25415
rect 14921 25375 14979 25381
rect 15105 25415 15163 25421
rect 15105 25381 15117 25415
rect 15151 25412 15163 25415
rect 16850 25412 16856 25424
rect 15151 25384 16856 25412
rect 15151 25381 15163 25384
rect 15105 25375 15163 25381
rect 15120 25344 15148 25375
rect 16850 25372 16856 25384
rect 16908 25372 16914 25424
rect 18322 25421 18328 25424
rect 18049 25415 18107 25421
rect 18049 25381 18061 25415
rect 18095 25381 18107 25415
rect 18049 25375 18107 25381
rect 18265 25415 18328 25421
rect 18265 25381 18277 25415
rect 18311 25381 18328 25415
rect 18265 25375 18328 25381
rect 14844 25316 15148 25344
rect 16758 25304 16764 25356
rect 16816 25304 16822 25356
rect 18064 25344 18092 25375
rect 18322 25372 18328 25375
rect 18380 25372 18386 25424
rect 18598 25372 18604 25424
rect 18656 25412 18662 25424
rect 18656 25384 21312 25412
rect 18656 25372 18662 25384
rect 19610 25353 19616 25356
rect 18509 25347 18567 25353
rect 18509 25344 18521 25347
rect 18064 25316 18521 25344
rect 18509 25313 18521 25316
rect 18555 25313 18567 25347
rect 18509 25307 18567 25313
rect 19604 25307 19616 25353
rect 19610 25304 19616 25307
rect 19668 25304 19674 25356
rect 21284 25353 21312 25384
rect 23842 25372 23848 25424
rect 23900 25412 23906 25424
rect 23900 25384 24348 25412
rect 23900 25372 23906 25384
rect 21269 25347 21327 25353
rect 21269 25313 21281 25347
rect 21315 25313 21327 25347
rect 21269 25307 21327 25313
rect 14550 25276 14556 25288
rect 3620 25180 13768 25208
rect 13924 25248 14556 25276
rect 3513 25171 3571 25177
rect 3881 25143 3939 25149
rect 3881 25109 3893 25143
rect 3927 25140 3939 25143
rect 4338 25140 4344 25152
rect 3927 25112 4344 25140
rect 3927 25109 3939 25112
rect 3881 25103 3939 25109
rect 4338 25100 4344 25112
rect 4396 25140 4402 25152
rect 5350 25140 5356 25152
rect 4396 25112 5356 25140
rect 4396 25100 4402 25112
rect 5350 25100 5356 25112
rect 5408 25100 5414 25152
rect 5442 25100 5448 25152
rect 5500 25140 5506 25152
rect 9582 25140 9588 25152
rect 5500 25112 9588 25140
rect 5500 25100 5506 25112
rect 9582 25100 9588 25112
rect 9640 25100 9646 25152
rect 12621 25143 12679 25149
rect 12621 25109 12633 25143
rect 12667 25140 12679 25143
rect 12710 25140 12716 25152
rect 12667 25112 12716 25140
rect 12667 25109 12679 25112
rect 12621 25103 12679 25109
rect 12710 25100 12716 25112
rect 12768 25100 12774 25152
rect 13078 25100 13084 25152
rect 13136 25140 13142 25152
rect 13817 25143 13875 25149
rect 13817 25140 13829 25143
rect 13136 25112 13829 25140
rect 13136 25100 13142 25112
rect 13817 25109 13829 25112
rect 13863 25140 13875 25143
rect 13924 25140 13952 25248
rect 14550 25236 14556 25248
rect 14608 25236 14614 25288
rect 14918 25236 14924 25288
rect 14976 25236 14982 25288
rect 16853 25279 16911 25285
rect 16853 25245 16865 25279
rect 16899 25276 16911 25279
rect 18690 25276 18696 25288
rect 16899 25248 18696 25276
rect 16899 25245 16911 25248
rect 16853 25239 16911 25245
rect 18690 25236 18696 25248
rect 18748 25276 18754 25288
rect 19061 25279 19119 25285
rect 19061 25276 19073 25279
rect 18748 25248 19073 25276
rect 18748 25236 18754 25248
rect 19061 25245 19073 25248
rect 19107 25245 19119 25279
rect 19061 25239 19119 25245
rect 19337 25279 19395 25285
rect 19337 25245 19349 25279
rect 19383 25245 19395 25279
rect 21284 25276 21312 25307
rect 21450 25304 21456 25356
rect 21508 25304 21514 25356
rect 21637 25347 21695 25353
rect 21637 25313 21649 25347
rect 21683 25344 21695 25347
rect 21913 25347 21971 25353
rect 21913 25344 21925 25347
rect 21683 25316 21925 25344
rect 21683 25313 21695 25316
rect 21637 25307 21695 25313
rect 21913 25313 21925 25316
rect 21959 25313 21971 25347
rect 21913 25307 21971 25313
rect 24049 25347 24107 25353
rect 24049 25313 24061 25347
rect 24095 25344 24107 25347
rect 24210 25344 24216 25356
rect 24095 25316 24216 25344
rect 24095 25313 24107 25316
rect 24049 25307 24107 25313
rect 24210 25304 24216 25316
rect 24268 25304 24274 25356
rect 24320 25353 24348 25384
rect 24305 25347 24363 25353
rect 24305 25313 24317 25347
rect 24351 25313 24363 25347
rect 24305 25307 24363 25313
rect 23198 25276 23204 25288
rect 21284 25248 23204 25276
rect 19337 25239 19395 25245
rect 14001 25211 14059 25217
rect 14001 25177 14013 25211
rect 14047 25208 14059 25211
rect 14936 25208 14964 25236
rect 14047 25180 14964 25208
rect 14047 25177 14059 25180
rect 14001 25171 14059 25177
rect 13863 25112 13952 25140
rect 13863 25109 13875 25112
rect 13817 25103 13875 25109
rect 14090 25100 14096 25152
rect 14148 25140 14154 25152
rect 14369 25143 14427 25149
rect 14369 25140 14381 25143
rect 14148 25112 14381 25140
rect 14148 25100 14154 25112
rect 14369 25109 14381 25112
rect 14415 25109 14427 25143
rect 14369 25103 14427 25109
rect 17126 25100 17132 25152
rect 17184 25100 17190 25152
rect 18138 25100 18144 25152
rect 18196 25140 18202 25152
rect 18233 25143 18291 25149
rect 18233 25140 18245 25143
rect 18196 25112 18245 25140
rect 18196 25100 18202 25112
rect 18233 25109 18245 25112
rect 18279 25109 18291 25143
rect 19352 25140 19380 25239
rect 23198 25236 23204 25248
rect 23256 25236 23262 25288
rect 19978 25140 19984 25152
rect 19352 25112 19984 25140
rect 18233 25103 18291 25109
rect 19978 25100 19984 25112
rect 20036 25100 20042 25152
rect 20717 25143 20775 25149
rect 20717 25109 20729 25143
rect 20763 25140 20775 25143
rect 20990 25140 20996 25152
rect 20763 25112 20996 25140
rect 20763 25109 20775 25112
rect 20717 25103 20775 25109
rect 20990 25100 20996 25112
rect 21048 25100 21054 25152
rect 22922 25100 22928 25152
rect 22980 25100 22986 25152
rect 552 25050 28428 25072
rect 552 24998 3882 25050
rect 3934 24998 3946 25050
rect 3998 24998 4010 25050
rect 4062 24998 4074 25050
rect 4126 24998 4138 25050
rect 4190 24998 10851 25050
rect 10903 24998 10915 25050
rect 10967 24998 10979 25050
rect 11031 24998 11043 25050
rect 11095 24998 11107 25050
rect 11159 24998 17820 25050
rect 17872 24998 17884 25050
rect 17936 24998 17948 25050
rect 18000 24998 18012 25050
rect 18064 24998 18076 25050
rect 18128 24998 24789 25050
rect 24841 24998 24853 25050
rect 24905 24998 24917 25050
rect 24969 24998 24981 25050
rect 25033 24998 25045 25050
rect 25097 24998 28428 25050
rect 552 24976 28428 24998
rect 6638 24936 6644 24948
rect 6288 24908 6644 24936
rect 3786 24828 3792 24880
rect 3844 24868 3850 24880
rect 6288 24877 6316 24908
rect 6638 24896 6644 24908
rect 6696 24896 6702 24948
rect 7006 24896 7012 24948
rect 7064 24936 7070 24948
rect 7193 24939 7251 24945
rect 7193 24936 7205 24939
rect 7064 24908 7205 24936
rect 7064 24896 7070 24908
rect 7193 24905 7205 24908
rect 7239 24905 7251 24939
rect 7193 24899 7251 24905
rect 9858 24896 9864 24948
rect 9916 24936 9922 24948
rect 10229 24939 10287 24945
rect 10229 24936 10241 24939
rect 9916 24908 10241 24936
rect 9916 24896 9922 24908
rect 10229 24905 10241 24908
rect 10275 24936 10287 24939
rect 11882 24936 11888 24948
rect 10275 24908 11888 24936
rect 10275 24905 10287 24908
rect 10229 24899 10287 24905
rect 11882 24896 11888 24908
rect 11940 24896 11946 24948
rect 12526 24896 12532 24948
rect 12584 24896 12590 24948
rect 14182 24896 14188 24948
rect 14240 24896 14246 24948
rect 14734 24896 14740 24948
rect 14792 24936 14798 24948
rect 15197 24939 15255 24945
rect 15197 24936 15209 24939
rect 14792 24908 15209 24936
rect 14792 24896 14798 24908
rect 15197 24905 15209 24908
rect 15243 24905 15255 24939
rect 15197 24899 15255 24905
rect 18322 24896 18328 24948
rect 18380 24936 18386 24948
rect 18877 24939 18935 24945
rect 18877 24936 18889 24939
rect 18380 24908 18889 24936
rect 18380 24896 18386 24908
rect 18877 24905 18889 24908
rect 18923 24936 18935 24939
rect 19242 24936 19248 24948
rect 18923 24908 19248 24936
rect 18923 24905 18935 24908
rect 18877 24899 18935 24905
rect 19242 24896 19248 24908
rect 19300 24896 19306 24948
rect 19610 24896 19616 24948
rect 19668 24896 19674 24948
rect 21450 24896 21456 24948
rect 21508 24936 21514 24948
rect 21545 24939 21603 24945
rect 21545 24936 21557 24939
rect 21508 24908 21557 24936
rect 21508 24896 21514 24908
rect 21545 24905 21557 24908
rect 21591 24905 21603 24939
rect 21545 24899 21603 24905
rect 22465 24939 22523 24945
rect 22465 24905 22477 24939
rect 22511 24936 22523 24939
rect 22646 24936 22652 24948
rect 22511 24908 22652 24936
rect 22511 24905 22523 24908
rect 22465 24899 22523 24905
rect 22646 24896 22652 24908
rect 22704 24896 22710 24948
rect 6273 24871 6331 24877
rect 6273 24868 6285 24871
rect 3844 24840 6285 24868
rect 3844 24828 3850 24840
rect 6273 24837 6285 24840
rect 6319 24837 6331 24871
rect 6273 24831 6331 24837
rect 11698 24828 11704 24880
rect 11756 24868 11762 24880
rect 12544 24868 12572 24896
rect 11756 24840 12572 24868
rect 11756 24828 11762 24840
rect 6457 24803 6515 24809
rect 6457 24769 6469 24803
rect 6503 24800 6515 24803
rect 7009 24803 7067 24809
rect 6503 24772 6868 24800
rect 6503 24769 6515 24772
rect 6457 24763 6515 24769
rect 6549 24735 6607 24741
rect 6549 24701 6561 24735
rect 6595 24701 6607 24735
rect 6840 24732 6868 24772
rect 7009 24769 7021 24803
rect 7055 24800 7067 24803
rect 7101 24803 7159 24809
rect 7101 24800 7113 24803
rect 7055 24772 7113 24800
rect 7055 24769 7067 24772
rect 7009 24763 7067 24769
rect 7101 24769 7113 24772
rect 7147 24769 7159 24803
rect 10505 24803 10563 24809
rect 10505 24800 10517 24803
rect 7101 24763 7159 24769
rect 9508 24772 10517 24800
rect 9508 24744 9536 24772
rect 10505 24769 10517 24772
rect 10551 24769 10563 24803
rect 10505 24763 10563 24769
rect 12342 24760 12348 24812
rect 12400 24760 12406 24812
rect 14200 24800 14228 24896
rect 14826 24828 14832 24880
rect 14884 24828 14890 24880
rect 13924 24772 14228 24800
rect 15304 24772 16068 24800
rect 13924 24744 13952 24772
rect 7285 24735 7343 24741
rect 7285 24732 7297 24735
rect 6840 24704 7297 24732
rect 6549 24695 6607 24701
rect 7285 24701 7297 24704
rect 7331 24701 7343 24735
rect 7285 24695 7343 24701
rect 7377 24735 7435 24741
rect 7377 24701 7389 24735
rect 7423 24701 7435 24735
rect 7377 24695 7435 24701
rect 5902 24624 5908 24676
rect 5960 24664 5966 24676
rect 5997 24667 6055 24673
rect 5997 24664 6009 24667
rect 5960 24636 6009 24664
rect 5960 24624 5966 24636
rect 5997 24633 6009 24636
rect 6043 24664 6055 24667
rect 6564 24664 6592 24695
rect 6043 24636 6592 24664
rect 6043 24633 6055 24636
rect 5997 24627 6055 24633
rect 7282 24556 7288 24608
rect 7340 24596 7346 24608
rect 7392 24596 7420 24695
rect 9490 24692 9496 24744
rect 9548 24692 9554 24744
rect 9582 24692 9588 24744
rect 9640 24732 9646 24744
rect 9861 24735 9919 24741
rect 9861 24732 9873 24735
rect 9640 24704 9873 24732
rect 9640 24692 9646 24704
rect 9861 24701 9873 24704
rect 9907 24701 9919 24735
rect 9861 24695 9919 24701
rect 11054 24692 11060 24744
rect 11112 24732 11118 24744
rect 12618 24732 12624 24744
rect 11112 24704 12624 24732
rect 11112 24692 11118 24704
rect 12618 24692 12624 24704
rect 12676 24692 12682 24744
rect 12710 24692 12716 24744
rect 12768 24732 12774 24744
rect 12805 24735 12863 24741
rect 12805 24732 12817 24735
rect 12768 24704 12817 24732
rect 12768 24692 12774 24704
rect 12805 24701 12817 24704
rect 12851 24701 12863 24735
rect 12805 24695 12863 24701
rect 13906 24692 13912 24744
rect 13964 24692 13970 24744
rect 13998 24692 14004 24744
rect 14056 24732 14062 24744
rect 14369 24735 14427 24741
rect 14369 24732 14381 24735
rect 14056 24704 14381 24732
rect 14056 24692 14062 24704
rect 14369 24701 14381 24704
rect 14415 24701 14427 24735
rect 14369 24695 14427 24701
rect 10229 24667 10287 24673
rect 10229 24633 10241 24667
rect 10275 24664 10287 24667
rect 10594 24664 10600 24676
rect 10275 24636 10600 24664
rect 10275 24633 10287 24636
rect 10229 24627 10287 24633
rect 10594 24624 10600 24636
rect 10652 24624 10658 24676
rect 10778 24673 10784 24676
rect 10772 24627 10784 24673
rect 10778 24624 10784 24627
rect 10836 24624 10842 24676
rect 14090 24624 14096 24676
rect 14148 24624 14154 24676
rect 14550 24624 14556 24676
rect 14608 24664 14614 24676
rect 15304 24664 15332 24772
rect 15933 24735 15991 24741
rect 15933 24732 15945 24735
rect 14608 24636 15332 24664
rect 15396 24704 15945 24732
rect 14608 24624 14614 24636
rect 7340 24568 7420 24596
rect 7340 24556 7346 24568
rect 10410 24556 10416 24608
rect 10468 24556 10474 24608
rect 10962 24556 10968 24608
rect 11020 24596 11026 24608
rect 11698 24596 11704 24608
rect 11020 24568 11704 24596
rect 11020 24556 11026 24568
rect 11698 24556 11704 24568
rect 11756 24596 11762 24608
rect 11885 24599 11943 24605
rect 11885 24596 11897 24599
rect 11756 24568 11897 24596
rect 11756 24556 11762 24568
rect 11885 24565 11897 24568
rect 11931 24565 11943 24599
rect 11885 24559 11943 24565
rect 14182 24556 14188 24608
rect 14240 24596 14246 24608
rect 15396 24605 15424 24704
rect 15933 24701 15945 24704
rect 15979 24701 15991 24735
rect 16040 24732 16068 24772
rect 16114 24760 16120 24812
rect 16172 24800 16178 24812
rect 16209 24803 16267 24809
rect 16209 24800 16221 24803
rect 16172 24772 16221 24800
rect 16172 24760 16178 24772
rect 16209 24769 16221 24772
rect 16255 24769 16267 24803
rect 16209 24763 16267 24769
rect 20806 24760 20812 24812
rect 20864 24800 20870 24812
rect 20901 24803 20959 24809
rect 20901 24800 20913 24803
rect 20864 24772 20913 24800
rect 20864 24760 20870 24772
rect 20901 24769 20913 24772
rect 20947 24769 20959 24803
rect 20901 24763 20959 24769
rect 22002 24760 22008 24812
rect 22060 24800 22066 24812
rect 22649 24803 22707 24809
rect 22649 24800 22661 24803
rect 22060 24772 22661 24800
rect 22060 24760 22066 24772
rect 22649 24769 22661 24772
rect 22695 24769 22707 24803
rect 22649 24763 22707 24769
rect 19797 24735 19855 24741
rect 19797 24732 19809 24735
rect 16040 24704 17632 24732
rect 15933 24695 15991 24701
rect 16454 24667 16512 24673
rect 16454 24664 16466 24667
rect 16132 24636 16466 24664
rect 16132 24605 16160 24636
rect 16454 24633 16466 24636
rect 16500 24633 16512 24667
rect 16454 24627 16512 24633
rect 17604 24605 17632 24704
rect 19076 24704 19809 24732
rect 18138 24624 18144 24676
rect 18196 24664 18202 24676
rect 18693 24667 18751 24673
rect 18693 24664 18705 24667
rect 18196 24636 18705 24664
rect 18196 24624 18202 24636
rect 18693 24633 18705 24636
rect 18739 24633 18751 24667
rect 18693 24627 18751 24633
rect 14277 24599 14335 24605
rect 14277 24596 14289 24599
rect 14240 24568 14289 24596
rect 14240 24556 14246 24568
rect 14277 24565 14289 24568
rect 14323 24565 14335 24599
rect 14277 24559 14335 24565
rect 14737 24599 14795 24605
rect 14737 24565 14749 24599
rect 14783 24596 14795 24599
rect 15197 24599 15255 24605
rect 15197 24596 15209 24599
rect 14783 24568 15209 24596
rect 14783 24565 14795 24568
rect 14737 24559 14795 24565
rect 15197 24565 15209 24568
rect 15243 24565 15255 24599
rect 15197 24559 15255 24565
rect 15381 24599 15439 24605
rect 15381 24565 15393 24599
rect 15427 24565 15439 24599
rect 15381 24559 15439 24565
rect 16117 24599 16175 24605
rect 16117 24565 16129 24599
rect 16163 24565 16175 24599
rect 16117 24559 16175 24565
rect 17589 24599 17647 24605
rect 17589 24565 17601 24599
rect 17635 24596 17647 24599
rect 18506 24596 18512 24608
rect 17635 24568 18512 24596
rect 17635 24565 17647 24568
rect 17589 24559 17647 24565
rect 18506 24556 18512 24568
rect 18564 24556 18570 24608
rect 18782 24556 18788 24608
rect 18840 24596 18846 24608
rect 19076 24605 19104 24704
rect 19797 24701 19809 24704
rect 19843 24701 19855 24735
rect 19797 24695 19855 24701
rect 21818 24692 21824 24744
rect 21876 24732 21882 24744
rect 22373 24735 22431 24741
rect 22373 24732 22385 24735
rect 21876 24704 22385 24732
rect 21876 24692 21882 24704
rect 22373 24701 22385 24704
rect 22419 24701 22431 24735
rect 22373 24695 22431 24701
rect 19337 24667 19395 24673
rect 19337 24633 19349 24667
rect 19383 24633 19395 24667
rect 19337 24627 19395 24633
rect 19521 24667 19579 24673
rect 19521 24633 19533 24667
rect 19567 24664 19579 24667
rect 19610 24664 19616 24676
rect 19567 24636 19616 24664
rect 19567 24633 19579 24636
rect 19521 24627 19579 24633
rect 18893 24599 18951 24605
rect 18893 24596 18905 24599
rect 18840 24568 18905 24596
rect 18840 24556 18846 24568
rect 18893 24565 18905 24568
rect 18939 24565 18951 24599
rect 18893 24559 18951 24565
rect 19061 24599 19119 24605
rect 19061 24565 19073 24599
rect 19107 24565 19119 24599
rect 19061 24559 19119 24565
rect 19153 24599 19211 24605
rect 19153 24565 19165 24599
rect 19199 24596 19211 24599
rect 19242 24596 19248 24608
rect 19199 24568 19248 24596
rect 19199 24565 19211 24568
rect 19153 24559 19211 24565
rect 19242 24556 19248 24568
rect 19300 24556 19306 24608
rect 19352 24596 19380 24627
rect 19610 24624 19616 24636
rect 19668 24664 19674 24676
rect 21177 24667 21235 24673
rect 21177 24664 21189 24667
rect 19668 24636 21189 24664
rect 19668 24624 19674 24636
rect 21177 24633 21189 24636
rect 21223 24633 21235 24667
rect 21177 24627 21235 24633
rect 19426 24596 19432 24608
rect 19352 24568 19432 24596
rect 19426 24556 19432 24568
rect 19484 24596 19490 24608
rect 20622 24596 20628 24608
rect 19484 24568 20628 24596
rect 19484 24556 19490 24568
rect 20622 24556 20628 24568
rect 20680 24556 20686 24608
rect 21082 24556 21088 24608
rect 21140 24556 21146 24608
rect 22646 24556 22652 24608
rect 22704 24556 22710 24608
rect 552 24506 28587 24528
rect 552 24454 7366 24506
rect 7418 24454 7430 24506
rect 7482 24454 7494 24506
rect 7546 24454 7558 24506
rect 7610 24454 7622 24506
rect 7674 24454 14335 24506
rect 14387 24454 14399 24506
rect 14451 24454 14463 24506
rect 14515 24454 14527 24506
rect 14579 24454 14591 24506
rect 14643 24454 21304 24506
rect 21356 24454 21368 24506
rect 21420 24454 21432 24506
rect 21484 24454 21496 24506
rect 21548 24454 21560 24506
rect 21612 24454 28273 24506
rect 28325 24454 28337 24506
rect 28389 24454 28401 24506
rect 28453 24454 28465 24506
rect 28517 24454 28529 24506
rect 28581 24454 28587 24506
rect 552 24432 28587 24454
rect 4341 24395 4399 24401
rect 4341 24361 4353 24395
rect 4387 24392 4399 24395
rect 4801 24395 4859 24401
rect 4801 24392 4813 24395
rect 4387 24364 4813 24392
rect 4387 24361 4399 24364
rect 4341 24355 4399 24361
rect 4801 24361 4813 24364
rect 4847 24361 4859 24395
rect 4801 24355 4859 24361
rect 1504 24296 2774 24324
rect 1302 24216 1308 24268
rect 1360 24216 1366 24268
rect 1394 24148 1400 24200
rect 1452 24188 1458 24200
rect 1504 24197 1532 24296
rect 1756 24259 1814 24265
rect 1756 24225 1768 24259
rect 1802 24256 1814 24259
rect 2130 24256 2136 24268
rect 1802 24228 2136 24256
rect 1802 24225 1814 24228
rect 1756 24219 1814 24225
rect 2130 24216 2136 24228
rect 2188 24216 2194 24268
rect 2746 24256 2774 24296
rect 2961 24259 3019 24265
rect 2961 24256 2973 24259
rect 2746 24228 2973 24256
rect 2961 24225 2973 24228
rect 3007 24225 3019 24259
rect 2961 24219 3019 24225
rect 3228 24259 3286 24265
rect 3228 24225 3240 24259
rect 3274 24256 3286 24259
rect 3510 24256 3516 24268
rect 3274 24228 3516 24256
rect 3274 24225 3286 24228
rect 3228 24219 3286 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 3694 24216 3700 24268
rect 3752 24256 3758 24268
rect 4617 24259 4675 24265
rect 4617 24256 4629 24259
rect 3752 24228 4629 24256
rect 3752 24216 3758 24228
rect 4617 24225 4629 24228
rect 4663 24225 4675 24259
rect 4617 24219 4675 24225
rect 4709 24259 4767 24265
rect 4709 24225 4721 24259
rect 4755 24225 4767 24259
rect 4816 24256 4844 24355
rect 5350 24352 5356 24404
rect 5408 24392 5414 24404
rect 7742 24392 7748 24404
rect 5408 24364 7748 24392
rect 5408 24352 5414 24364
rect 6932 24333 6960 24364
rect 7742 24352 7748 24364
rect 7800 24352 7806 24404
rect 8297 24395 8355 24401
rect 8297 24361 8309 24395
rect 8343 24392 8355 24395
rect 8662 24392 8668 24404
rect 8343 24364 8668 24392
rect 8343 24361 8355 24364
rect 8297 24355 8355 24361
rect 8662 24352 8668 24364
rect 8720 24352 8726 24404
rect 9214 24352 9220 24404
rect 9272 24392 9278 24404
rect 9743 24395 9801 24401
rect 9743 24392 9755 24395
rect 9272 24364 9755 24392
rect 9272 24352 9278 24364
rect 9743 24361 9755 24364
rect 9789 24361 9801 24395
rect 9743 24355 9801 24361
rect 10410 24352 10416 24404
rect 10468 24352 10474 24404
rect 10594 24352 10600 24404
rect 10652 24352 10658 24404
rect 10689 24395 10747 24401
rect 10689 24361 10701 24395
rect 10735 24392 10747 24395
rect 10778 24392 10784 24404
rect 10735 24364 10784 24392
rect 10735 24361 10747 24364
rect 10689 24355 10747 24361
rect 10778 24352 10784 24364
rect 10836 24352 10842 24404
rect 10965 24395 11023 24401
rect 10965 24361 10977 24395
rect 11011 24361 11023 24395
rect 10965 24355 11023 24361
rect 6917 24327 6975 24333
rect 6012 24296 6776 24324
rect 5169 24259 5227 24265
rect 5169 24256 5181 24259
rect 4816 24228 5181 24256
rect 4709 24219 4767 24225
rect 5169 24225 5181 24228
rect 5215 24225 5227 24259
rect 5169 24219 5227 24225
rect 1489 24191 1547 24197
rect 1489 24188 1501 24191
rect 1452 24160 1501 24188
rect 1452 24148 1458 24160
rect 1489 24157 1501 24160
rect 1535 24157 1547 24191
rect 1489 24151 1547 24157
rect 4433 24123 4491 24129
rect 4433 24089 4445 24123
rect 4479 24089 4491 24123
rect 4724 24120 4752 24219
rect 5350 24148 5356 24200
rect 5408 24188 5414 24200
rect 5902 24188 5908 24200
rect 5408 24160 5908 24188
rect 5408 24148 5414 24160
rect 5902 24148 5908 24160
rect 5960 24188 5966 24200
rect 6012 24197 6040 24296
rect 6181 24259 6239 24265
rect 6181 24225 6193 24259
rect 6227 24256 6239 24259
rect 6362 24256 6368 24268
rect 6227 24228 6368 24256
rect 6227 24225 6239 24228
rect 6181 24219 6239 24225
rect 6362 24216 6368 24228
rect 6420 24256 6426 24268
rect 6420 24228 6684 24256
rect 6420 24216 6426 24228
rect 5997 24191 6055 24197
rect 5997 24188 6009 24191
rect 5960 24160 6009 24188
rect 5960 24148 5966 24160
rect 5997 24157 6009 24160
rect 6043 24157 6055 24191
rect 5997 24151 6055 24157
rect 6089 24191 6147 24197
rect 6089 24157 6101 24191
rect 6135 24157 6147 24191
rect 6273 24191 6331 24197
rect 6273 24188 6285 24191
rect 6089 24151 6147 24157
rect 6196 24160 6285 24188
rect 4724 24092 6040 24120
rect 4433 24083 4491 24089
rect 1118 24012 1124 24064
rect 1176 24012 1182 24064
rect 2869 24055 2927 24061
rect 2869 24021 2881 24055
rect 2915 24052 2927 24055
rect 4246 24052 4252 24064
rect 2915 24024 4252 24052
rect 2915 24021 2927 24024
rect 2869 24015 2927 24021
rect 4246 24012 4252 24024
rect 4304 24052 4310 24064
rect 4448 24052 4476 24083
rect 6012 24064 6040 24092
rect 6104 24064 6132 24151
rect 6196 24132 6224 24160
rect 6273 24157 6285 24160
rect 6319 24157 6331 24191
rect 6273 24151 6331 24157
rect 6178 24080 6184 24132
rect 6236 24080 6242 24132
rect 6656 24129 6684 24228
rect 6748 24188 6776 24296
rect 6917 24293 6929 24327
rect 6963 24293 6975 24327
rect 6917 24287 6975 24293
rect 9953 24327 10011 24333
rect 9953 24293 9965 24327
rect 9999 24293 10011 24327
rect 9953 24287 10011 24293
rect 7285 24259 7343 24265
rect 7285 24225 7297 24259
rect 7331 24256 7343 24259
rect 7742 24256 7748 24268
rect 7331 24228 7748 24256
rect 7331 24225 7343 24228
rect 7285 24219 7343 24225
rect 7742 24216 7748 24228
rect 7800 24216 7806 24268
rect 7929 24259 7987 24265
rect 7929 24225 7941 24259
rect 7975 24225 7987 24259
rect 7929 24219 7987 24225
rect 9493 24259 9551 24265
rect 9493 24225 9505 24259
rect 9539 24256 9551 24259
rect 9968 24256 9996 24287
rect 9539 24228 9996 24256
rect 10428 24256 10456 24352
rect 10612 24324 10640 24352
rect 10980 24324 11008 24355
rect 11146 24352 11152 24404
rect 11204 24392 11210 24404
rect 12986 24392 12992 24404
rect 11204 24364 12992 24392
rect 11204 24352 11210 24364
rect 12986 24352 12992 24364
rect 13044 24352 13050 24404
rect 13906 24352 13912 24404
rect 13964 24352 13970 24404
rect 13998 24352 14004 24404
rect 14056 24392 14062 24404
rect 14093 24395 14151 24401
rect 14093 24392 14105 24395
rect 14056 24364 14105 24392
rect 14056 24352 14062 24364
rect 14093 24361 14105 24364
rect 14139 24361 14151 24395
rect 14093 24355 14151 24361
rect 10612 24296 11008 24324
rect 11532 24296 11744 24324
rect 10505 24259 10563 24265
rect 10505 24256 10517 24259
rect 10428 24228 10517 24256
rect 9539 24225 9551 24228
rect 9493 24219 9551 24225
rect 7193 24191 7251 24197
rect 7193 24188 7205 24191
rect 6748 24160 7205 24188
rect 7193 24157 7205 24160
rect 7239 24157 7251 24191
rect 7193 24151 7251 24157
rect 7653 24191 7711 24197
rect 7653 24157 7665 24191
rect 7699 24188 7711 24191
rect 7837 24191 7895 24197
rect 7837 24188 7849 24191
rect 7699 24160 7849 24188
rect 7699 24157 7711 24160
rect 7653 24151 7711 24157
rect 7837 24157 7849 24160
rect 7883 24157 7895 24191
rect 7837 24151 7895 24157
rect 6641 24123 6699 24129
rect 6288 24092 6592 24120
rect 4304 24024 4476 24052
rect 4985 24055 5043 24061
rect 4304 24012 4310 24024
rect 4985 24021 4997 24055
rect 5031 24052 5043 24055
rect 5258 24052 5264 24064
rect 5031 24024 5264 24052
rect 5031 24021 5043 24024
rect 4985 24015 5043 24021
rect 5258 24012 5264 24024
rect 5316 24012 5322 24064
rect 5350 24012 5356 24064
rect 5408 24012 5414 24064
rect 5810 24012 5816 24064
rect 5868 24012 5874 24064
rect 5994 24012 6000 24064
rect 6052 24012 6058 24064
rect 6086 24012 6092 24064
rect 6144 24052 6150 24064
rect 6288 24052 6316 24092
rect 6144 24024 6316 24052
rect 6144 24012 6150 24024
rect 6454 24012 6460 24064
rect 6512 24012 6518 24064
rect 6564 24052 6592 24092
rect 6641 24089 6653 24123
rect 6687 24089 6699 24123
rect 6641 24083 6699 24089
rect 7282 24080 7288 24132
rect 7340 24120 7346 24132
rect 7944 24120 7972 24219
rect 9968 24188 9996 24228
rect 10505 24225 10517 24228
rect 10551 24225 10563 24259
rect 10505 24219 10563 24225
rect 11242 24262 11300 24265
rect 11532 24262 11560 24296
rect 11242 24259 11560 24262
rect 11242 24225 11254 24259
rect 11288 24234 11560 24259
rect 11288 24225 11300 24234
rect 11242 24219 11300 24225
rect 11606 24216 11612 24268
rect 11664 24216 11670 24268
rect 10962 24188 10968 24200
rect 9968 24160 10968 24188
rect 10962 24148 10968 24160
rect 11020 24148 11026 24200
rect 11054 24148 11060 24200
rect 11112 24148 11118 24200
rect 11146 24148 11152 24200
rect 11204 24148 11210 24200
rect 11333 24191 11391 24197
rect 11333 24157 11345 24191
rect 11379 24157 11391 24191
rect 11333 24151 11391 24157
rect 11425 24191 11483 24197
rect 11425 24157 11437 24191
rect 11471 24157 11483 24191
rect 11716 24188 11744 24296
rect 11790 24216 11796 24268
rect 11848 24256 11854 24268
rect 12437 24259 12495 24265
rect 12437 24256 12449 24259
rect 11848 24228 12449 24256
rect 11848 24216 11854 24228
rect 12437 24225 12449 24228
rect 12483 24225 12495 24259
rect 12437 24219 12495 24225
rect 12529 24259 12587 24265
rect 12529 24225 12541 24259
rect 12575 24256 12587 24259
rect 13078 24256 13084 24268
rect 12575 24228 13084 24256
rect 12575 24225 12587 24228
rect 12529 24219 12587 24225
rect 13078 24216 13084 24228
rect 13136 24216 13142 24268
rect 13924 24265 13952 24352
rect 13909 24259 13967 24265
rect 13909 24225 13921 24259
rect 13955 24225 13967 24259
rect 14108 24256 14136 24355
rect 14182 24352 14188 24404
rect 14240 24392 14246 24404
rect 14645 24395 14703 24401
rect 14645 24392 14657 24395
rect 14240 24364 14657 24392
rect 14240 24352 14246 24364
rect 14645 24361 14657 24364
rect 14691 24361 14703 24395
rect 14645 24355 14703 24361
rect 15381 24395 15439 24401
rect 15381 24361 15393 24395
rect 15427 24361 15439 24395
rect 15381 24355 15439 24361
rect 15396 24324 15424 24355
rect 15562 24352 15568 24404
rect 15620 24392 15626 24404
rect 15620 24364 18736 24392
rect 15620 24352 15626 24364
rect 16362 24327 16420 24333
rect 16362 24324 16374 24327
rect 15396 24296 16374 24324
rect 16362 24293 16374 24296
rect 16408 24293 16420 24327
rect 16362 24287 16420 24293
rect 18248 24296 18644 24324
rect 14277 24259 14335 24265
rect 14277 24256 14289 24259
rect 14108 24228 14289 24256
rect 13909 24219 13967 24225
rect 14277 24225 14289 24228
rect 14323 24225 14335 24259
rect 15197 24259 15255 24265
rect 15197 24256 15209 24259
rect 14277 24219 14335 24225
rect 14844 24228 15209 24256
rect 12066 24188 12072 24200
rect 11716 24160 12072 24188
rect 11425 24151 11483 24157
rect 7340 24092 7972 24120
rect 8036 24092 9444 24120
rect 7340 24080 7346 24092
rect 7742 24052 7748 24064
rect 6564 24024 7748 24052
rect 7742 24012 7748 24024
rect 7800 24052 7806 24064
rect 8036 24052 8064 24092
rect 7800 24024 8064 24052
rect 7800 24012 7806 24024
rect 9030 24012 9036 24064
rect 9088 24012 9094 24064
rect 9416 24061 9444 24092
rect 9582 24080 9588 24132
rect 9640 24080 9646 24132
rect 11072 24120 11100 24148
rect 9692 24092 11100 24120
rect 9401 24055 9459 24061
rect 9401 24021 9413 24055
rect 9447 24052 9459 24055
rect 9692 24052 9720 24092
rect 9447 24024 9720 24052
rect 9447 24021 9459 24024
rect 9401 24015 9459 24021
rect 9766 24012 9772 24064
rect 9824 24052 9830 24064
rect 10686 24052 10692 24064
rect 9824 24024 10692 24052
rect 9824 24012 9830 24024
rect 10686 24012 10692 24024
rect 10744 24052 10750 24064
rect 11348 24052 11376 24151
rect 11440 24120 11468 24151
rect 12066 24148 12072 24160
rect 12124 24148 12130 24200
rect 12802 24148 12808 24200
rect 12860 24188 12866 24200
rect 13725 24191 13783 24197
rect 13725 24188 13737 24191
rect 12860 24160 13737 24188
rect 12860 24148 12866 24160
rect 13725 24157 13737 24160
rect 13771 24188 13783 24191
rect 14090 24188 14096 24200
rect 13771 24160 14096 24188
rect 13771 24157 13783 24160
rect 13725 24151 13783 24157
rect 14090 24148 14096 24160
rect 14148 24188 14154 24200
rect 14148 24160 14780 24188
rect 14148 24148 14154 24160
rect 11698 24120 11704 24132
rect 11440 24092 11704 24120
rect 11698 24080 11704 24092
rect 11756 24080 11762 24132
rect 10744 24024 11376 24052
rect 10744 24012 10750 24024
rect 11790 24012 11796 24064
rect 11848 24012 11854 24064
rect 13906 24012 13912 24064
rect 13964 24052 13970 24064
rect 14642 24052 14648 24064
rect 13964 24024 14648 24052
rect 13964 24012 13970 24024
rect 14642 24012 14648 24024
rect 14700 24012 14706 24064
rect 14752 24052 14780 24160
rect 14844 24129 14872 24228
rect 15197 24225 15209 24228
rect 15243 24225 15255 24259
rect 15197 24219 15255 24225
rect 16114 24216 16120 24268
rect 16172 24216 16178 24268
rect 17957 24259 18015 24265
rect 17957 24225 17969 24259
rect 18003 24256 18015 24259
rect 18046 24256 18052 24268
rect 18003 24228 18052 24256
rect 18003 24225 18015 24228
rect 17957 24219 18015 24225
rect 18046 24216 18052 24228
rect 18104 24216 18110 24268
rect 18248 24265 18276 24296
rect 18616 24268 18644 24296
rect 18141 24259 18199 24265
rect 18141 24225 18153 24259
rect 18187 24225 18199 24259
rect 18141 24219 18199 24225
rect 18233 24259 18291 24265
rect 18233 24225 18245 24259
rect 18279 24225 18291 24259
rect 18233 24219 18291 24225
rect 18156 24188 18184 24219
rect 18506 24216 18512 24268
rect 18564 24216 18570 24268
rect 18598 24216 18604 24268
rect 18656 24216 18662 24268
rect 18708 24256 18736 24364
rect 18782 24352 18788 24404
rect 18840 24352 18846 24404
rect 18969 24395 19027 24401
rect 18969 24361 18981 24395
rect 19015 24392 19027 24395
rect 19981 24395 20039 24401
rect 19981 24392 19993 24395
rect 19015 24364 19993 24392
rect 19015 24361 19027 24364
rect 18969 24355 19027 24361
rect 19981 24361 19993 24364
rect 20027 24361 20039 24395
rect 19981 24355 20039 24361
rect 20441 24395 20499 24401
rect 20441 24361 20453 24395
rect 20487 24392 20499 24395
rect 22462 24392 22468 24404
rect 20487 24364 22468 24392
rect 20487 24361 20499 24364
rect 20441 24355 20499 24361
rect 22462 24352 22468 24364
rect 22520 24352 22526 24404
rect 22646 24352 22652 24404
rect 22704 24352 22710 24404
rect 22020 24296 22600 24324
rect 18910 24259 18968 24265
rect 18910 24256 18922 24259
rect 18708 24228 18922 24256
rect 18910 24225 18922 24228
rect 18956 24225 18968 24259
rect 18910 24219 18968 24225
rect 20346 24216 20352 24268
rect 20404 24216 20410 24268
rect 21634 24216 21640 24268
rect 21692 24256 21698 24268
rect 22020 24265 22048 24296
rect 22572 24268 22600 24296
rect 22005 24259 22063 24265
rect 22005 24256 22017 24259
rect 21692 24228 22017 24256
rect 21692 24216 21698 24228
rect 22005 24225 22017 24228
rect 22051 24225 22063 24259
rect 22005 24219 22063 24225
rect 22097 24259 22155 24265
rect 22097 24225 22109 24259
rect 22143 24225 22155 24259
rect 22281 24259 22339 24265
rect 22281 24256 22293 24259
rect 22097 24219 22155 24225
rect 22204 24228 22293 24256
rect 18782 24188 18788 24200
rect 18156 24160 18788 24188
rect 18782 24148 18788 24160
rect 18840 24148 18846 24200
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24188 19487 24191
rect 19610 24188 19616 24200
rect 19475 24160 19616 24188
rect 19475 24157 19487 24160
rect 19429 24151 19487 24157
rect 19610 24148 19616 24160
rect 19668 24148 19674 24200
rect 20530 24148 20536 24200
rect 20588 24148 20594 24200
rect 14829 24123 14887 24129
rect 14829 24089 14841 24123
rect 14875 24089 14887 24123
rect 19337 24123 19395 24129
rect 19337 24120 19349 24123
rect 14829 24083 14887 24089
rect 17696 24092 19349 24120
rect 17696 24064 17724 24092
rect 19337 24089 19349 24092
rect 19383 24120 19395 24123
rect 20990 24120 20996 24132
rect 19383 24092 20996 24120
rect 19383 24089 19395 24092
rect 19337 24083 19395 24089
rect 20990 24080 20996 24092
rect 21048 24120 21054 24132
rect 21818 24120 21824 24132
rect 21048 24092 21824 24120
rect 21048 24080 21054 24092
rect 21818 24080 21824 24092
rect 21876 24120 21882 24132
rect 22112 24120 22140 24219
rect 22204 24200 22232 24228
rect 22281 24225 22293 24228
rect 22327 24225 22339 24259
rect 22281 24219 22339 24225
rect 22554 24216 22560 24268
rect 22612 24216 22618 24268
rect 22664 24256 22692 24352
rect 23216 24296 23428 24324
rect 23216 24268 23244 24296
rect 23109 24259 23167 24265
rect 23109 24256 23121 24259
rect 22664 24228 23121 24256
rect 23109 24225 23121 24228
rect 23155 24225 23167 24259
rect 23109 24219 23167 24225
rect 23198 24216 23204 24268
rect 23256 24216 23262 24268
rect 23400 24265 23428 24296
rect 23293 24259 23351 24265
rect 23293 24225 23305 24259
rect 23339 24225 23351 24259
rect 23293 24219 23351 24225
rect 23385 24259 23443 24265
rect 23385 24225 23397 24259
rect 23431 24225 23443 24259
rect 23385 24219 23443 24225
rect 22186 24148 22192 24200
rect 22244 24188 22250 24200
rect 22649 24191 22707 24197
rect 22649 24188 22661 24191
rect 22244 24160 22661 24188
rect 22244 24148 22250 24160
rect 22649 24157 22661 24160
rect 22695 24157 22707 24191
rect 22649 24151 22707 24157
rect 22925 24123 22983 24129
rect 21876 24092 22600 24120
rect 21876 24080 21882 24092
rect 17034 24052 17040 24064
rect 14752 24024 17040 24052
rect 17034 24012 17040 24024
rect 17092 24052 17098 24064
rect 17497 24055 17555 24061
rect 17497 24052 17509 24055
rect 17092 24024 17509 24052
rect 17092 24012 17098 24024
rect 17497 24021 17509 24024
rect 17543 24021 17555 24055
rect 17497 24015 17555 24021
rect 17678 24012 17684 24064
rect 17736 24012 17742 24064
rect 18322 24012 18328 24064
rect 18380 24012 18386 24064
rect 18414 24012 18420 24064
rect 18472 24012 18478 24064
rect 22462 24012 22468 24064
rect 22520 24012 22526 24064
rect 22572 24061 22600 24092
rect 22925 24089 22937 24123
rect 22971 24120 22983 24123
rect 23106 24120 23112 24132
rect 22971 24092 23112 24120
rect 22971 24089 22983 24092
rect 22925 24083 22983 24089
rect 23106 24080 23112 24092
rect 23164 24120 23170 24132
rect 23308 24120 23336 24219
rect 23566 24216 23572 24268
rect 23624 24216 23630 24268
rect 24112 24259 24170 24265
rect 24112 24225 24124 24259
rect 24158 24256 24170 24259
rect 24486 24256 24492 24268
rect 24158 24228 24492 24256
rect 24158 24225 24170 24228
rect 24112 24219 24170 24225
rect 24486 24216 24492 24228
rect 24544 24216 24550 24268
rect 23842 24148 23848 24200
rect 23900 24148 23906 24200
rect 23164 24092 23336 24120
rect 23164 24080 23170 24092
rect 22557 24055 22615 24061
rect 22557 24021 22569 24055
rect 22603 24021 22615 24055
rect 22557 24015 22615 24021
rect 23198 24012 23204 24064
rect 23256 24012 23262 24064
rect 23753 24055 23811 24061
rect 23753 24021 23765 24055
rect 23799 24052 23811 24055
rect 24210 24052 24216 24064
rect 23799 24024 24216 24052
rect 23799 24021 23811 24024
rect 23753 24015 23811 24021
rect 24210 24012 24216 24024
rect 24268 24012 24274 24064
rect 24578 24012 24584 24064
rect 24636 24052 24642 24064
rect 25225 24055 25283 24061
rect 25225 24052 25237 24055
rect 24636 24024 25237 24052
rect 24636 24012 24642 24024
rect 25225 24021 25237 24024
rect 25271 24021 25283 24055
rect 25225 24015 25283 24021
rect 552 23962 28428 23984
rect 552 23910 3882 23962
rect 3934 23910 3946 23962
rect 3998 23910 4010 23962
rect 4062 23910 4074 23962
rect 4126 23910 4138 23962
rect 4190 23910 10851 23962
rect 10903 23910 10915 23962
rect 10967 23910 10979 23962
rect 11031 23910 11043 23962
rect 11095 23910 11107 23962
rect 11159 23910 17820 23962
rect 17872 23910 17884 23962
rect 17936 23910 17948 23962
rect 18000 23910 18012 23962
rect 18064 23910 18076 23962
rect 18128 23910 24789 23962
rect 24841 23910 24853 23962
rect 24905 23910 24917 23962
rect 24969 23910 24981 23962
rect 25033 23910 25045 23962
rect 25097 23910 28428 23962
rect 552 23888 28428 23910
rect 2130 23808 2136 23860
rect 2188 23848 2194 23860
rect 2685 23851 2743 23857
rect 2685 23848 2697 23851
rect 2188 23820 2697 23848
rect 2188 23808 2194 23820
rect 2685 23817 2697 23820
rect 2731 23817 2743 23851
rect 2685 23811 2743 23817
rect 3694 23808 3700 23860
rect 3752 23808 3758 23860
rect 4246 23808 4252 23860
rect 4304 23808 4310 23860
rect 4801 23851 4859 23857
rect 4801 23817 4813 23851
rect 4847 23848 4859 23851
rect 4890 23848 4896 23860
rect 4847 23820 4896 23848
rect 4847 23817 4859 23820
rect 4801 23811 4859 23817
rect 4890 23808 4896 23820
rect 4948 23808 4954 23860
rect 4985 23851 5043 23857
rect 4985 23817 4997 23851
rect 5031 23848 5043 23851
rect 5810 23848 5816 23860
rect 5031 23820 5816 23848
rect 5031 23817 5043 23820
rect 4985 23811 5043 23817
rect 5810 23808 5816 23820
rect 5868 23808 5874 23860
rect 6086 23808 6092 23860
rect 6144 23808 6150 23860
rect 6457 23851 6515 23857
rect 6457 23817 6469 23851
rect 6503 23848 6515 23851
rect 7282 23848 7288 23860
rect 6503 23820 7288 23848
rect 6503 23817 6515 23820
rect 6457 23811 6515 23817
rect 7282 23808 7288 23820
rect 7340 23808 7346 23860
rect 9030 23808 9036 23860
rect 9088 23808 9094 23860
rect 9122 23808 9128 23860
rect 9180 23848 9186 23860
rect 11514 23848 11520 23860
rect 9180 23820 11520 23848
rect 9180 23808 9186 23820
rect 11514 23808 11520 23820
rect 11572 23808 11578 23860
rect 12710 23808 12716 23860
rect 12768 23848 12774 23860
rect 14090 23848 14096 23860
rect 12768 23820 14096 23848
rect 12768 23808 12774 23820
rect 14090 23808 14096 23820
rect 14148 23808 14154 23860
rect 15654 23808 15660 23860
rect 15712 23848 15718 23860
rect 16114 23848 16120 23860
rect 15712 23820 16120 23848
rect 15712 23808 15718 23820
rect 16114 23808 16120 23820
rect 16172 23808 16178 23860
rect 19978 23808 19984 23860
rect 20036 23808 20042 23860
rect 20530 23808 20536 23860
rect 20588 23808 20594 23860
rect 23566 23808 23572 23860
rect 23624 23848 23630 23860
rect 23845 23851 23903 23857
rect 23845 23848 23857 23851
rect 23624 23820 23857 23848
rect 23624 23808 23630 23820
rect 23845 23817 23857 23820
rect 23891 23817 23903 23851
rect 23845 23811 23903 23817
rect 24210 23808 24216 23860
rect 24268 23808 24274 23860
rect 24486 23808 24492 23860
rect 24544 23808 24550 23860
rect 2225 23783 2283 23789
rect 2225 23749 2237 23783
rect 2271 23749 2283 23783
rect 2225 23743 2283 23749
rect 2240 23712 2268 23743
rect 3712 23712 3740 23808
rect 4264 23712 4292 23808
rect 6104 23712 6132 23808
rect 9048 23712 9076 23808
rect 9214 23740 9220 23792
rect 9272 23780 9278 23792
rect 15562 23780 15568 23792
rect 9272 23752 15568 23780
rect 9272 23740 9278 23752
rect 15562 23740 15568 23752
rect 15620 23740 15626 23792
rect 16758 23740 16764 23792
rect 16816 23780 16822 23792
rect 17678 23780 17684 23792
rect 16816 23752 17684 23780
rect 16816 23740 16822 23752
rect 17678 23740 17684 23752
rect 17736 23780 17742 23792
rect 17736 23752 17816 23780
rect 17736 23740 17742 23752
rect 9766 23712 9772 23724
rect 2240 23684 3740 23712
rect 4080 23684 4292 23712
rect 4356 23684 6132 23712
rect 6196 23684 9076 23712
rect 9140 23684 9772 23712
rect 845 23647 903 23653
rect 845 23613 857 23647
rect 891 23644 903 23647
rect 1394 23644 1400 23656
rect 891 23616 1400 23644
rect 891 23613 903 23616
rect 845 23607 903 23613
rect 1118 23585 1124 23588
rect 1112 23576 1124 23585
rect 1079 23548 1124 23576
rect 1112 23539 1124 23548
rect 1118 23536 1124 23539
rect 1176 23536 1182 23588
rect 1228 23520 1256 23616
rect 1394 23604 1400 23616
rect 1452 23604 1458 23656
rect 2608 23653 2636 23684
rect 2593 23647 2651 23653
rect 2593 23613 2605 23647
rect 2639 23644 2651 23647
rect 2639 23616 2673 23644
rect 2639 23613 2651 23616
rect 2593 23607 2651 23613
rect 2866 23604 2872 23656
rect 2924 23604 2930 23656
rect 4080 23653 4108 23684
rect 4065 23647 4123 23653
rect 4065 23613 4077 23647
rect 4111 23613 4123 23647
rect 4065 23607 4123 23613
rect 4157 23647 4215 23653
rect 4157 23613 4169 23647
rect 4203 23644 4215 23647
rect 4246 23644 4252 23656
rect 4203 23616 4252 23644
rect 4203 23613 4215 23616
rect 4157 23607 4215 23613
rect 4246 23604 4252 23616
rect 4304 23604 4310 23656
rect 3694 23536 3700 23588
rect 3752 23576 3758 23588
rect 4356 23576 4384 23684
rect 5258 23604 5264 23656
rect 5316 23644 5322 23656
rect 6196 23653 6224 23684
rect 5353 23647 5411 23653
rect 5353 23644 5365 23647
rect 5316 23616 5365 23644
rect 5316 23604 5322 23616
rect 5353 23613 5365 23616
rect 5399 23613 5411 23647
rect 5353 23607 5411 23613
rect 6181 23647 6239 23653
rect 6181 23613 6193 23647
rect 6227 23613 6239 23647
rect 6181 23607 6239 23613
rect 6454 23604 6460 23656
rect 6512 23604 6518 23656
rect 9030 23604 9036 23656
rect 9088 23644 9094 23656
rect 9140 23653 9168 23684
rect 9766 23672 9772 23684
rect 9824 23672 9830 23724
rect 12986 23672 12992 23724
rect 13044 23712 13050 23724
rect 13814 23712 13820 23724
rect 13044 23684 13820 23712
rect 13044 23672 13050 23684
rect 13814 23672 13820 23684
rect 13872 23712 13878 23724
rect 13872 23684 14044 23712
rect 13872 23672 13878 23684
rect 9125 23647 9183 23653
rect 9125 23644 9137 23647
rect 9088 23616 9137 23644
rect 9088 23604 9094 23616
rect 9125 23613 9137 23616
rect 9171 23613 9183 23647
rect 9125 23607 9183 23613
rect 9214 23604 9220 23656
rect 9272 23644 9278 23656
rect 9309 23647 9367 23653
rect 9309 23644 9321 23647
rect 9272 23616 9321 23644
rect 9272 23604 9278 23616
rect 9309 23613 9321 23616
rect 9355 23613 9367 23647
rect 9309 23607 9367 23613
rect 9398 23604 9404 23656
rect 9456 23604 9462 23656
rect 12345 23647 12403 23653
rect 12345 23613 12357 23647
rect 12391 23644 12403 23647
rect 12537 23649 12595 23655
rect 12391 23616 12425 23644
rect 12391 23613 12403 23616
rect 12345 23607 12403 23613
rect 12537 23615 12549 23649
rect 12583 23644 12595 23649
rect 13078 23644 13084 23656
rect 12583 23616 13084 23644
rect 12583 23615 12595 23616
rect 12537 23609 12595 23615
rect 6273 23579 6331 23585
rect 6273 23576 6285 23579
rect 3752 23548 4384 23576
rect 4632 23548 6285 23576
rect 3752 23536 3758 23548
rect 1210 23468 1216 23520
rect 1268 23468 1274 23520
rect 2406 23468 2412 23520
rect 2464 23468 2470 23520
rect 3602 23468 3608 23520
rect 3660 23508 3666 23520
rect 4632 23517 4660 23548
rect 6273 23545 6285 23548
rect 6319 23545 6331 23579
rect 6273 23539 6331 23545
rect 7834 23536 7840 23588
rect 7892 23576 7898 23588
rect 12360 23576 12388 23607
rect 13078 23604 13084 23616
rect 13136 23604 13142 23656
rect 14016 23653 14044 23684
rect 16960 23684 17633 23712
rect 14001 23647 14059 23653
rect 14001 23613 14013 23647
rect 14047 23613 14059 23647
rect 14001 23607 14059 23613
rect 12802 23576 12808 23588
rect 7892 23548 12808 23576
rect 7892 23536 7898 23548
rect 12802 23536 12808 23548
rect 12860 23536 12866 23588
rect 12986 23536 12992 23588
rect 13044 23576 13050 23588
rect 16850 23576 16856 23588
rect 13044 23548 16856 23576
rect 13044 23536 13050 23548
rect 16850 23536 16856 23548
rect 16908 23576 16914 23588
rect 16960 23576 16988 23684
rect 17126 23604 17132 23656
rect 17184 23644 17190 23656
rect 17605 23653 17633 23684
rect 17788 23653 17816 23752
rect 22388 23752 24164 23780
rect 18782 23672 18788 23724
rect 18840 23712 18846 23724
rect 20806 23712 20812 23724
rect 18840 23684 20812 23712
rect 18840 23672 18846 23684
rect 20806 23672 20812 23684
rect 20864 23712 20870 23724
rect 21634 23712 21640 23724
rect 20864 23684 21640 23712
rect 20864 23672 20870 23684
rect 21634 23672 21640 23684
rect 21692 23672 21698 23724
rect 22388 23712 22416 23752
rect 22204 23684 22416 23712
rect 17497 23647 17555 23653
rect 17497 23644 17509 23647
rect 17184 23616 17509 23644
rect 17184 23604 17190 23616
rect 17497 23613 17509 23616
rect 17543 23613 17555 23647
rect 17497 23607 17555 23613
rect 17590 23647 17648 23653
rect 17590 23613 17602 23647
rect 17636 23613 17648 23647
rect 17590 23607 17648 23613
rect 17773 23647 17831 23653
rect 17773 23613 17785 23647
rect 17819 23613 17831 23647
rect 17773 23607 17831 23613
rect 18003 23647 18061 23653
rect 18003 23613 18015 23647
rect 18049 23644 18061 23647
rect 18966 23644 18972 23656
rect 18049 23616 18972 23644
rect 18049 23613 18061 23616
rect 18003 23607 18061 23613
rect 18966 23604 18972 23616
rect 19024 23604 19030 23656
rect 20901 23647 20959 23653
rect 20901 23613 20913 23647
rect 20947 23644 20959 23647
rect 20990 23644 20996 23656
rect 20947 23616 20996 23644
rect 20947 23613 20959 23616
rect 20901 23607 20959 23613
rect 20990 23604 20996 23616
rect 21048 23644 21054 23656
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 21048 23616 21833 23644
rect 21048 23604 21054 23616
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 21821 23607 21879 23613
rect 21910 23604 21916 23656
rect 21968 23644 21974 23656
rect 22204 23653 22232 23684
rect 22462 23672 22468 23724
rect 22520 23712 22526 23724
rect 22520 23684 22600 23712
rect 22520 23672 22526 23684
rect 22189 23647 22247 23653
rect 21968 23616 22094 23644
rect 21968 23604 21974 23616
rect 16908 23548 16988 23576
rect 16908 23536 16914 23548
rect 17402 23536 17408 23588
rect 17460 23536 17466 23588
rect 17862 23536 17868 23588
rect 17920 23536 17926 23588
rect 18693 23579 18751 23585
rect 18693 23576 18705 23579
rect 17972 23548 18705 23576
rect 3881 23511 3939 23517
rect 3881 23508 3893 23511
rect 3660 23480 3893 23508
rect 3660 23468 3666 23480
rect 3881 23477 3893 23480
rect 3927 23477 3939 23511
rect 3881 23471 3939 23477
rect 4617 23511 4675 23517
rect 4617 23477 4629 23511
rect 4663 23477 4675 23511
rect 4617 23471 4675 23477
rect 4985 23511 5043 23517
rect 4985 23477 4997 23511
rect 5031 23508 5043 23511
rect 8846 23508 8852 23520
rect 5031 23480 8852 23508
rect 5031 23477 5043 23480
rect 4985 23471 5043 23477
rect 8846 23468 8852 23480
rect 8904 23468 8910 23520
rect 8938 23468 8944 23520
rect 8996 23468 9002 23520
rect 9585 23511 9643 23517
rect 9585 23477 9597 23511
rect 9631 23508 9643 23511
rect 9674 23508 9680 23520
rect 9631 23480 9680 23508
rect 9631 23477 9643 23480
rect 9585 23471 9643 23477
rect 9674 23468 9680 23480
rect 9732 23468 9738 23520
rect 11606 23468 11612 23520
rect 11664 23508 11670 23520
rect 12250 23508 12256 23520
rect 11664 23480 12256 23508
rect 11664 23468 11670 23480
rect 12250 23468 12256 23480
rect 12308 23468 12314 23520
rect 12526 23468 12532 23520
rect 12584 23508 12590 23520
rect 13630 23508 13636 23520
rect 12584 23480 13636 23508
rect 12584 23468 12590 23480
rect 13630 23468 13636 23480
rect 13688 23468 13694 23520
rect 14182 23468 14188 23520
rect 14240 23468 14246 23520
rect 17420 23508 17448 23536
rect 17972 23508 18000 23548
rect 18693 23545 18705 23548
rect 18739 23545 18751 23579
rect 22066 23576 22094 23616
rect 22189 23613 22201 23647
rect 22235 23613 22247 23647
rect 22189 23607 22247 23613
rect 22204 23576 22232 23607
rect 22370 23604 22376 23656
rect 22428 23604 22434 23656
rect 22572 23653 22600 23684
rect 22557 23647 22615 23653
rect 22557 23613 22569 23647
rect 22603 23613 22615 23647
rect 22557 23607 22615 23613
rect 22925 23647 22983 23653
rect 22925 23613 22937 23647
rect 22971 23644 22983 23647
rect 23198 23644 23204 23656
rect 22971 23616 23204 23644
rect 22971 23613 22983 23616
rect 22925 23607 22983 23613
rect 23198 23604 23204 23616
rect 23256 23604 23262 23656
rect 23382 23604 23388 23656
rect 23440 23644 23446 23656
rect 24136 23653 24164 23752
rect 24228 23712 24256 23808
rect 24228 23684 24716 23712
rect 24029 23647 24087 23653
rect 24029 23644 24041 23647
rect 23440 23616 24041 23644
rect 23440 23604 23446 23616
rect 24029 23613 24041 23616
rect 24075 23613 24087 23647
rect 24029 23607 24087 23613
rect 24121 23647 24179 23653
rect 24121 23613 24133 23647
rect 24167 23644 24179 23647
rect 24167 23616 24348 23644
rect 24167 23613 24179 23616
rect 24121 23607 24179 23613
rect 22741 23579 22799 23585
rect 22741 23576 22753 23579
rect 22066 23548 22232 23576
rect 22572 23548 22753 23576
rect 18693 23539 18751 23545
rect 22572 23520 22600 23548
rect 22741 23545 22753 23548
rect 22787 23545 22799 23579
rect 22741 23539 22799 23545
rect 22833 23579 22891 23585
rect 22833 23545 22845 23579
rect 22879 23545 22891 23579
rect 24213 23579 24271 23585
rect 22833 23539 22891 23545
rect 23124 23548 24072 23576
rect 17420 23480 18000 23508
rect 18138 23468 18144 23520
rect 18196 23468 18202 23520
rect 22465 23511 22523 23517
rect 22465 23477 22477 23511
rect 22511 23508 22523 23511
rect 22554 23508 22560 23520
rect 22511 23480 22560 23508
rect 22511 23477 22523 23480
rect 22465 23471 22523 23477
rect 22554 23468 22560 23480
rect 22612 23468 22618 23520
rect 22646 23468 22652 23520
rect 22704 23508 22710 23520
rect 22848 23508 22876 23539
rect 23124 23517 23152 23548
rect 22704 23480 22876 23508
rect 23109 23511 23167 23517
rect 22704 23468 22710 23480
rect 23109 23477 23121 23511
rect 23155 23477 23167 23511
rect 24044 23508 24072 23548
rect 24213 23545 24225 23579
rect 24259 23545 24271 23579
rect 24320 23576 24348 23616
rect 24394 23604 24400 23656
rect 24452 23604 24458 23656
rect 24578 23604 24584 23656
rect 24636 23604 24642 23656
rect 24688 23653 24716 23684
rect 24673 23647 24731 23653
rect 24673 23613 24685 23647
rect 24719 23613 24731 23647
rect 24673 23607 24731 23613
rect 24596 23576 24624 23604
rect 24320 23548 24624 23576
rect 24213 23539 24271 23545
rect 24228 23508 24256 23539
rect 24044 23480 24256 23508
rect 23109 23471 23167 23477
rect 552 23418 28587 23440
rect 552 23366 7366 23418
rect 7418 23366 7430 23418
rect 7482 23366 7494 23418
rect 7546 23366 7558 23418
rect 7610 23366 7622 23418
rect 7674 23366 14335 23418
rect 14387 23366 14399 23418
rect 14451 23366 14463 23418
rect 14515 23366 14527 23418
rect 14579 23366 14591 23418
rect 14643 23366 21304 23418
rect 21356 23366 21368 23418
rect 21420 23366 21432 23418
rect 21484 23366 21496 23418
rect 21548 23366 21560 23418
rect 21612 23366 28273 23418
rect 28325 23366 28337 23418
rect 28389 23366 28401 23418
rect 28453 23366 28465 23418
rect 28517 23366 28529 23418
rect 28581 23366 28587 23418
rect 552 23344 28587 23366
rect 1121 23307 1179 23313
rect 1121 23273 1133 23307
rect 1167 23304 1179 23307
rect 1302 23304 1308 23316
rect 1167 23276 1308 23304
rect 1167 23273 1179 23276
rect 1121 23267 1179 23273
rect 1302 23264 1308 23276
rect 1360 23264 1366 23316
rect 3421 23307 3479 23313
rect 3421 23273 3433 23307
rect 3467 23273 3479 23307
rect 3421 23267 3479 23273
rect 1762 23196 1768 23248
rect 1820 23196 1826 23248
rect 1981 23239 2039 23245
rect 1981 23205 1993 23239
rect 2027 23236 2039 23239
rect 2130 23236 2136 23248
rect 2027 23208 2136 23236
rect 2027 23205 2039 23208
rect 1981 23199 2039 23205
rect 2130 23196 2136 23208
rect 2188 23196 2194 23248
rect 3053 23239 3111 23245
rect 3053 23205 3065 23239
rect 3099 23205 3111 23239
rect 3053 23199 3111 23205
rect 1581 23103 1639 23109
rect 1581 23069 1593 23103
rect 1627 23100 1639 23103
rect 2406 23100 2412 23112
rect 1627 23072 2412 23100
rect 1627 23069 1639 23072
rect 1581 23063 1639 23069
rect 2406 23060 2412 23072
rect 2464 23060 2470 23112
rect 3068 23100 3096 23199
rect 3234 23196 3240 23248
rect 3292 23245 3298 23248
rect 3292 23239 3311 23245
rect 3299 23205 3311 23239
rect 3292 23199 3311 23205
rect 3292 23196 3298 23199
rect 3436 23168 3464 23267
rect 3510 23264 3516 23316
rect 3568 23264 3574 23316
rect 8849 23307 8907 23313
rect 8849 23273 8861 23307
rect 8895 23304 8907 23307
rect 9141 23307 9199 23313
rect 9141 23304 9153 23307
rect 8895 23276 9153 23304
rect 8895 23273 8907 23276
rect 8849 23267 8907 23273
rect 9141 23273 9153 23276
rect 9187 23273 9199 23307
rect 9141 23267 9199 23273
rect 9309 23307 9367 23313
rect 9309 23273 9321 23307
rect 9355 23304 9367 23307
rect 9398 23304 9404 23316
rect 9355 23276 9404 23304
rect 9355 23273 9367 23276
rect 9309 23267 9367 23273
rect 9398 23264 9404 23276
rect 9456 23264 9462 23316
rect 9508 23276 10640 23304
rect 4522 23236 4528 23248
rect 4172 23208 4528 23236
rect 3697 23171 3755 23177
rect 3697 23168 3709 23171
rect 3436 23140 3709 23168
rect 3697 23137 3709 23140
rect 3743 23137 3755 23171
rect 3697 23131 3755 23137
rect 4172 23100 4200 23208
rect 4522 23196 4528 23208
rect 4580 23236 4586 23248
rect 8754 23236 8760 23248
rect 4580 23208 8760 23236
rect 4580 23196 4586 23208
rect 8754 23196 8760 23208
rect 8812 23236 8818 23248
rect 8941 23239 8999 23245
rect 8941 23236 8953 23239
rect 8812 23208 8953 23236
rect 8812 23196 8818 23208
rect 8941 23205 8953 23208
rect 8987 23205 8999 23239
rect 8941 23199 8999 23205
rect 9030 23196 9036 23248
rect 9088 23196 9094 23248
rect 9508 23236 9536 23276
rect 9674 23245 9680 23248
rect 9668 23236 9680 23245
rect 9140 23208 9536 23236
rect 9635 23208 9680 23236
rect 4430 23128 4436 23180
rect 4488 23128 4494 23180
rect 4614 23128 4620 23180
rect 4672 23168 4678 23180
rect 5350 23168 5356 23180
rect 4672 23140 5356 23168
rect 4672 23128 4678 23140
rect 5350 23128 5356 23140
rect 5408 23128 5414 23180
rect 6638 23128 6644 23180
rect 6696 23128 6702 23180
rect 7834 23128 7840 23180
rect 7892 23168 7898 23180
rect 8389 23171 8447 23177
rect 8389 23168 8401 23171
rect 7892 23140 8401 23168
rect 7892 23128 7898 23140
rect 8389 23137 8401 23140
rect 8435 23137 8447 23171
rect 8389 23131 8447 23137
rect 8662 23128 8668 23180
rect 8720 23128 8726 23180
rect 8849 23171 8907 23177
rect 8849 23137 8861 23171
rect 8895 23168 8907 23171
rect 9048 23168 9076 23196
rect 8895 23140 9076 23168
rect 8895 23137 8907 23140
rect 8849 23131 8907 23137
rect 3068 23072 4200 23100
rect 6730 23060 6736 23112
rect 6788 23060 6794 23112
rect 8294 23060 8300 23112
rect 8352 23100 8358 23112
rect 9140 23100 9168 23208
rect 9668 23199 9680 23208
rect 9674 23196 9680 23199
rect 9732 23196 9738 23248
rect 9401 23171 9459 23177
rect 9401 23137 9413 23171
rect 9447 23168 9459 23171
rect 9490 23168 9496 23180
rect 9447 23140 9496 23168
rect 9447 23137 9459 23140
rect 9401 23131 9459 23137
rect 9490 23128 9496 23140
rect 9548 23128 9554 23180
rect 10612 23168 10640 23276
rect 10686 23264 10692 23316
rect 10744 23304 10750 23316
rect 10781 23307 10839 23313
rect 10781 23304 10793 23307
rect 10744 23276 10793 23304
rect 10744 23264 10750 23276
rect 10781 23273 10793 23276
rect 10827 23273 10839 23307
rect 10781 23267 10839 23273
rect 11330 23264 11336 23316
rect 11388 23304 11394 23316
rect 11882 23304 11888 23316
rect 11388 23276 11888 23304
rect 11388 23264 11394 23276
rect 11882 23264 11888 23276
rect 11940 23264 11946 23316
rect 12986 23304 12992 23316
rect 11992 23276 12992 23304
rect 11124 23239 11182 23245
rect 11124 23205 11136 23239
rect 11170 23236 11182 23239
rect 11348 23236 11376 23264
rect 11992 23236 12020 23276
rect 12986 23264 12992 23276
rect 13044 23264 13050 23316
rect 13081 23307 13139 23313
rect 13081 23273 13093 23307
rect 13127 23273 13139 23307
rect 13081 23267 13139 23273
rect 13096 23236 13124 23267
rect 13814 23264 13820 23316
rect 13872 23264 13878 23316
rect 13998 23304 14004 23316
rect 13924 23276 14004 23304
rect 13924 23245 13952 23276
rect 13998 23264 14004 23276
rect 14056 23264 14062 23316
rect 14090 23264 14096 23316
rect 14148 23304 14154 23316
rect 17313 23307 17371 23313
rect 14148 23276 14596 23304
rect 14148 23264 14154 23276
rect 13909 23239 13967 23245
rect 11170 23208 11376 23236
rect 11716 23208 12020 23236
rect 12048 23208 12572 23236
rect 13096 23208 13216 23236
rect 11170 23205 11182 23208
rect 11124 23199 11182 23205
rect 11241 23171 11299 23177
rect 11241 23168 11253 23171
rect 10612 23140 11253 23168
rect 11241 23137 11253 23140
rect 11287 23168 11299 23171
rect 11716 23168 11744 23208
rect 11287 23140 11744 23168
rect 11287 23137 11299 23140
rect 11241 23131 11299 23137
rect 11790 23128 11796 23180
rect 11848 23168 11854 23180
rect 12048 23177 12076 23208
rect 12544 23180 12572 23208
rect 11885 23171 11943 23177
rect 11885 23168 11897 23171
rect 11848 23140 11897 23168
rect 11848 23128 11854 23140
rect 11885 23137 11897 23140
rect 11931 23137 11943 23171
rect 11885 23131 11943 23137
rect 12033 23171 12091 23177
rect 12033 23137 12045 23171
rect 12079 23137 12091 23171
rect 12033 23131 12091 23137
rect 12158 23128 12164 23180
rect 12216 23128 12222 23180
rect 12250 23128 12256 23180
rect 12308 23128 12314 23180
rect 12342 23128 12348 23180
rect 12400 23177 12406 23180
rect 12400 23171 12447 23177
rect 12400 23137 12401 23171
rect 12435 23137 12447 23171
rect 12400 23131 12447 23137
rect 12400 23128 12406 23131
rect 12526 23128 12532 23180
rect 12584 23128 12590 23180
rect 12894 23177 12900 23180
rect 12621 23171 12679 23177
rect 12621 23137 12633 23171
rect 12667 23137 12679 23171
rect 12621 23131 12679 23137
rect 12890 23131 12900 23177
rect 12952 23168 12958 23180
rect 12952 23140 12990 23168
rect 8352 23072 9168 23100
rect 8352 23060 8358 23072
rect 11330 23060 11336 23112
rect 11388 23060 11394 23112
rect 11609 23103 11667 23109
rect 11609 23069 11621 23103
rect 11655 23100 11667 23103
rect 11698 23100 11704 23112
rect 11655 23072 11704 23100
rect 11655 23069 11667 23072
rect 11609 23063 11667 23069
rect 11698 23060 11704 23072
rect 11756 23060 11762 23112
rect 12625 23044 12653 23131
rect 12894 23128 12900 23131
rect 12952 23128 12958 23140
rect 13078 23128 13084 23180
rect 13136 23128 13142 23180
rect 13188 23177 13216 23208
rect 13909 23205 13921 23239
rect 13955 23205 13967 23239
rect 13909 23199 13967 23205
rect 13179 23171 13237 23177
rect 13179 23137 13191 23171
rect 13225 23137 13237 23171
rect 13179 23131 13237 23137
rect 13354 23128 13360 23180
rect 13412 23168 13418 23180
rect 14568 23177 14596 23276
rect 17313 23273 17325 23307
rect 17359 23304 17371 23307
rect 17862 23304 17868 23316
rect 17359 23276 17868 23304
rect 17359 23273 17371 23276
rect 17313 23267 17371 23273
rect 14921 23239 14979 23245
rect 14921 23205 14933 23239
rect 14967 23236 14979 23239
rect 15010 23236 15016 23248
rect 14967 23208 15016 23236
rect 14967 23205 14979 23208
rect 14921 23199 14979 23205
rect 15010 23196 15016 23208
rect 15068 23196 15074 23248
rect 15105 23239 15163 23245
rect 15105 23205 15117 23239
rect 15151 23236 15163 23239
rect 15286 23236 15292 23248
rect 15151 23208 15292 23236
rect 15151 23205 15163 23208
rect 15105 23199 15163 23205
rect 15286 23196 15292 23208
rect 15344 23196 15350 23248
rect 15562 23196 15568 23248
rect 15620 23196 15626 23248
rect 17328 23236 17356 23267
rect 17862 23264 17868 23276
rect 17920 23264 17926 23316
rect 18417 23307 18475 23313
rect 18417 23273 18429 23307
rect 18463 23273 18475 23307
rect 18417 23267 18475 23273
rect 17144 23208 17356 23236
rect 18049 23239 18107 23245
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 13412 23140 13553 23168
rect 13412 23128 13418 23140
rect 13541 23137 13553 23140
rect 13587 23137 13599 23171
rect 14369 23171 14427 23177
rect 13541 23131 13599 23137
rect 13648 23140 13892 23168
rect 12805 23103 12863 23109
rect 12805 23069 12817 23103
rect 12851 23100 12863 23103
rect 13096 23100 13124 23128
rect 13648 23100 13676 23140
rect 12851 23072 13124 23100
rect 13556 23072 13676 23100
rect 13864 23100 13892 23140
rect 14369 23137 14381 23171
rect 14415 23137 14427 23171
rect 14369 23131 14427 23137
rect 14553 23171 14611 23177
rect 14553 23137 14565 23171
rect 14599 23137 14611 23171
rect 14553 23131 14611 23137
rect 14384 23100 14412 23131
rect 14826 23128 14832 23180
rect 14884 23128 14890 23180
rect 15381 23171 15439 23177
rect 15381 23137 15393 23171
rect 15427 23168 15439 23171
rect 15580 23168 15608 23196
rect 15427 23140 15608 23168
rect 15933 23171 15991 23177
rect 15427 23137 15439 23140
rect 15381 23131 15439 23137
rect 15933 23137 15945 23171
rect 15979 23137 15991 23171
rect 15933 23131 15991 23137
rect 14734 23100 14740 23112
rect 13864 23072 14740 23100
rect 12851 23069 12863 23072
rect 12805 23063 12863 23069
rect 1305 23035 1363 23041
rect 1305 23001 1317 23035
rect 1351 23032 1363 23035
rect 2133 23035 2191 23041
rect 1351 23004 1716 23032
rect 1351 23001 1363 23004
rect 1305 22995 1363 23001
rect 1688 22976 1716 23004
rect 2133 23001 2145 23035
rect 2179 23032 2191 23035
rect 2866 23032 2872 23044
rect 2179 23004 2872 23032
rect 2179 23001 2191 23004
rect 2133 22995 2191 23001
rect 2866 22992 2872 23004
rect 2924 22992 2930 23044
rect 7009 23035 7067 23041
rect 7009 23001 7021 23035
rect 7055 23032 7067 23035
rect 12529 23035 12587 23041
rect 7055 23004 9260 23032
rect 7055 23001 7067 23004
rect 7009 22995 7067 23001
rect 1670 22924 1676 22976
rect 1728 22964 1734 22976
rect 1949 22967 2007 22973
rect 1949 22964 1961 22967
rect 1728 22936 1961 22964
rect 1728 22924 1734 22936
rect 1949 22933 1961 22936
rect 1995 22933 2007 22967
rect 1949 22927 2007 22933
rect 3237 22967 3295 22973
rect 3237 22933 3249 22967
rect 3283 22964 3295 22967
rect 3786 22964 3792 22976
rect 3283 22936 3792 22964
rect 3283 22933 3295 22936
rect 3237 22927 3295 22933
rect 3786 22924 3792 22936
rect 3844 22924 3850 22976
rect 4522 22924 4528 22976
rect 4580 22924 4586 22976
rect 8938 22924 8944 22976
rect 8996 22964 9002 22976
rect 9125 22967 9183 22973
rect 9125 22964 9137 22967
rect 8996 22936 9137 22964
rect 8996 22924 9002 22936
rect 9125 22933 9137 22936
rect 9171 22933 9183 22967
rect 9232 22964 9260 23004
rect 12529 23001 12541 23035
rect 12575 23001 12587 23035
rect 12529 22995 12587 23001
rect 10042 22964 10048 22976
rect 9232 22936 10048 22964
rect 9125 22927 9183 22933
rect 10042 22924 10048 22936
rect 10100 22924 10106 22976
rect 10686 22924 10692 22976
rect 10744 22964 10750 22976
rect 10965 22967 11023 22973
rect 10965 22964 10977 22967
rect 10744 22936 10977 22964
rect 10744 22924 10750 22936
rect 10965 22933 10977 22936
rect 11011 22933 11023 22967
rect 10965 22927 11023 22933
rect 11606 22924 11612 22976
rect 11664 22964 11670 22976
rect 12544 22964 12572 22995
rect 12618 22992 12624 23044
rect 12676 22992 12682 23044
rect 13170 22992 13176 23044
rect 13228 22992 13234 23044
rect 11664 22936 12572 22964
rect 12897 22967 12955 22973
rect 11664 22924 11670 22936
rect 12897 22933 12909 22967
rect 12943 22964 12955 22967
rect 13556 22964 13584 23072
rect 14734 23060 14740 23072
rect 14792 23060 14798 23112
rect 13998 22992 14004 23044
rect 14056 23032 14062 23044
rect 14185 23035 14243 23041
rect 14185 23032 14197 23035
rect 14056 23004 14197 23032
rect 14056 22992 14062 23004
rect 14185 23001 14197 23004
rect 14231 23001 14243 23035
rect 15948 23032 15976 23131
rect 16758 23128 16764 23180
rect 16816 23128 16822 23180
rect 16850 23128 16856 23180
rect 16908 23168 16914 23180
rect 17144 23177 17172 23208
rect 18049 23205 18061 23239
rect 18095 23236 18107 23239
rect 18432 23236 18460 23267
rect 20990 23264 20996 23316
rect 21048 23304 21054 23316
rect 21545 23307 21603 23313
rect 21545 23304 21557 23307
rect 21048 23276 21557 23304
rect 21048 23264 21054 23276
rect 21545 23273 21557 23276
rect 21591 23273 21603 23307
rect 21545 23267 21603 23273
rect 21634 23264 21640 23316
rect 21692 23264 21698 23316
rect 19521 23239 19579 23245
rect 19521 23236 19533 23239
rect 18095 23208 18460 23236
rect 18570 23208 19533 23236
rect 18095 23205 18107 23208
rect 18049 23199 18107 23205
rect 17129 23171 17187 23177
rect 16908 23140 16953 23168
rect 16908 23128 16914 23140
rect 17129 23137 17141 23171
rect 17175 23137 17187 23171
rect 17129 23131 17187 23137
rect 17218 23128 17224 23180
rect 17276 23128 17282 23180
rect 17310 23128 17316 23180
rect 17368 23168 17374 23180
rect 17773 23171 17831 23177
rect 17773 23168 17785 23171
rect 17368 23140 17785 23168
rect 17368 23128 17374 23140
rect 17773 23137 17785 23140
rect 17819 23137 17831 23171
rect 17773 23131 17831 23137
rect 17865 23171 17923 23177
rect 17865 23137 17877 23171
rect 17911 23168 17923 23171
rect 18322 23168 18328 23180
rect 17911 23140 18328 23168
rect 17911 23137 17923 23140
rect 17865 23131 17923 23137
rect 18322 23128 18328 23140
rect 18380 23128 18386 23180
rect 18414 23128 18420 23180
rect 18472 23168 18478 23180
rect 18570 23177 18598 23208
rect 19521 23205 19533 23208
rect 19567 23205 19579 23239
rect 21910 23236 21916 23248
rect 19521 23199 19579 23205
rect 21468 23208 21916 23236
rect 18555 23171 18613 23177
rect 18555 23168 18567 23171
rect 18472 23140 18567 23168
rect 18472 23128 18478 23140
rect 18555 23137 18567 23140
rect 18601 23137 18613 23171
rect 18555 23131 18613 23137
rect 18690 23128 18696 23180
rect 18748 23128 18754 23180
rect 18782 23128 18788 23180
rect 18840 23128 18846 23180
rect 18874 23128 18880 23180
rect 18932 23177 18938 23180
rect 18932 23171 18971 23177
rect 18959 23137 18971 23171
rect 18932 23131 18971 23137
rect 18932 23128 18938 23131
rect 19058 23128 19064 23180
rect 19116 23128 19122 23180
rect 21468 23177 21496 23208
rect 21910 23196 21916 23208
rect 21968 23196 21974 23248
rect 19613 23171 19671 23177
rect 19613 23137 19625 23171
rect 19659 23168 19671 23171
rect 21453 23171 21511 23177
rect 21453 23168 21465 23171
rect 19659 23140 21465 23168
rect 19659 23137 19671 23140
rect 19613 23131 19671 23137
rect 21453 23137 21465 23140
rect 21499 23137 21511 23171
rect 21453 23131 21511 23137
rect 16577 23103 16635 23109
rect 16577 23069 16589 23103
rect 16623 23100 16635 23103
rect 18046 23100 18052 23112
rect 16623 23072 18052 23100
rect 16623 23069 16635 23072
rect 16577 23063 16635 23069
rect 18046 23060 18052 23072
rect 18104 23060 18110 23112
rect 17037 23035 17095 23041
rect 14185 22995 14243 23001
rect 15028 23004 16896 23032
rect 12943 22936 13584 22964
rect 12943 22933 12955 22936
rect 12897 22927 12955 22933
rect 13630 22924 13636 22976
rect 13688 22924 13694 22976
rect 13722 22924 13728 22976
rect 13780 22924 13786 22976
rect 14458 22924 14464 22976
rect 14516 22964 14522 22976
rect 14737 22967 14795 22973
rect 14737 22964 14749 22967
rect 14516 22936 14749 22964
rect 14516 22924 14522 22936
rect 14737 22933 14749 22936
rect 14783 22964 14795 22967
rect 15028 22964 15056 23004
rect 16868 22976 16896 23004
rect 17037 23001 17049 23035
rect 17083 23032 17095 23035
rect 21269 23035 21327 23041
rect 21269 23032 21281 23035
rect 17083 23004 19012 23032
rect 17083 23001 17095 23004
rect 17037 22995 17095 23001
rect 18984 22976 19012 23004
rect 19168 23004 21281 23032
rect 19168 22976 19196 23004
rect 21269 23001 21281 23004
rect 21315 23032 21327 23035
rect 21726 23032 21732 23044
rect 21315 23004 21732 23032
rect 21315 23001 21327 23004
rect 21269 22995 21327 23001
rect 21726 22992 21732 23004
rect 21784 22992 21790 23044
rect 14783 22936 15056 22964
rect 14783 22933 14795 22936
rect 14737 22927 14795 22933
rect 15102 22924 15108 22976
rect 15160 22924 15166 22976
rect 15838 22924 15844 22976
rect 15896 22924 15902 22976
rect 16850 22924 16856 22976
rect 16908 22924 16914 22976
rect 17586 22924 17592 22976
rect 17644 22924 17650 22976
rect 18049 22967 18107 22973
rect 18049 22933 18061 22967
rect 18095 22964 18107 22967
rect 18138 22964 18144 22976
rect 18095 22936 18144 22964
rect 18095 22933 18107 22936
rect 18049 22927 18107 22933
rect 18138 22924 18144 22936
rect 18196 22924 18202 22976
rect 18966 22924 18972 22976
rect 19024 22924 19030 22976
rect 19150 22924 19156 22976
rect 19208 22924 19214 22976
rect 21818 22924 21824 22976
rect 21876 22924 21882 22976
rect 552 22874 28428 22896
rect 552 22822 3882 22874
rect 3934 22822 3946 22874
rect 3998 22822 4010 22874
rect 4062 22822 4074 22874
rect 4126 22822 4138 22874
rect 4190 22822 10851 22874
rect 10903 22822 10915 22874
rect 10967 22822 10979 22874
rect 11031 22822 11043 22874
rect 11095 22822 11107 22874
rect 11159 22822 17820 22874
rect 17872 22822 17884 22874
rect 17936 22822 17948 22874
rect 18000 22822 18012 22874
rect 18064 22822 18076 22874
rect 18128 22822 24789 22874
rect 24841 22822 24853 22874
rect 24905 22822 24917 22874
rect 24969 22822 24981 22874
rect 25033 22822 25045 22874
rect 25097 22822 28428 22874
rect 552 22800 28428 22822
rect 1762 22720 1768 22772
rect 1820 22720 1826 22772
rect 2130 22720 2136 22772
rect 2188 22720 2194 22772
rect 3234 22720 3240 22772
rect 3292 22720 3298 22772
rect 3694 22720 3700 22772
rect 3752 22720 3758 22772
rect 3786 22720 3792 22772
rect 3844 22720 3850 22772
rect 4522 22720 4528 22772
rect 4580 22720 4586 22772
rect 5368 22732 5948 22760
rect 1780 22692 1808 22720
rect 2317 22695 2375 22701
rect 2317 22692 2329 22695
rect 1780 22664 2329 22692
rect 2317 22661 2329 22664
rect 2363 22661 2375 22695
rect 2317 22655 2375 22661
rect 3712 22624 3740 22720
rect 1780 22596 2452 22624
rect 1780 22565 1808 22596
rect 2424 22568 2452 22596
rect 2792 22596 3924 22624
rect 1765 22559 1823 22565
rect 1765 22525 1777 22559
rect 1811 22525 1823 22559
rect 1765 22519 1823 22525
rect 1949 22559 2007 22565
rect 1949 22525 1961 22559
rect 1995 22556 2007 22559
rect 2225 22559 2283 22565
rect 2225 22556 2237 22559
rect 1995 22528 2237 22556
rect 1995 22525 2007 22528
rect 1949 22519 2007 22525
rect 2225 22525 2237 22528
rect 2271 22525 2283 22559
rect 2225 22519 2283 22525
rect 2240 22488 2268 22519
rect 2406 22516 2412 22568
rect 2464 22556 2470 22568
rect 2792 22556 2820 22596
rect 2464 22528 2820 22556
rect 2464 22516 2470 22528
rect 3418 22516 3424 22568
rect 3476 22516 3482 22568
rect 3712 22565 3740 22596
rect 3896 22565 3924 22596
rect 3697 22559 3755 22565
rect 3697 22525 3709 22559
rect 3743 22525 3755 22559
rect 3697 22519 3755 22525
rect 3789 22559 3847 22565
rect 3789 22525 3801 22559
rect 3835 22525 3847 22559
rect 3789 22519 3847 22525
rect 3881 22559 3939 22565
rect 3881 22525 3893 22559
rect 3927 22525 3939 22559
rect 4540 22556 4568 22720
rect 5368 22701 5396 22732
rect 5353 22695 5411 22701
rect 5353 22661 5365 22695
rect 5399 22661 5411 22695
rect 5920 22692 5948 22732
rect 5994 22720 6000 22772
rect 6052 22760 6058 22772
rect 6178 22760 6184 22772
rect 6052 22732 6184 22760
rect 6052 22720 6058 22732
rect 6178 22720 6184 22732
rect 6236 22760 6242 22772
rect 6365 22763 6423 22769
rect 6365 22760 6377 22763
rect 6236 22732 6377 22760
rect 6236 22720 6242 22732
rect 6365 22729 6377 22732
rect 6411 22729 6423 22763
rect 6365 22723 6423 22729
rect 6914 22720 6920 22772
rect 6972 22760 6978 22772
rect 7929 22763 7987 22769
rect 7929 22760 7941 22763
rect 6972 22732 7941 22760
rect 6972 22720 6978 22732
rect 7929 22729 7941 22732
rect 7975 22729 7987 22763
rect 7929 22723 7987 22729
rect 8938 22720 8944 22772
rect 8996 22760 9002 22772
rect 9858 22760 9864 22772
rect 8996 22732 9864 22760
rect 8996 22720 9002 22732
rect 9858 22720 9864 22732
rect 9916 22760 9922 22772
rect 10410 22760 10416 22772
rect 9916 22732 10416 22760
rect 9916 22720 9922 22732
rect 10410 22720 10416 22732
rect 10468 22720 10474 22772
rect 11241 22763 11299 22769
rect 11241 22729 11253 22763
rect 11287 22760 11299 22763
rect 11422 22760 11428 22772
rect 11287 22732 11428 22760
rect 11287 22729 11299 22732
rect 11241 22723 11299 22729
rect 11422 22720 11428 22732
rect 11480 22720 11486 22772
rect 11790 22720 11796 22772
rect 11848 22720 11854 22772
rect 11882 22720 11888 22772
rect 11940 22720 11946 22772
rect 12158 22720 12164 22772
rect 12216 22720 12222 22772
rect 12529 22763 12587 22769
rect 12529 22729 12541 22763
rect 12575 22760 12587 22763
rect 12618 22760 12624 22772
rect 12575 22732 12624 22760
rect 12575 22729 12587 22732
rect 12529 22723 12587 22729
rect 12618 22720 12624 22732
rect 12676 22720 12682 22772
rect 12897 22763 12955 22769
rect 12897 22729 12909 22763
rect 12943 22760 12955 22763
rect 13817 22763 13875 22769
rect 12943 22732 13584 22760
rect 12943 22729 12955 22732
rect 12897 22723 12955 22729
rect 6546 22692 6552 22704
rect 5920 22664 6552 22692
rect 5353 22655 5411 22661
rect 6546 22652 6552 22664
rect 6604 22652 6610 22704
rect 6825 22695 6883 22701
rect 6825 22661 6837 22695
rect 6871 22692 6883 22695
rect 7745 22695 7803 22701
rect 7745 22692 7757 22695
rect 6871 22664 7757 22692
rect 6871 22661 6883 22664
rect 6825 22655 6883 22661
rect 7745 22661 7757 22664
rect 7791 22661 7803 22695
rect 11606 22692 11612 22704
rect 7745 22655 7803 22661
rect 8680 22664 11612 22692
rect 4709 22627 4767 22633
rect 4709 22593 4721 22627
rect 4755 22624 4767 22627
rect 5537 22627 5595 22633
rect 5537 22624 5549 22627
rect 4755 22596 5120 22624
rect 4755 22593 4767 22596
rect 4709 22587 4767 22593
rect 4801 22559 4859 22565
rect 4801 22556 4813 22559
rect 3881 22519 3939 22525
rect 3988 22528 4467 22556
rect 4540 22528 4813 22556
rect 3602 22488 3608 22500
rect 2240 22460 3608 22488
rect 3602 22448 3608 22460
rect 3660 22488 3666 22500
rect 3804 22488 3832 22519
rect 3988 22488 4016 22528
rect 3660 22460 4016 22488
rect 4065 22491 4123 22497
rect 3660 22448 3666 22460
rect 4065 22457 4077 22491
rect 4111 22457 4123 22491
rect 4065 22451 4123 22457
rect 3418 22380 3424 22432
rect 3476 22420 3482 22432
rect 4080 22420 4108 22451
rect 4338 22448 4344 22500
rect 4396 22448 4402 22500
rect 4439 22488 4467 22528
rect 4801 22525 4813 22528
rect 4847 22525 4859 22559
rect 4801 22519 4859 22525
rect 4890 22516 4896 22568
rect 4948 22556 4954 22568
rect 5092 22565 5120 22596
rect 5276 22596 5549 22624
rect 4985 22559 5043 22565
rect 4985 22556 4997 22559
rect 4948 22528 4997 22556
rect 4948 22516 4954 22528
rect 4985 22525 4997 22528
rect 5031 22525 5043 22559
rect 4985 22519 5043 22525
rect 5077 22559 5135 22565
rect 5077 22525 5089 22559
rect 5123 22525 5135 22559
rect 5077 22519 5135 22525
rect 5169 22559 5227 22565
rect 5169 22525 5181 22559
rect 5215 22558 5227 22559
rect 5276 22558 5304 22596
rect 5537 22593 5549 22596
rect 5583 22593 5595 22627
rect 6362 22624 6368 22636
rect 5537 22587 5595 22593
rect 5644 22596 6368 22624
rect 5215 22530 5304 22558
rect 5215 22525 5227 22530
rect 5169 22519 5227 22525
rect 5350 22516 5356 22568
rect 5408 22556 5414 22568
rect 5644 22565 5672 22596
rect 6362 22584 6368 22596
rect 6420 22584 6426 22636
rect 6454 22584 6460 22636
rect 6512 22584 6518 22636
rect 7760 22624 7788 22655
rect 8680 22633 8708 22664
rect 11606 22652 11612 22664
rect 11664 22652 11670 22704
rect 8665 22627 8723 22633
rect 7760 22596 8616 22624
rect 5445 22559 5503 22565
rect 5445 22556 5457 22559
rect 5408 22528 5457 22556
rect 5408 22516 5414 22528
rect 5445 22525 5457 22528
rect 5491 22525 5503 22559
rect 5445 22519 5503 22525
rect 5629 22559 5687 22565
rect 5629 22525 5641 22559
rect 5675 22525 5687 22559
rect 5629 22519 5687 22525
rect 5813 22559 5871 22565
rect 5813 22525 5825 22559
rect 5859 22525 5871 22559
rect 5813 22519 5871 22525
rect 6181 22559 6239 22565
rect 6181 22525 6193 22559
rect 6227 22556 6239 22559
rect 6380 22556 6408 22584
rect 6641 22559 6699 22565
rect 6641 22556 6653 22559
rect 6227 22528 6653 22556
rect 6227 22525 6239 22528
rect 6181 22519 6239 22525
rect 6641 22525 6653 22528
rect 6687 22525 6699 22559
rect 6641 22519 6699 22525
rect 7653 22559 7711 22565
rect 7653 22525 7665 22559
rect 7699 22556 7711 22559
rect 8018 22556 8024 22568
rect 7699 22528 8024 22556
rect 7699 22525 7711 22528
rect 7653 22519 7711 22525
rect 4525 22491 4583 22497
rect 4525 22488 4537 22491
rect 4439 22460 4537 22488
rect 4525 22457 4537 22460
rect 4571 22488 4583 22491
rect 5644 22488 5672 22519
rect 4571 22460 5672 22488
rect 5828 22488 5856 22519
rect 8018 22516 8024 22528
rect 8076 22516 8082 22568
rect 8588 22565 8616 22596
rect 8665 22593 8677 22627
rect 8711 22593 8723 22627
rect 8665 22587 8723 22593
rect 8754 22584 8760 22636
rect 8812 22584 8818 22636
rect 11808 22624 11836 22720
rect 11164 22596 11836 22624
rect 11900 22692 11928 22720
rect 12912 22692 12940 22723
rect 11900 22664 12940 22692
rect 8481 22559 8539 22565
rect 8481 22558 8493 22559
rect 8404 22530 8493 22558
rect 6365 22491 6423 22497
rect 6365 22488 6377 22491
rect 5828 22460 6377 22488
rect 4571 22457 4583 22460
rect 4525 22451 4583 22457
rect 6365 22457 6377 22460
rect 6411 22488 6423 22491
rect 6730 22488 6736 22500
rect 6411 22460 6736 22488
rect 6411 22457 6423 22460
rect 6365 22451 6423 22457
rect 6730 22448 6736 22460
rect 6788 22448 6794 22500
rect 7561 22491 7619 22497
rect 7561 22457 7573 22491
rect 7607 22488 7619 22491
rect 7742 22488 7748 22500
rect 7607 22460 7748 22488
rect 7607 22457 7619 22460
rect 7561 22451 7619 22457
rect 7742 22448 7748 22460
rect 7800 22448 7806 22500
rect 7929 22491 7987 22497
rect 7929 22457 7941 22491
rect 7975 22488 7987 22491
rect 8294 22488 8300 22500
rect 7975 22460 8300 22488
rect 7975 22457 7987 22460
rect 7929 22451 7987 22457
rect 8294 22448 8300 22460
rect 8352 22448 8358 22500
rect 8404 22488 8432 22530
rect 8481 22525 8493 22530
rect 8527 22525 8539 22559
rect 8481 22519 8539 22525
rect 8573 22559 8631 22565
rect 8573 22525 8585 22559
rect 8619 22525 8631 22559
rect 9674 22556 9680 22568
rect 8956 22534 9680 22556
rect 8573 22519 8631 22525
rect 8680 22528 9680 22534
rect 8680 22506 8984 22528
rect 9674 22516 9680 22528
rect 9732 22516 9738 22568
rect 10686 22516 10692 22568
rect 10744 22556 10750 22568
rect 11164 22565 11192 22596
rect 10965 22559 11023 22565
rect 10965 22556 10977 22559
rect 10744 22528 10977 22556
rect 10744 22516 10750 22528
rect 10965 22525 10977 22528
rect 11011 22525 11023 22559
rect 10965 22519 11023 22525
rect 11149 22559 11207 22565
rect 11149 22525 11161 22559
rect 11195 22525 11207 22559
rect 11149 22519 11207 22525
rect 11241 22559 11299 22565
rect 11241 22525 11253 22559
rect 11287 22525 11299 22559
rect 11241 22519 11299 22525
rect 11793 22559 11851 22565
rect 11793 22525 11805 22559
rect 11839 22556 11851 22559
rect 11900 22556 11928 22664
rect 12710 22584 12716 22636
rect 12768 22624 12774 22636
rect 13556 22624 13584 22732
rect 13817 22729 13829 22763
rect 13863 22760 13875 22763
rect 13863 22732 14320 22760
rect 13863 22729 13875 22732
rect 13817 22723 13875 22729
rect 13630 22652 13636 22704
rect 13688 22692 13694 22704
rect 13909 22695 13967 22701
rect 13909 22692 13921 22695
rect 13688 22664 13921 22692
rect 13688 22652 13694 22664
rect 13909 22661 13921 22664
rect 13955 22661 13967 22695
rect 13909 22655 13967 22661
rect 13998 22652 14004 22704
rect 14056 22652 14062 22704
rect 14292 22692 14320 22732
rect 16390 22720 16396 22772
rect 16448 22720 16454 22772
rect 18693 22763 18751 22769
rect 18693 22729 18705 22763
rect 18739 22760 18751 22763
rect 19058 22760 19064 22772
rect 18739 22732 19064 22760
rect 18739 22729 18751 22732
rect 18693 22723 18751 22729
rect 19058 22720 19064 22732
rect 19116 22720 19122 22772
rect 20165 22763 20223 22769
rect 20165 22760 20177 22763
rect 19168 22732 20177 22760
rect 15286 22692 15292 22704
rect 14292 22664 15292 22692
rect 15286 22652 15292 22664
rect 15344 22652 15350 22704
rect 16209 22695 16267 22701
rect 16209 22692 16221 22695
rect 15580 22664 16221 22692
rect 12768 22596 12940 22624
rect 13556 22596 13860 22624
rect 12768 22584 12774 22596
rect 11839 22528 11928 22556
rect 11977 22559 12035 22565
rect 11839 22525 11851 22528
rect 11793 22519 11851 22525
rect 11977 22525 11989 22559
rect 12023 22556 12035 22559
rect 12802 22556 12808 22568
rect 12023 22528 12808 22556
rect 12023 22525 12035 22528
rect 11977 22519 12035 22525
rect 8680 22488 8708 22506
rect 8404 22460 8708 22488
rect 4614 22420 4620 22432
rect 3476 22392 4620 22420
rect 3476 22380 3482 22392
rect 4614 22380 4620 22392
rect 4672 22420 4678 22432
rect 5810 22420 5816 22432
rect 4672 22392 5816 22420
rect 4672 22380 4678 22392
rect 5810 22380 5816 22392
rect 5868 22420 5874 22432
rect 5905 22423 5963 22429
rect 5905 22420 5917 22423
rect 5868 22392 5917 22420
rect 5868 22380 5874 22392
rect 5905 22389 5917 22392
rect 5951 22389 5963 22423
rect 5905 22383 5963 22389
rect 5994 22380 6000 22432
rect 6052 22380 6058 22432
rect 6181 22423 6239 22429
rect 6181 22389 6193 22423
rect 6227 22420 6239 22423
rect 8754 22420 8760 22432
rect 6227 22392 8760 22420
rect 6227 22389 6239 22392
rect 6181 22383 6239 22389
rect 8754 22380 8760 22392
rect 8812 22380 8818 22432
rect 8938 22380 8944 22432
rect 8996 22380 9002 22432
rect 11256 22420 11284 22519
rect 12802 22516 12808 22528
rect 12860 22516 12866 22568
rect 12912 22565 12940 22596
rect 12897 22559 12955 22565
rect 12897 22525 12909 22559
rect 12943 22525 12955 22559
rect 12897 22519 12955 22525
rect 11698 22448 11704 22500
rect 11756 22488 11762 22500
rect 11756 22460 12653 22488
rect 11756 22448 11762 22460
rect 12526 22420 12532 22432
rect 11256 22392 12532 22420
rect 12526 22380 12532 22392
rect 12584 22380 12590 22432
rect 12625 22420 12653 22460
rect 13354 22448 13360 22500
rect 13412 22488 13418 22500
rect 13725 22491 13783 22497
rect 13725 22488 13737 22491
rect 13412 22460 13737 22488
rect 13412 22448 13418 22460
rect 13725 22457 13737 22460
rect 13771 22457 13783 22491
rect 13832 22488 13860 22596
rect 14016 22565 14044 22652
rect 15580 22633 15608 22664
rect 16209 22661 16221 22664
rect 16255 22661 16267 22695
rect 16209 22655 16267 22661
rect 18966 22652 18972 22704
rect 19024 22692 19030 22704
rect 19168 22692 19196 22732
rect 20165 22729 20177 22732
rect 20211 22760 20223 22763
rect 20806 22760 20812 22772
rect 20211 22732 20812 22760
rect 20211 22729 20223 22732
rect 20165 22723 20223 22729
rect 20806 22720 20812 22732
rect 20864 22720 20870 22772
rect 22370 22720 22376 22772
rect 22428 22720 22434 22772
rect 19024 22664 19196 22692
rect 19024 22652 19030 22664
rect 19334 22652 19340 22704
rect 19392 22692 19398 22704
rect 20073 22695 20131 22701
rect 20073 22692 20085 22695
rect 19392 22664 20085 22692
rect 19392 22652 19398 22664
rect 20073 22661 20085 22664
rect 20119 22661 20131 22695
rect 20073 22655 20131 22661
rect 20254 22652 20260 22704
rect 20312 22652 20318 22704
rect 20714 22692 20720 22704
rect 20364 22664 20720 22692
rect 15565 22627 15623 22633
rect 15565 22593 15577 22627
rect 15611 22593 15623 22627
rect 15565 22587 15623 22593
rect 15838 22584 15844 22636
rect 15896 22584 15902 22636
rect 18230 22584 18236 22636
rect 18288 22624 18294 22636
rect 18288 22596 19104 22624
rect 18288 22584 18294 22596
rect 19076 22568 19104 22596
rect 19150 22584 19156 22636
rect 19208 22584 19214 22636
rect 20364 22624 20392 22664
rect 20714 22652 20720 22664
rect 20772 22652 20778 22704
rect 21174 22652 21180 22704
rect 21232 22692 21238 22704
rect 22388 22692 22416 22720
rect 21232 22664 22508 22692
rect 21232 22652 21238 22664
rect 20272 22596 20392 22624
rect 20625 22627 20683 22633
rect 14001 22559 14059 22565
rect 14001 22525 14013 22559
rect 14047 22525 14059 22559
rect 14001 22519 14059 22525
rect 14093 22559 14151 22565
rect 14093 22525 14105 22559
rect 14139 22556 14151 22559
rect 14182 22556 14188 22568
rect 14139 22528 14188 22556
rect 14139 22525 14151 22528
rect 14093 22519 14151 22525
rect 14182 22516 14188 22528
rect 14240 22556 14246 22568
rect 14826 22556 14832 22568
rect 14240 22528 14832 22556
rect 14240 22516 14246 22528
rect 14826 22516 14832 22528
rect 14884 22516 14890 22568
rect 15473 22559 15531 22565
rect 15473 22525 15485 22559
rect 15519 22525 15531 22559
rect 15473 22519 15531 22525
rect 14458 22488 14464 22500
rect 13832 22460 14464 22488
rect 13725 22451 13783 22457
rect 14458 22448 14464 22460
rect 14516 22448 14522 22500
rect 12894 22420 12900 22432
rect 12625 22392 12900 22420
rect 12894 22380 12900 22392
rect 12952 22420 12958 22432
rect 14277 22423 14335 22429
rect 14277 22420 14289 22423
rect 12952 22392 14289 22420
rect 12952 22380 12958 22392
rect 14277 22389 14289 22392
rect 14323 22420 14335 22423
rect 15488 22420 15516 22519
rect 19058 22516 19064 22568
rect 19116 22516 19122 22568
rect 19957 22559 20015 22565
rect 19957 22556 19969 22559
rect 19306 22528 19969 22556
rect 16577 22491 16635 22497
rect 16577 22457 16589 22491
rect 16623 22488 16635 22491
rect 18138 22488 18144 22500
rect 16623 22460 18144 22488
rect 16623 22457 16635 22460
rect 16577 22451 16635 22457
rect 18138 22448 18144 22460
rect 18196 22488 18202 22500
rect 19306 22488 19334 22528
rect 19957 22525 19969 22528
rect 20003 22556 20015 22559
rect 20272 22558 20300 22596
rect 20625 22593 20637 22627
rect 20671 22624 20683 22627
rect 22186 22624 22192 22636
rect 20671 22596 22192 22624
rect 20671 22593 20683 22596
rect 20625 22587 20683 22593
rect 20374 22559 20432 22565
rect 20374 22558 20386 22559
rect 20003 22528 20208 22556
rect 20272 22530 20386 22558
rect 20364 22528 20386 22530
rect 20003 22525 20015 22528
rect 19957 22519 20015 22525
rect 18196 22460 19334 22488
rect 18196 22448 18202 22460
rect 14323 22392 15516 22420
rect 16377 22423 16435 22429
rect 14323 22389 14335 22392
rect 14277 22383 14335 22389
rect 16377 22389 16389 22423
rect 16423 22420 16435 22423
rect 16482 22420 16488 22432
rect 16423 22392 16488 22420
rect 16423 22389 16435 22392
rect 16377 22383 16435 22389
rect 16482 22380 16488 22392
rect 16540 22380 16546 22432
rect 20180 22420 20208 22528
rect 20374 22525 20386 22528
rect 20420 22525 20432 22559
rect 20374 22519 20432 22525
rect 20530 22516 20536 22568
rect 20588 22556 20594 22568
rect 20588 22528 20944 22556
rect 20588 22516 20594 22528
rect 20254 22448 20260 22500
rect 20312 22488 20318 22500
rect 20717 22491 20775 22497
rect 20717 22488 20729 22491
rect 20312 22460 20729 22488
rect 20312 22448 20318 22460
rect 20717 22457 20729 22460
rect 20763 22457 20775 22491
rect 20916 22488 20944 22528
rect 20990 22516 20996 22568
rect 21048 22516 21054 22568
rect 21560 22565 21588 22596
rect 22186 22584 22192 22596
rect 22244 22624 22250 22636
rect 22480 22633 22508 22664
rect 22373 22627 22431 22633
rect 22373 22624 22385 22627
rect 22244 22596 22385 22624
rect 22244 22584 22250 22596
rect 22373 22593 22385 22596
rect 22419 22593 22431 22627
rect 22373 22587 22431 22593
rect 22465 22627 22523 22633
rect 22465 22593 22477 22627
rect 22511 22624 22523 22627
rect 22646 22624 22652 22636
rect 22511 22596 22652 22624
rect 22511 22593 22523 22596
rect 22465 22587 22523 22593
rect 22646 22584 22652 22596
rect 22704 22584 22710 22636
rect 23290 22584 23296 22636
rect 23348 22584 23354 22636
rect 23842 22584 23848 22636
rect 23900 22584 23906 22636
rect 21361 22559 21419 22565
rect 21361 22525 21373 22559
rect 21407 22525 21419 22559
rect 21361 22519 21419 22525
rect 21545 22559 21603 22565
rect 21545 22525 21557 22559
rect 21591 22525 21603 22559
rect 21545 22519 21603 22525
rect 22281 22559 22339 22565
rect 22281 22525 22293 22559
rect 22327 22525 22339 22559
rect 22281 22519 22339 22525
rect 21376 22488 21404 22519
rect 20916 22460 21404 22488
rect 20717 22451 20775 22457
rect 22296 22432 22324 22519
rect 22554 22516 22560 22568
rect 22612 22516 22618 22568
rect 23474 22516 23480 22568
rect 23532 22516 23538 22568
rect 23106 22448 23112 22500
rect 23164 22448 23170 22500
rect 24112 22491 24170 22497
rect 24112 22457 24124 22491
rect 24158 22488 24170 22491
rect 24302 22488 24308 22500
rect 24158 22460 24308 22488
rect 24158 22457 24170 22460
rect 24112 22451 24170 22457
rect 24302 22448 24308 22460
rect 24360 22448 24366 22500
rect 20530 22420 20536 22432
rect 20180 22392 20536 22420
rect 20530 22380 20536 22392
rect 20588 22420 20594 22432
rect 20809 22423 20867 22429
rect 20809 22420 20821 22423
rect 20588 22392 20821 22420
rect 20588 22380 20594 22392
rect 20809 22389 20821 22392
rect 20855 22389 20867 22423
rect 20809 22383 20867 22389
rect 21453 22423 21511 22429
rect 21453 22389 21465 22423
rect 21499 22420 21511 22423
rect 21634 22420 21640 22432
rect 21499 22392 21640 22420
rect 21499 22389 21511 22392
rect 21453 22383 21511 22389
rect 21634 22380 21640 22392
rect 21692 22380 21698 22432
rect 22094 22380 22100 22432
rect 22152 22380 22158 22432
rect 22278 22380 22284 22432
rect 22336 22420 22342 22432
rect 23124 22420 23152 22448
rect 22336 22392 23152 22420
rect 22336 22380 22342 22392
rect 23658 22380 23664 22432
rect 23716 22380 23722 22432
rect 25222 22380 25228 22432
rect 25280 22380 25286 22432
rect 552 22330 28587 22352
rect 552 22278 7366 22330
rect 7418 22278 7430 22330
rect 7482 22278 7494 22330
rect 7546 22278 7558 22330
rect 7610 22278 7622 22330
rect 7674 22278 14335 22330
rect 14387 22278 14399 22330
rect 14451 22278 14463 22330
rect 14515 22278 14527 22330
rect 14579 22278 14591 22330
rect 14643 22278 21304 22330
rect 21356 22278 21368 22330
rect 21420 22278 21432 22330
rect 21484 22278 21496 22330
rect 21548 22278 21560 22330
rect 21612 22278 28273 22330
rect 28325 22278 28337 22330
rect 28389 22278 28401 22330
rect 28453 22278 28465 22330
rect 28517 22278 28529 22330
rect 28581 22278 28587 22330
rect 552 22256 28587 22278
rect 4801 22219 4859 22225
rect 4801 22185 4813 22219
rect 4847 22216 4859 22219
rect 4890 22216 4896 22228
rect 4847 22188 4896 22216
rect 4847 22185 4859 22188
rect 4801 22179 4859 22185
rect 4890 22176 4896 22188
rect 4948 22176 4954 22228
rect 5810 22176 5816 22228
rect 5868 22216 5874 22228
rect 6454 22216 6460 22228
rect 5868 22188 6460 22216
rect 5868 22176 5874 22188
rect 6454 22176 6460 22188
rect 6512 22176 6518 22228
rect 8938 22176 8944 22228
rect 8996 22176 9002 22228
rect 9600 22188 10824 22216
rect 4430 22108 4436 22160
rect 4488 22148 4494 22160
rect 5350 22148 5356 22160
rect 4488 22120 5356 22148
rect 4488 22108 4494 22120
rect 5350 22108 5356 22120
rect 5408 22108 5414 22160
rect 1486 22040 1492 22092
rect 1544 22040 1550 22092
rect 1581 22083 1639 22089
rect 1581 22049 1593 22083
rect 1627 22049 1639 22083
rect 1581 22043 1639 22049
rect 1765 22083 1823 22089
rect 1765 22049 1777 22083
rect 1811 22080 1823 22083
rect 1854 22080 1860 22092
rect 1811 22052 1860 22080
rect 1811 22049 1823 22052
rect 1765 22043 1823 22049
rect 1596 22012 1624 22043
rect 1854 22040 1860 22052
rect 1912 22040 1918 22092
rect 4617 22083 4675 22089
rect 4617 22049 4629 22083
rect 4663 22049 4675 22083
rect 4617 22043 4675 22049
rect 2593 22015 2651 22021
rect 2593 22012 2605 22015
rect 1596 21984 2084 22012
rect 2056 21888 2084 21984
rect 2424 21984 2605 22012
rect 2424 21888 2452 21984
rect 2593 21981 2605 21984
rect 2639 22012 2651 22015
rect 2639 21984 2774 22012
rect 2639 21981 2651 21984
rect 2593 21975 2651 21981
rect 2746 21944 2774 21984
rect 3418 21972 3424 22024
rect 3476 22012 3482 22024
rect 4632 22012 4660 22043
rect 6730 22040 6736 22092
rect 6788 22080 6794 22092
rect 7101 22083 7159 22089
rect 7101 22080 7113 22083
rect 6788 22052 7113 22080
rect 6788 22040 6794 22052
rect 7101 22049 7113 22052
rect 7147 22049 7159 22083
rect 7101 22043 7159 22049
rect 8478 22040 8484 22092
rect 8536 22040 8542 22092
rect 8665 22083 8723 22089
rect 8665 22049 8677 22083
rect 8711 22049 8723 22083
rect 8956 22080 8984 22176
rect 9600 22092 9628 22188
rect 9674 22108 9680 22160
rect 9732 22148 9738 22160
rect 10594 22148 10600 22160
rect 9732 22120 10600 22148
rect 9732 22108 9738 22120
rect 10594 22108 10600 22120
rect 10652 22108 10658 22160
rect 10796 22157 10824 22188
rect 13004 22188 13584 22216
rect 10781 22151 10839 22157
rect 10781 22117 10793 22151
rect 10827 22148 10839 22151
rect 10827 22120 11376 22148
rect 10827 22117 10839 22120
rect 10781 22111 10839 22117
rect 9309 22083 9367 22089
rect 9309 22080 9321 22083
rect 8956 22052 9321 22080
rect 8665 22043 8723 22049
rect 9309 22049 9321 22052
rect 9355 22049 9367 22083
rect 9309 22043 9367 22049
rect 9401 22083 9459 22089
rect 9401 22049 9413 22083
rect 9447 22049 9459 22083
rect 9582 22080 9588 22092
rect 9543 22052 9588 22080
rect 9401 22043 9459 22049
rect 3476 21984 4660 22012
rect 8680 22012 8708 22043
rect 9416 22012 9444 22043
rect 9582 22040 9588 22052
rect 9640 22040 9646 22092
rect 10502 22040 10508 22092
rect 10560 22080 10566 22092
rect 10965 22083 11023 22089
rect 10965 22080 10977 22083
rect 10560 22052 10977 22080
rect 10560 22040 10566 22052
rect 10965 22049 10977 22052
rect 11011 22049 11023 22083
rect 10965 22043 11023 22049
rect 11054 22040 11060 22092
rect 11112 22080 11118 22092
rect 11348 22089 11376 22120
rect 12250 22108 12256 22160
rect 12308 22148 12314 22160
rect 13004 22148 13032 22188
rect 12308 22120 13032 22148
rect 12308 22108 12314 22120
rect 13354 22108 13360 22160
rect 13412 22108 13418 22160
rect 13556 22157 13584 22188
rect 17328 22188 19334 22216
rect 13541 22151 13599 22157
rect 13541 22117 13553 22151
rect 13587 22117 13599 22151
rect 13541 22111 13599 22117
rect 13630 22108 13636 22160
rect 13688 22148 13694 22160
rect 13725 22151 13783 22157
rect 13725 22148 13737 22151
rect 13688 22120 13737 22148
rect 13688 22108 13694 22120
rect 13725 22117 13737 22120
rect 13771 22117 13783 22151
rect 13725 22111 13783 22117
rect 16114 22108 16120 22160
rect 16172 22148 16178 22160
rect 17218 22148 17224 22160
rect 16172 22120 17224 22148
rect 16172 22108 16178 22120
rect 17218 22108 17224 22120
rect 17276 22108 17282 22160
rect 11149 22083 11207 22089
rect 11149 22080 11161 22083
rect 11112 22052 11161 22080
rect 11112 22040 11118 22052
rect 11149 22049 11161 22052
rect 11195 22049 11207 22083
rect 11149 22043 11207 22049
rect 11241 22083 11299 22089
rect 11241 22049 11253 22083
rect 11287 22049 11299 22083
rect 11241 22043 11299 22049
rect 11333 22083 11391 22089
rect 11333 22049 11345 22083
rect 11379 22080 11391 22083
rect 11379 22052 11413 22080
rect 11379 22049 11391 22052
rect 11333 22043 11391 22049
rect 11256 22012 11284 22043
rect 14734 22040 14740 22092
rect 14792 22080 14798 22092
rect 16393 22083 16451 22089
rect 16393 22080 16405 22083
rect 14792 22052 16405 22080
rect 14792 22040 14798 22052
rect 16393 22049 16405 22052
rect 16439 22049 16451 22083
rect 16393 22043 16451 22049
rect 8680 21984 9076 22012
rect 3476 21972 3482 21984
rect 6454 21944 6460 21956
rect 2746 21916 6460 21944
rect 6454 21904 6460 21916
rect 6512 21944 6518 21956
rect 6512 21916 8524 21944
rect 6512 21904 6518 21916
rect 1762 21836 1768 21888
rect 1820 21836 1826 21888
rect 2038 21836 2044 21888
rect 2096 21836 2102 21888
rect 2406 21836 2412 21888
rect 2464 21836 2470 21888
rect 6638 21836 6644 21888
rect 6696 21876 6702 21888
rect 6917 21879 6975 21885
rect 6917 21876 6929 21879
rect 6696 21848 6929 21876
rect 6696 21836 6702 21848
rect 6917 21845 6929 21848
rect 6963 21845 6975 21879
rect 6917 21839 6975 21845
rect 8294 21836 8300 21888
rect 8352 21836 8358 21888
rect 8496 21885 8524 21916
rect 9048 21888 9076 21984
rect 9324 21984 11284 22012
rect 11609 22015 11667 22021
rect 9324 21888 9352 21984
rect 11609 21981 11621 22015
rect 11655 22012 11667 22015
rect 12434 22012 12440 22024
rect 11655 21984 12440 22012
rect 11655 21981 11667 21984
rect 11609 21975 11667 21981
rect 12434 21972 12440 21984
rect 12492 21972 12498 22024
rect 12618 21972 12624 22024
rect 12676 22012 12682 22024
rect 15102 22012 15108 22024
rect 12676 21984 15108 22012
rect 12676 21972 12682 21984
rect 15102 21972 15108 21984
rect 15160 21972 15166 22024
rect 16482 21972 16488 22024
rect 16540 21972 16546 22024
rect 9585 21947 9643 21953
rect 9585 21913 9597 21947
rect 9631 21944 9643 21947
rect 9950 21944 9956 21956
rect 9631 21916 9956 21944
rect 9631 21913 9643 21916
rect 9585 21907 9643 21913
rect 9950 21904 9956 21916
rect 10008 21904 10014 21956
rect 10781 21947 10839 21953
rect 10781 21913 10793 21947
rect 10827 21944 10839 21947
rect 11146 21944 11152 21956
rect 10827 21916 11152 21944
rect 10827 21913 10839 21916
rect 10781 21907 10839 21913
rect 11146 21904 11152 21916
rect 11204 21904 11210 21956
rect 11974 21904 11980 21956
rect 12032 21944 12038 21956
rect 17328 21944 17356 22188
rect 18874 22108 18880 22160
rect 18932 22148 18938 22160
rect 19030 22151 19088 22157
rect 19030 22148 19042 22151
rect 18932 22120 19042 22148
rect 18932 22108 18938 22120
rect 19030 22117 19042 22120
rect 19076 22117 19088 22151
rect 19030 22111 19088 22117
rect 19306 22080 19334 22188
rect 19702 22176 19708 22228
rect 19760 22176 19766 22228
rect 20990 22216 20996 22228
rect 20640 22188 20996 22216
rect 19720 22148 19748 22176
rect 20640 22157 20668 22188
rect 20990 22176 20996 22188
rect 21048 22176 21054 22228
rect 22554 22176 22560 22228
rect 22612 22216 22618 22228
rect 22612 22188 22784 22216
rect 22612 22176 22618 22188
rect 20625 22151 20683 22157
rect 20625 22148 20637 22151
rect 19720 22120 20637 22148
rect 20625 22117 20637 22120
rect 20671 22117 20683 22151
rect 20625 22111 20683 22117
rect 21726 22108 21732 22160
rect 21784 22108 21790 22160
rect 22094 22148 22100 22160
rect 21928 22120 22100 22148
rect 19426 22080 19432 22092
rect 19306 22052 19432 22080
rect 19426 22040 19432 22052
rect 19484 22080 19490 22092
rect 19484 22052 20208 22080
rect 19484 22040 19490 22052
rect 18782 21972 18788 22024
rect 18840 21972 18846 22024
rect 20180 22012 20208 22052
rect 20254 22040 20260 22092
rect 20312 22080 20318 22092
rect 20349 22083 20407 22089
rect 20349 22080 20361 22083
rect 20312 22052 20361 22080
rect 20312 22040 20318 22052
rect 20349 22049 20361 22052
rect 20395 22049 20407 22083
rect 20349 22043 20407 22049
rect 20441 22083 20499 22089
rect 20441 22049 20453 22083
rect 20487 22080 20499 22083
rect 20530 22080 20536 22092
rect 20487 22052 20536 22080
rect 20487 22049 20499 22052
rect 20441 22043 20499 22049
rect 20530 22040 20536 22052
rect 20588 22040 20594 22092
rect 21637 22083 21695 22089
rect 21637 22049 21649 22083
rect 21683 22080 21695 22083
rect 21928 22080 21956 22120
rect 22094 22108 22100 22120
rect 22152 22108 22158 22160
rect 22278 22108 22284 22160
rect 22336 22148 22342 22160
rect 22336 22120 22508 22148
rect 22336 22108 22342 22120
rect 21683 22052 21956 22080
rect 22005 22083 22063 22089
rect 21683 22049 21695 22052
rect 21637 22043 21695 22049
rect 22005 22049 22017 22083
rect 22051 22080 22063 22083
rect 22373 22083 22431 22089
rect 22373 22080 22385 22083
rect 22051 22052 22385 22080
rect 22051 22049 22063 22052
rect 22005 22043 22063 22049
rect 22373 22049 22385 22052
rect 22419 22049 22431 22083
rect 22480 22080 22508 22120
rect 22756 22094 22784 22188
rect 23658 22176 23664 22228
rect 23716 22176 23722 22228
rect 24302 22176 24308 22228
rect 24360 22176 24366 22228
rect 22940 22120 23428 22148
rect 22557 22083 22615 22089
rect 22557 22080 22569 22083
rect 22480 22052 22569 22080
rect 22373 22043 22431 22049
rect 22557 22049 22569 22052
rect 22603 22049 22615 22083
rect 22557 22043 22615 22049
rect 22646 22040 22652 22092
rect 22704 22040 22710 22092
rect 22756 22089 22876 22094
rect 22940 22092 22968 22120
rect 22756 22083 22891 22089
rect 22756 22066 22845 22083
rect 22833 22049 22845 22066
rect 22879 22049 22891 22083
rect 22833 22043 22891 22049
rect 22922 22040 22928 22092
rect 22980 22040 22986 22092
rect 23400 22089 23428 22120
rect 23109 22083 23167 22089
rect 23109 22049 23121 22083
rect 23155 22049 23167 22083
rect 23109 22043 23167 22049
rect 23293 22083 23351 22089
rect 23293 22049 23305 22083
rect 23339 22049 23351 22083
rect 23293 22043 23351 22049
rect 23381 22083 23439 22089
rect 23381 22049 23393 22083
rect 23427 22049 23439 22083
rect 23381 22043 23439 22049
rect 20990 22012 20996 22024
rect 20180 21984 20996 22012
rect 20990 21972 20996 21984
rect 21048 21972 21054 22024
rect 22097 22015 22155 22021
rect 22097 21981 22109 22015
rect 22143 21981 22155 22015
rect 22097 21975 22155 21981
rect 12032 21916 17356 21944
rect 12032 21904 12038 21916
rect 20346 21904 20352 21956
rect 20404 21944 20410 21956
rect 20625 21947 20683 21953
rect 20625 21944 20637 21947
rect 20404 21916 20637 21944
rect 20404 21904 20410 21916
rect 20625 21913 20637 21916
rect 20671 21913 20683 21947
rect 20625 21907 20683 21913
rect 21634 21904 21640 21956
rect 21692 21944 21698 21956
rect 22112 21944 22140 21975
rect 22462 21972 22468 22024
rect 22520 22012 22526 22024
rect 23124 22012 23152 22043
rect 22520 21984 23152 22012
rect 22520 21972 22526 21984
rect 21692 21916 22140 21944
rect 22281 21947 22339 21953
rect 21692 21904 21698 21916
rect 22281 21913 22293 21947
rect 22327 21944 22339 21947
rect 23308 21944 23336 22043
rect 23474 22040 23480 22092
rect 23532 22040 23538 22092
rect 23676 22080 23704 22176
rect 24489 22083 24547 22089
rect 24489 22080 24501 22083
rect 23676 22052 24501 22080
rect 24489 22049 24501 22052
rect 24535 22049 24547 22083
rect 24489 22043 24547 22049
rect 22327 21916 23336 21944
rect 22327 21913 22339 21916
rect 22281 21907 22339 21913
rect 23566 21904 23572 21956
rect 23624 21944 23630 21956
rect 23661 21947 23719 21953
rect 23661 21944 23673 21947
rect 23624 21916 23673 21944
rect 23624 21904 23630 21916
rect 23661 21913 23673 21916
rect 23707 21913 23719 21947
rect 23661 21907 23719 21913
rect 8481 21879 8539 21885
rect 8481 21845 8493 21879
rect 8527 21876 8539 21879
rect 8662 21876 8668 21888
rect 8527 21848 8668 21876
rect 8527 21845 8539 21848
rect 8481 21839 8539 21845
rect 8662 21836 8668 21848
rect 8720 21836 8726 21888
rect 9030 21836 9036 21888
rect 9088 21836 9094 21888
rect 9306 21836 9312 21888
rect 9364 21836 9370 21888
rect 9858 21836 9864 21888
rect 9916 21876 9922 21888
rect 11422 21876 11428 21888
rect 9916 21848 11428 21876
rect 9916 21836 9922 21848
rect 11422 21836 11428 21848
rect 11480 21836 11486 21888
rect 15102 21836 15108 21888
rect 15160 21876 15166 21888
rect 16666 21876 16672 21888
rect 15160 21848 16672 21876
rect 15160 21836 15166 21848
rect 16666 21836 16672 21848
rect 16724 21836 16730 21888
rect 16761 21879 16819 21885
rect 16761 21845 16773 21879
rect 16807 21876 16819 21879
rect 17678 21876 17684 21888
rect 16807 21848 17684 21876
rect 16807 21845 16819 21848
rect 16761 21839 16819 21845
rect 17678 21836 17684 21848
rect 17736 21836 17742 21888
rect 20165 21879 20223 21885
rect 20165 21845 20177 21879
rect 20211 21876 20223 21879
rect 20254 21876 20260 21888
rect 20211 21848 20260 21876
rect 20211 21845 20223 21848
rect 20165 21839 20223 21845
rect 20254 21836 20260 21848
rect 20312 21836 20318 21888
rect 21726 21836 21732 21888
rect 21784 21876 21790 21888
rect 22922 21876 22928 21888
rect 21784 21848 22928 21876
rect 21784 21836 21790 21848
rect 22922 21836 22928 21848
rect 22980 21836 22986 21888
rect 552 21786 28428 21808
rect 552 21734 3882 21786
rect 3934 21734 3946 21786
rect 3998 21734 4010 21786
rect 4062 21734 4074 21786
rect 4126 21734 4138 21786
rect 4190 21734 10851 21786
rect 10903 21734 10915 21786
rect 10967 21734 10979 21786
rect 11031 21734 11043 21786
rect 11095 21734 11107 21786
rect 11159 21734 17820 21786
rect 17872 21734 17884 21786
rect 17936 21734 17948 21786
rect 18000 21734 18012 21786
rect 18064 21734 18076 21786
rect 18128 21734 24789 21786
rect 24841 21734 24853 21786
rect 24905 21734 24917 21786
rect 24969 21734 24981 21786
rect 25033 21734 25045 21786
rect 25097 21734 28428 21786
rect 552 21712 28428 21734
rect 2406 21632 2412 21684
rect 2464 21632 2470 21684
rect 5445 21675 5503 21681
rect 5445 21641 5457 21675
rect 5491 21672 5503 21675
rect 6914 21672 6920 21684
rect 5491 21644 6920 21672
rect 5491 21641 5503 21644
rect 5445 21635 5503 21641
rect 6914 21632 6920 21644
rect 6972 21672 6978 21684
rect 6972 21644 7512 21672
rect 6972 21632 6978 21644
rect 3053 21607 3111 21613
rect 3053 21573 3065 21607
rect 3099 21573 3111 21607
rect 3053 21567 3111 21573
rect 1029 21471 1087 21477
rect 1029 21437 1041 21471
rect 1075 21468 1087 21471
rect 1118 21468 1124 21480
rect 1075 21440 1124 21468
rect 1075 21437 1087 21440
rect 1029 21431 1087 21437
rect 1118 21428 1124 21440
rect 1176 21428 1182 21480
rect 1296 21471 1354 21477
rect 1296 21437 1308 21471
rect 1342 21468 1354 21471
rect 1762 21468 1768 21480
rect 1342 21440 1768 21468
rect 1342 21437 1354 21440
rect 1296 21431 1354 21437
rect 1762 21428 1768 21440
rect 1820 21428 1826 21480
rect 2777 21471 2835 21477
rect 2777 21437 2789 21471
rect 2823 21468 2835 21471
rect 3068 21468 3096 21567
rect 5166 21564 5172 21616
rect 5224 21604 5230 21616
rect 5350 21604 5356 21616
rect 5224 21576 5356 21604
rect 5224 21564 5230 21576
rect 5350 21564 5356 21576
rect 5408 21564 5414 21616
rect 5534 21536 5540 21548
rect 4908 21508 5540 21536
rect 3237 21471 3295 21477
rect 2823 21440 3004 21468
rect 3068 21440 3188 21468
rect 2823 21437 2835 21440
rect 2777 21431 2835 21437
rect 2866 21292 2872 21344
rect 2924 21292 2930 21344
rect 2976 21332 3004 21440
rect 3050 21360 3056 21412
rect 3108 21360 3114 21412
rect 3160 21400 3188 21440
rect 3237 21437 3249 21471
rect 3283 21468 3295 21471
rect 4908 21468 4936 21508
rect 5534 21496 5540 21508
rect 5592 21496 5598 21548
rect 7024 21508 7236 21536
rect 7024 21480 7052 21508
rect 3283 21440 4936 21468
rect 4985 21471 5043 21477
rect 3283 21437 3295 21440
rect 3237 21431 3295 21437
rect 4985 21437 4997 21471
rect 5031 21468 5043 21471
rect 5261 21471 5319 21477
rect 5261 21468 5273 21471
rect 5031 21440 5273 21468
rect 5031 21437 5043 21440
rect 4985 21431 5043 21437
rect 5261 21437 5273 21440
rect 5307 21437 5319 21471
rect 5261 21431 5319 21437
rect 3482 21403 3540 21409
rect 3482 21400 3494 21403
rect 3160 21372 3494 21400
rect 3482 21369 3494 21372
rect 3528 21369 3540 21403
rect 5000 21400 5028 21431
rect 5350 21428 5356 21480
rect 5408 21468 5414 21480
rect 5445 21471 5503 21477
rect 5445 21468 5457 21471
rect 5408 21440 5457 21468
rect 5408 21428 5414 21440
rect 5445 21437 5457 21440
rect 5491 21437 5503 21471
rect 5445 21431 5503 21437
rect 7006 21428 7012 21480
rect 7064 21428 7070 21480
rect 7098 21428 7104 21480
rect 7156 21428 7162 21480
rect 7208 21477 7236 21508
rect 7484 21477 7512 21644
rect 8294 21632 8300 21684
rect 8352 21672 8358 21684
rect 8573 21675 8631 21681
rect 8573 21672 8585 21675
rect 8352 21644 8585 21672
rect 8352 21632 8358 21644
rect 8573 21641 8585 21644
rect 8619 21641 8631 21675
rect 9306 21672 9312 21684
rect 8573 21635 8631 21641
rect 8864 21644 9312 21672
rect 8389 21607 8447 21613
rect 8389 21573 8401 21607
rect 8435 21604 8447 21607
rect 8864 21604 8892 21644
rect 9306 21632 9312 21644
rect 9364 21632 9370 21684
rect 9401 21675 9459 21681
rect 9401 21641 9413 21675
rect 9447 21672 9459 21675
rect 9582 21672 9588 21684
rect 9447 21644 9588 21672
rect 9447 21641 9459 21644
rect 9401 21635 9459 21641
rect 9582 21632 9588 21644
rect 9640 21632 9646 21684
rect 13998 21632 14004 21684
rect 14056 21672 14062 21684
rect 14185 21675 14243 21681
rect 14185 21672 14197 21675
rect 14056 21644 14197 21672
rect 14056 21632 14062 21644
rect 14185 21641 14197 21644
rect 14231 21641 14243 21675
rect 15654 21672 15660 21684
rect 14185 21635 14243 21641
rect 14384 21644 15660 21672
rect 8435 21576 8892 21604
rect 8956 21576 11744 21604
rect 8435 21573 8447 21576
rect 8389 21567 8447 21573
rect 8018 21496 8024 21548
rect 8076 21496 8082 21548
rect 7193 21471 7251 21477
rect 7193 21437 7205 21471
rect 7239 21437 7251 21471
rect 7193 21431 7251 21437
rect 7469 21471 7527 21477
rect 7469 21437 7481 21471
rect 7515 21437 7527 21471
rect 7469 21431 7527 21437
rect 7742 21428 7748 21480
rect 7800 21428 7806 21480
rect 7837 21471 7895 21477
rect 7837 21437 7849 21471
rect 7883 21437 7895 21471
rect 8036 21468 8064 21496
rect 8386 21468 8392 21480
rect 8036 21440 8392 21468
rect 7837 21431 7895 21437
rect 5810 21409 5816 21412
rect 3482 21363 3540 21369
rect 4632 21372 5028 21400
rect 3326 21332 3332 21344
rect 2976 21304 3332 21332
rect 3326 21292 3332 21304
rect 3384 21292 3390 21344
rect 4632 21341 4660 21372
rect 5804 21363 5816 21409
rect 5810 21360 5816 21363
rect 5868 21360 5874 21412
rect 4617 21335 4675 21341
rect 4617 21301 4629 21335
rect 4663 21301 4675 21335
rect 4617 21295 4675 21301
rect 4798 21292 4804 21344
rect 4856 21292 4862 21344
rect 6730 21292 6736 21344
rect 6788 21332 6794 21344
rect 6917 21335 6975 21341
rect 6917 21332 6929 21335
rect 6788 21304 6929 21332
rect 6788 21292 6794 21304
rect 6917 21301 6929 21304
rect 6963 21332 6975 21335
rect 7852 21332 7880 21431
rect 8386 21428 8392 21440
rect 8444 21468 8450 21480
rect 8573 21471 8631 21477
rect 8573 21468 8585 21471
rect 8444 21440 8585 21468
rect 8444 21428 8450 21440
rect 8573 21437 8585 21440
rect 8619 21437 8631 21471
rect 8573 21431 8631 21437
rect 8662 21428 8668 21480
rect 8720 21428 8726 21480
rect 8956 21477 8984 21576
rect 9306 21496 9312 21548
rect 9364 21536 9370 21548
rect 9364 21508 9812 21536
rect 9364 21496 9370 21508
rect 8941 21471 8999 21477
rect 8941 21437 8953 21471
rect 8987 21437 8999 21471
rect 8941 21431 8999 21437
rect 9030 21428 9036 21480
rect 9088 21468 9094 21480
rect 9539 21471 9597 21477
rect 9539 21468 9551 21471
rect 9088 21440 9551 21468
rect 9088 21428 9094 21440
rect 9539 21437 9551 21440
rect 9585 21437 9597 21471
rect 9784 21468 9812 21508
rect 9858 21496 9864 21548
rect 9916 21536 9922 21548
rect 9916 21508 9996 21536
rect 9916 21496 9922 21508
rect 9968 21477 9996 21508
rect 9952 21471 10010 21477
rect 9784 21440 9904 21468
rect 9539 21431 9597 21437
rect 8680 21400 8708 21428
rect 9677 21403 9735 21409
rect 9677 21400 9689 21403
rect 8680 21372 9689 21400
rect 9600 21344 9628 21372
rect 9677 21369 9689 21372
rect 9723 21369 9735 21403
rect 9677 21363 9735 21369
rect 9769 21403 9827 21409
rect 9769 21369 9781 21403
rect 9815 21369 9827 21403
rect 9876 21400 9904 21440
rect 9952 21437 9964 21471
rect 9998 21437 10010 21471
rect 9952 21431 10010 21437
rect 10042 21428 10048 21480
rect 10100 21428 10106 21480
rect 10321 21471 10379 21477
rect 10321 21468 10333 21471
rect 10152 21440 10333 21468
rect 10152 21400 10180 21440
rect 10321 21437 10333 21440
rect 10367 21437 10379 21471
rect 10321 21431 10379 21437
rect 10502 21428 10508 21480
rect 10560 21428 10566 21480
rect 9876 21372 10180 21400
rect 9769 21363 9827 21369
rect 6963 21304 7880 21332
rect 6963 21301 6975 21304
rect 6917 21295 6975 21301
rect 9582 21292 9588 21344
rect 9640 21292 9646 21344
rect 9784 21332 9812 21363
rect 10226 21360 10232 21412
rect 10284 21400 10290 21412
rect 10413 21403 10471 21409
rect 10413 21400 10425 21403
rect 10284 21372 10425 21400
rect 10284 21360 10290 21372
rect 10413 21369 10425 21372
rect 10459 21369 10471 21403
rect 10413 21363 10471 21369
rect 10318 21332 10324 21344
rect 9784 21304 10324 21332
rect 10318 21292 10324 21304
rect 10376 21292 10382 21344
rect 10520 21332 10548 21428
rect 11716 21400 11744 21576
rect 11882 21564 11888 21616
rect 11940 21564 11946 21616
rect 12066 21536 12072 21548
rect 11808 21508 12072 21536
rect 11808 21477 11836 21508
rect 12066 21496 12072 21508
rect 12124 21536 12130 21548
rect 14384 21545 14412 21644
rect 15654 21632 15660 21644
rect 15712 21632 15718 21684
rect 15838 21632 15844 21684
rect 15896 21672 15902 21684
rect 16209 21675 16267 21681
rect 16209 21672 16221 21675
rect 15896 21644 16221 21672
rect 15896 21632 15902 21644
rect 16209 21641 16221 21644
rect 16255 21641 16267 21675
rect 17218 21672 17224 21684
rect 16209 21635 16267 21641
rect 16316 21644 17224 21672
rect 16316 21604 16344 21644
rect 17218 21632 17224 21644
rect 17276 21632 17282 21684
rect 18874 21632 18880 21684
rect 18932 21672 18938 21684
rect 19153 21675 19211 21681
rect 19153 21672 19165 21675
rect 18932 21644 19165 21672
rect 18932 21632 18938 21644
rect 19153 21641 19165 21644
rect 19199 21641 19211 21675
rect 19153 21635 19211 21641
rect 21082 21632 21088 21684
rect 21140 21672 21146 21684
rect 21269 21675 21327 21681
rect 21269 21672 21281 21675
rect 21140 21644 21281 21672
rect 21140 21632 21146 21644
rect 21269 21641 21281 21644
rect 21315 21641 21327 21675
rect 21269 21635 21327 21641
rect 22005 21675 22063 21681
rect 22005 21641 22017 21675
rect 22051 21672 22063 21675
rect 22738 21672 22744 21684
rect 22051 21644 22744 21672
rect 22051 21641 22063 21644
rect 22005 21635 22063 21641
rect 22738 21632 22744 21644
rect 22796 21632 22802 21684
rect 22830 21632 22836 21684
rect 22888 21672 22894 21684
rect 23201 21675 23259 21681
rect 23201 21672 23213 21675
rect 22888 21644 23213 21672
rect 22888 21632 22894 21644
rect 23201 21641 23213 21644
rect 23247 21672 23259 21675
rect 23247 21644 24155 21672
rect 23247 21641 23259 21644
rect 23201 21635 23259 21641
rect 15764 21576 16344 21604
rect 16393 21607 16451 21613
rect 14369 21539 14427 21545
rect 12124 21508 14320 21536
rect 12124 21496 12130 21508
rect 11793 21471 11851 21477
rect 11793 21437 11805 21471
rect 11839 21437 11851 21471
rect 11793 21431 11851 21437
rect 11977 21471 12035 21477
rect 11977 21437 11989 21471
rect 12023 21468 12035 21471
rect 12023 21440 12434 21468
rect 12023 21437 12035 21440
rect 11977 21431 12035 21437
rect 12406 21400 12434 21440
rect 12710 21428 12716 21480
rect 12768 21468 12774 21480
rect 14001 21471 14059 21477
rect 14001 21468 14013 21471
rect 12768 21440 14013 21468
rect 12768 21428 12774 21440
rect 14001 21437 14013 21440
rect 14047 21437 14059 21471
rect 14001 21431 14059 21437
rect 14185 21471 14243 21477
rect 14185 21437 14197 21471
rect 14231 21437 14243 21471
rect 14292 21468 14320 21508
rect 14369 21505 14381 21539
rect 14415 21505 14427 21539
rect 14369 21499 14427 21505
rect 15010 21468 15016 21480
rect 14292 21440 15016 21468
rect 14185 21431 14243 21437
rect 14090 21400 14096 21412
rect 11716 21372 12296 21400
rect 12406 21372 14096 21400
rect 11790 21332 11796 21344
rect 10520 21304 11796 21332
rect 11790 21292 11796 21304
rect 11848 21292 11854 21344
rect 12268 21332 12296 21372
rect 14090 21360 14096 21372
rect 14148 21400 14154 21412
rect 14200 21400 14228 21431
rect 15010 21428 15016 21440
rect 15068 21428 15074 21480
rect 14148 21372 14228 21400
rect 14636 21403 14694 21409
rect 14148 21360 14154 21372
rect 14636 21369 14648 21403
rect 14682 21400 14694 21403
rect 14826 21400 14832 21412
rect 14682 21372 14832 21400
rect 14682 21369 14694 21372
rect 14636 21363 14694 21369
rect 14826 21360 14832 21372
rect 14884 21360 14890 21412
rect 15764 21341 15792 21576
rect 16393 21573 16405 21607
rect 16439 21604 16451 21607
rect 17405 21607 17463 21613
rect 17405 21604 17417 21607
rect 16439 21576 17417 21604
rect 16439 21573 16451 21576
rect 16393 21567 16451 21573
rect 17405 21573 17417 21576
rect 17451 21573 17463 21607
rect 17405 21567 17463 21573
rect 22278 21564 22284 21616
rect 22336 21604 22342 21616
rect 24029 21607 24087 21613
rect 24029 21604 24041 21607
rect 22336 21576 24041 21604
rect 22336 21564 22342 21576
rect 17678 21496 17684 21548
rect 17736 21496 17742 21548
rect 18248 21508 19380 21536
rect 16117 21471 16175 21477
rect 16117 21437 16129 21471
rect 16163 21437 16175 21471
rect 16117 21431 16175 21437
rect 16132 21400 16160 21431
rect 16298 21428 16304 21480
rect 16356 21428 16362 21480
rect 16592 21477 16779 21484
rect 16577 21471 16779 21477
rect 16577 21437 16589 21471
rect 16623 21464 16779 21471
rect 16623 21456 16804 21464
rect 16623 21437 16635 21456
rect 16577 21431 16635 21437
rect 16751 21436 16804 21456
rect 16669 21403 16727 21409
rect 16132 21372 16552 21400
rect 15749 21335 15807 21341
rect 15749 21332 15761 21335
rect 12268 21304 15761 21332
rect 15749 21301 15761 21304
rect 15795 21301 15807 21335
rect 15749 21295 15807 21301
rect 15838 21292 15844 21344
rect 15896 21292 15902 21344
rect 16524 21332 16552 21372
rect 16669 21369 16681 21403
rect 16715 21369 16727 21403
rect 16776 21400 16804 21436
rect 17218 21428 17224 21480
rect 17276 21428 17282 21480
rect 17586 21428 17592 21480
rect 17644 21428 17650 21480
rect 17773 21471 17831 21477
rect 17773 21437 17785 21471
rect 17819 21437 17831 21471
rect 17773 21431 17831 21437
rect 17604 21400 17632 21428
rect 16776 21372 17632 21400
rect 17788 21400 17816 21431
rect 18046 21428 18052 21480
rect 18104 21428 18110 21480
rect 18248 21477 18276 21508
rect 19352 21480 19380 21508
rect 20714 21496 20720 21548
rect 20772 21536 20778 21548
rect 20901 21539 20959 21545
rect 20901 21536 20913 21539
rect 20772 21508 20913 21536
rect 20772 21496 20778 21508
rect 20901 21505 20913 21508
rect 20947 21536 20959 21539
rect 22373 21539 22431 21545
rect 20947 21508 21496 21536
rect 20947 21505 20959 21508
rect 20901 21499 20959 21505
rect 18233 21471 18291 21477
rect 18233 21437 18245 21471
rect 18279 21437 18291 21471
rect 18233 21431 18291 21437
rect 18966 21428 18972 21480
rect 19024 21428 19030 21480
rect 19334 21428 19340 21480
rect 19392 21428 19398 21480
rect 20346 21468 20352 21480
rect 19444 21440 20352 21468
rect 18141 21403 18199 21409
rect 18141 21400 18153 21403
rect 17788 21372 18153 21400
rect 16669 21363 16727 21369
rect 18141 21369 18153 21372
rect 18187 21369 18199 21403
rect 18141 21363 18199 21369
rect 16684 21332 16712 21363
rect 16524 21304 16712 21332
rect 16758 21292 16764 21344
rect 16816 21332 16822 21344
rect 19444 21332 19472 21440
rect 20346 21428 20352 21440
rect 20404 21468 20410 21480
rect 20809 21471 20867 21477
rect 20809 21468 20821 21471
rect 20404 21440 20821 21468
rect 20404 21428 20410 21440
rect 20809 21437 20821 21440
rect 20855 21437 20867 21471
rect 20809 21431 20867 21437
rect 19702 21360 19708 21412
rect 19760 21400 19766 21412
rect 19978 21400 19984 21412
rect 19760 21372 19984 21400
rect 19760 21360 19766 21372
rect 19978 21360 19984 21372
rect 20036 21400 20042 21412
rect 20824 21400 20852 21431
rect 20990 21428 20996 21480
rect 21048 21468 21054 21480
rect 21085 21471 21143 21477
rect 21085 21468 21097 21471
rect 21048 21440 21097 21468
rect 21048 21428 21054 21440
rect 21085 21437 21097 21440
rect 21131 21437 21143 21471
rect 21085 21431 21143 21437
rect 21361 21471 21419 21477
rect 21361 21437 21373 21471
rect 21407 21437 21419 21471
rect 21468 21468 21496 21508
rect 22373 21505 22385 21539
rect 22419 21536 22431 21539
rect 22646 21536 22652 21548
rect 22419 21508 22652 21536
rect 22419 21505 22431 21508
rect 22373 21499 22431 21505
rect 22646 21496 22652 21508
rect 22704 21496 22710 21548
rect 22922 21496 22928 21548
rect 22980 21536 22986 21548
rect 23293 21539 23351 21545
rect 23293 21536 23305 21539
rect 22980 21508 23305 21536
rect 22980 21496 22986 21508
rect 23293 21505 23305 21508
rect 23339 21505 23351 21539
rect 23293 21499 23351 21505
rect 21545 21471 21603 21477
rect 21545 21468 21557 21471
rect 21468 21440 21557 21468
rect 21361 21431 21419 21437
rect 21545 21437 21557 21440
rect 21591 21468 21603 21471
rect 21634 21468 21640 21480
rect 21591 21440 21640 21468
rect 21591 21437 21603 21440
rect 21545 21431 21603 21437
rect 21376 21400 21404 21431
rect 21634 21428 21640 21440
rect 21692 21428 21698 21480
rect 22186 21428 22192 21480
rect 22244 21428 22250 21480
rect 20036 21372 20392 21400
rect 20824 21372 21404 21400
rect 23308 21400 23336 21499
rect 23400 21477 23428 21576
rect 24029 21573 24041 21576
rect 24075 21573 24087 21607
rect 24029 21567 24087 21573
rect 23845 21539 23903 21545
rect 23845 21505 23857 21539
rect 23891 21536 23903 21539
rect 24127 21536 24155 21644
rect 24302 21536 24308 21548
rect 23891 21508 24308 21536
rect 23891 21505 23903 21508
rect 23845 21499 23903 21505
rect 24302 21496 24308 21508
rect 24360 21496 24366 21548
rect 23385 21471 23443 21477
rect 23385 21437 23397 21471
rect 23431 21437 23443 21471
rect 23385 21431 23443 21437
rect 24121 21471 24179 21477
rect 24121 21437 24133 21471
rect 24167 21468 24179 21471
rect 25222 21468 25228 21480
rect 24167 21440 25228 21468
rect 24167 21437 24179 21440
rect 24121 21431 24179 21437
rect 24136 21400 24164 21431
rect 25222 21428 25228 21440
rect 25280 21428 25286 21480
rect 23308 21372 24164 21400
rect 20036 21360 20042 21372
rect 16816 21304 19472 21332
rect 16816 21292 16822 21304
rect 19518 21292 19524 21344
rect 19576 21332 19582 21344
rect 20254 21332 20260 21344
rect 19576 21304 20260 21332
rect 19576 21292 19582 21304
rect 20254 21292 20260 21304
rect 20312 21292 20318 21344
rect 20364 21332 20392 21372
rect 21637 21335 21695 21341
rect 21637 21332 21649 21335
rect 20364 21304 21649 21332
rect 21637 21301 21649 21304
rect 21683 21332 21695 21335
rect 21910 21332 21916 21344
rect 21683 21304 21916 21332
rect 21683 21301 21695 21304
rect 21637 21295 21695 21301
rect 21910 21292 21916 21304
rect 21968 21292 21974 21344
rect 23014 21292 23020 21344
rect 23072 21292 23078 21344
rect 23842 21292 23848 21344
rect 23900 21292 23906 21344
rect 552 21242 28587 21264
rect 552 21190 7366 21242
rect 7418 21190 7430 21242
rect 7482 21190 7494 21242
rect 7546 21190 7558 21242
rect 7610 21190 7622 21242
rect 7674 21190 14335 21242
rect 14387 21190 14399 21242
rect 14451 21190 14463 21242
rect 14515 21190 14527 21242
rect 14579 21190 14591 21242
rect 14643 21190 21304 21242
rect 21356 21190 21368 21242
rect 21420 21190 21432 21242
rect 21484 21190 21496 21242
rect 21548 21190 21560 21242
rect 21612 21190 28273 21242
rect 28325 21190 28337 21242
rect 28389 21190 28401 21242
rect 28453 21190 28465 21242
rect 28517 21190 28529 21242
rect 28581 21190 28587 21242
rect 552 21168 28587 21190
rect 1765 21131 1823 21137
rect 1765 21097 1777 21131
rect 1811 21128 1823 21131
rect 1854 21128 1860 21140
rect 1811 21100 1860 21128
rect 1811 21097 1823 21100
rect 1765 21091 1823 21097
rect 1854 21088 1860 21100
rect 1912 21088 1918 21140
rect 3050 21088 3056 21140
rect 3108 21128 3114 21140
rect 3237 21131 3295 21137
rect 3237 21128 3249 21131
rect 3108 21100 3249 21128
rect 3108 21088 3114 21100
rect 3237 21097 3249 21100
rect 3283 21097 3295 21131
rect 3237 21091 3295 21097
rect 5258 21088 5264 21140
rect 5316 21128 5322 21140
rect 5316 21100 5396 21128
rect 5316 21088 5322 21100
rect 5368 21060 5396 21100
rect 5534 21088 5540 21140
rect 5592 21128 5598 21140
rect 9125 21131 9183 21137
rect 9125 21128 9137 21131
rect 5592 21100 9137 21128
rect 5592 21088 5598 21100
rect 9125 21097 9137 21100
rect 9171 21128 9183 21131
rect 9490 21128 9496 21140
rect 9171 21100 9496 21128
rect 9171 21097 9183 21100
rect 9125 21091 9183 21097
rect 9490 21088 9496 21100
rect 9548 21128 9554 21140
rect 9766 21128 9772 21140
rect 9548 21100 9772 21128
rect 9548 21088 9554 21100
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 10318 21088 10324 21140
rect 10376 21128 10382 21140
rect 12526 21128 12532 21140
rect 10376 21100 12532 21128
rect 10376 21088 10382 21100
rect 5000 21032 5396 21060
rect 5000 21004 5028 21032
rect 1670 20952 1676 21004
rect 1728 20992 1734 21004
rect 1728 20964 1808 20992
rect 1728 20952 1734 20964
rect 1780 20933 1808 20964
rect 2038 20952 2044 21004
rect 2096 20952 2102 21004
rect 2866 20952 2872 21004
rect 2924 20992 2930 21004
rect 3513 20995 3571 21001
rect 3513 20992 3525 20995
rect 2924 20964 3525 20992
rect 2924 20952 2930 20964
rect 3513 20961 3525 20964
rect 3559 20992 3571 20995
rect 4798 20992 4804 21004
rect 3559 20964 4804 20992
rect 3559 20961 3571 20964
rect 3513 20955 3571 20961
rect 4798 20952 4804 20964
rect 4856 20952 4862 21004
rect 4982 20952 4988 21004
rect 5040 20952 5046 21004
rect 5368 21001 5396 21032
rect 9674 21020 9680 21072
rect 9732 21020 9738 21072
rect 10428 21069 10456 21100
rect 12526 21088 12532 21100
rect 12584 21088 12590 21140
rect 13538 21088 13544 21140
rect 13596 21128 13602 21140
rect 13596 21100 14412 21128
rect 13596 21088 13602 21100
rect 10413 21063 10471 21069
rect 10413 21029 10425 21063
rect 10459 21029 10471 21063
rect 10413 21023 10471 21029
rect 11149 21063 11207 21069
rect 11149 21029 11161 21063
rect 11195 21060 11207 21063
rect 11514 21060 11520 21072
rect 11195 21032 11520 21060
rect 11195 21029 11207 21032
rect 11149 21023 11207 21029
rect 11514 21020 11520 21032
rect 11572 21020 11578 21072
rect 11974 21020 11980 21072
rect 12032 21020 12038 21072
rect 13906 21060 13912 21072
rect 12544 21032 13912 21060
rect 5261 20995 5319 21001
rect 5261 20961 5273 20995
rect 5307 20961 5319 20995
rect 5261 20955 5319 20961
rect 5353 20995 5411 21001
rect 5353 20961 5365 20995
rect 5399 20961 5411 20995
rect 5353 20955 5411 20961
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20924 1823 20927
rect 3237 20927 3295 20933
rect 3237 20924 3249 20927
rect 1811 20896 3249 20924
rect 1811 20893 1823 20896
rect 1765 20887 1823 20893
rect 3237 20893 3249 20896
rect 3283 20893 3295 20927
rect 3237 20887 3295 20893
rect 1486 20748 1492 20800
rect 1544 20788 1550 20800
rect 1949 20791 2007 20797
rect 1949 20788 1961 20791
rect 1544 20760 1961 20788
rect 1544 20748 1550 20760
rect 1949 20757 1961 20760
rect 1995 20757 2007 20791
rect 3252 20788 3280 20887
rect 5074 20884 5080 20936
rect 5132 20924 5138 20936
rect 5169 20927 5227 20933
rect 5169 20924 5181 20927
rect 5132 20896 5181 20924
rect 5132 20884 5138 20896
rect 5169 20893 5181 20896
rect 5215 20924 5227 20927
rect 5276 20924 5304 20955
rect 5442 20952 5448 21004
rect 5500 20992 5506 21004
rect 5813 20995 5871 21001
rect 5813 20992 5825 20995
rect 5500 20964 5825 20992
rect 5500 20952 5506 20964
rect 5813 20961 5825 20964
rect 5859 20992 5871 20995
rect 6270 20992 6276 21004
rect 5859 20964 6276 20992
rect 5859 20961 5871 20964
rect 5813 20955 5871 20961
rect 6270 20952 6276 20964
rect 6328 20952 6334 21004
rect 7561 20995 7619 21001
rect 7561 20961 7573 20995
rect 7607 20992 7619 20995
rect 7837 20995 7895 21001
rect 7837 20992 7849 20995
rect 7607 20964 7849 20992
rect 7607 20961 7619 20964
rect 7561 20955 7619 20961
rect 7837 20961 7849 20964
rect 7883 20992 7895 20995
rect 8202 20992 8208 21004
rect 7883 20964 8208 20992
rect 7883 20961 7895 20964
rect 7837 20955 7895 20961
rect 8202 20952 8208 20964
rect 8260 20952 8266 21004
rect 10226 20952 10232 21004
rect 10284 20992 10290 21004
rect 12544 21001 12572 21032
rect 13906 21020 13912 21032
rect 13964 21020 13970 21072
rect 14108 21032 14320 21060
rect 12802 21001 12808 21004
rect 11793 20995 11851 21001
rect 11793 20992 11805 20995
rect 10284 20964 11805 20992
rect 10284 20952 10290 20964
rect 11793 20961 11805 20964
rect 11839 20961 11851 20995
rect 11793 20955 11851 20961
rect 12069 20995 12127 21001
rect 12069 20961 12081 20995
rect 12115 20961 12127 20995
rect 12069 20955 12127 20961
rect 12529 20995 12587 21001
rect 12529 20961 12541 20995
rect 12575 20961 12587 20995
rect 12796 20992 12808 21001
rect 12763 20964 12808 20992
rect 12529 20955 12587 20961
rect 12796 20955 12808 20964
rect 5215 20896 5304 20924
rect 5215 20893 5227 20896
rect 5169 20887 5227 20893
rect 5534 20884 5540 20936
rect 5592 20924 5598 20936
rect 5592 20896 6132 20924
rect 5592 20884 5598 20896
rect 6104 20868 6132 20896
rect 9858 20884 9864 20936
rect 9916 20884 9922 20936
rect 9950 20884 9956 20936
rect 10008 20884 10014 20936
rect 10042 20884 10048 20936
rect 10100 20924 10106 20936
rect 11698 20924 11704 20936
rect 10100 20896 11704 20924
rect 10100 20884 10106 20896
rect 3326 20816 3332 20868
rect 3384 20856 3390 20868
rect 3421 20859 3479 20865
rect 3421 20856 3433 20859
rect 3384 20828 3433 20856
rect 3384 20816 3390 20828
rect 3421 20825 3433 20828
rect 3467 20856 3479 20859
rect 4801 20859 4859 20865
rect 4801 20856 4813 20859
rect 3467 20828 4813 20856
rect 3467 20825 3479 20828
rect 3421 20819 3479 20825
rect 4801 20825 4813 20828
rect 4847 20856 4859 20859
rect 4847 20828 6040 20856
rect 4847 20825 4859 20828
rect 4801 20819 4859 20825
rect 6012 20800 6040 20828
rect 6086 20816 6092 20868
rect 6144 20816 6150 20868
rect 10428 20865 10456 20896
rect 11698 20884 11704 20896
rect 11756 20884 11762 20936
rect 11974 20884 11980 20936
rect 12032 20924 12038 20936
rect 12084 20924 12112 20955
rect 12802 20952 12808 20955
rect 12860 20952 12866 21004
rect 14108 20992 14136 21032
rect 13832 20964 14136 20992
rect 12032 20896 12112 20924
rect 12032 20884 12038 20896
rect 10413 20859 10471 20865
rect 10413 20825 10425 20859
rect 10459 20825 10471 20859
rect 10413 20819 10471 20825
rect 10965 20859 11023 20865
rect 10965 20825 10977 20859
rect 11011 20856 11023 20859
rect 11238 20856 11244 20868
rect 11011 20828 11244 20856
rect 11011 20825 11023 20828
rect 10965 20819 11023 20825
rect 11238 20816 11244 20828
rect 11296 20816 11302 20868
rect 11517 20859 11575 20865
rect 11517 20825 11529 20859
rect 11563 20856 11575 20859
rect 11563 20828 12434 20856
rect 11563 20825 11575 20828
rect 11517 20819 11575 20825
rect 3694 20788 3700 20800
rect 3252 20760 3700 20788
rect 1949 20751 2007 20757
rect 3694 20748 3700 20760
rect 3752 20748 3758 20800
rect 5445 20791 5503 20797
rect 5445 20757 5457 20791
rect 5491 20788 5503 20791
rect 5626 20788 5632 20800
rect 5491 20760 5632 20788
rect 5491 20757 5503 20760
rect 5445 20751 5503 20757
rect 5626 20748 5632 20760
rect 5684 20748 5690 20800
rect 5994 20748 6000 20800
rect 6052 20748 6058 20800
rect 11149 20791 11207 20797
rect 11149 20757 11161 20791
rect 11195 20788 11207 20791
rect 11609 20791 11667 20797
rect 11609 20788 11621 20791
rect 11195 20760 11621 20788
rect 11195 20757 11207 20760
rect 11149 20751 11207 20757
rect 11609 20757 11621 20760
rect 11655 20757 11667 20791
rect 12406 20788 12434 20828
rect 13832 20788 13860 20964
rect 14182 20952 14188 21004
rect 14240 20952 14246 21004
rect 13909 20859 13967 20865
rect 13909 20825 13921 20859
rect 13955 20856 13967 20859
rect 14200 20856 14228 20952
rect 14292 20924 14320 21032
rect 14384 21001 14412 21100
rect 14826 21088 14832 21140
rect 14884 21088 14890 21140
rect 15838 21088 15844 21140
rect 15896 21088 15902 21140
rect 16482 21088 16488 21140
rect 16540 21128 16546 21140
rect 18785 21131 18843 21137
rect 16540 21100 18736 21128
rect 16540 21088 16546 21100
rect 14369 20995 14427 21001
rect 14369 20961 14381 20995
rect 14415 20961 14427 20995
rect 14369 20955 14427 20961
rect 15010 20952 15016 21004
rect 15068 20952 15074 21004
rect 15197 20995 15255 21001
rect 15197 20961 15209 20995
rect 15243 20992 15255 20995
rect 15856 20992 15884 21088
rect 16736 21063 16794 21069
rect 16736 21029 16748 21063
rect 16782 21060 16794 21063
rect 17405 21063 17463 21069
rect 17405 21060 17417 21063
rect 16782 21032 17417 21060
rect 16782 21029 16794 21032
rect 16736 21023 16794 21029
rect 17405 21029 17417 21032
rect 17451 21029 17463 21063
rect 17405 21023 17463 21029
rect 17512 21032 17724 21060
rect 15243 20964 15884 20992
rect 15243 20961 15255 20964
rect 15197 20955 15255 20961
rect 17126 20952 17132 21004
rect 17184 20992 17190 21004
rect 17512 21001 17540 21032
rect 17696 21004 17724 21032
rect 17313 20995 17371 21001
rect 17313 20992 17325 20995
rect 17184 20964 17325 20992
rect 17184 20952 17190 20964
rect 17313 20961 17325 20964
rect 17359 20961 17371 20995
rect 17313 20955 17371 20961
rect 17497 20995 17555 21001
rect 17497 20961 17509 20995
rect 17543 20961 17555 20995
rect 17497 20955 17555 20961
rect 17586 20952 17592 21004
rect 17644 20952 17650 21004
rect 17678 20952 17684 21004
rect 17736 20952 17742 21004
rect 18708 20992 18736 21100
rect 18785 21097 18797 21131
rect 18831 21128 18843 21131
rect 18966 21128 18972 21140
rect 18831 21100 18972 21128
rect 18831 21097 18843 21100
rect 18785 21091 18843 21097
rect 18966 21088 18972 21100
rect 19024 21088 19030 21140
rect 19245 21131 19303 21137
rect 19245 21097 19257 21131
rect 19291 21097 19303 21131
rect 19245 21091 19303 21097
rect 19260 21060 19288 21091
rect 20806 21088 20812 21140
rect 20864 21088 20870 21140
rect 22738 21088 22744 21140
rect 22796 21088 22802 21140
rect 23842 21088 23848 21140
rect 23900 21088 23906 21140
rect 19429 21063 19487 21069
rect 19260 21032 19380 21060
rect 19153 20995 19211 21001
rect 19153 20992 19165 20995
rect 18708 20964 19165 20992
rect 19153 20961 19165 20964
rect 19199 20961 19211 20995
rect 19352 20992 19380 21032
rect 19429 21029 19441 21063
rect 19475 21060 19487 21063
rect 19518 21060 19524 21072
rect 19475 21032 19524 21060
rect 19475 21029 19487 21032
rect 19429 21023 19487 21029
rect 19518 21020 19524 21032
rect 19576 21060 19582 21072
rect 19889 21063 19947 21069
rect 19889 21060 19901 21063
rect 19576 21032 19901 21060
rect 19576 21020 19582 21032
rect 19889 21029 19901 21032
rect 19935 21029 19947 21063
rect 19889 21023 19947 21029
rect 19978 21020 19984 21072
rect 20036 21060 20042 21072
rect 20824 21060 20852 21088
rect 21726 21060 21732 21072
rect 20036 21032 20081 21060
rect 20824 21032 21732 21060
rect 20036 21020 20042 21032
rect 21726 21020 21732 21032
rect 21784 21060 21790 21072
rect 22830 21060 22836 21072
rect 21784 21032 22836 21060
rect 21784 21020 21790 21032
rect 19702 20998 19708 21004
rect 19628 20992 19708 20998
rect 19352 20970 19708 20992
rect 19352 20964 19656 20970
rect 19153 20955 19211 20961
rect 15289 20927 15347 20933
rect 15289 20924 15301 20927
rect 14292 20896 15301 20924
rect 15289 20893 15301 20896
rect 15335 20924 15347 20927
rect 15335 20896 16620 20924
rect 15335 20893 15347 20896
rect 15289 20887 15347 20893
rect 16592 20865 16620 20896
rect 16758 20884 16764 20936
rect 16816 20924 16822 20936
rect 16853 20927 16911 20933
rect 16853 20924 16865 20927
rect 16816 20896 16865 20924
rect 16816 20884 16822 20896
rect 16853 20893 16865 20896
rect 16899 20893 16911 20927
rect 16853 20887 16911 20893
rect 16945 20927 17003 20933
rect 16945 20893 16957 20927
rect 16991 20893 17003 20927
rect 16945 20887 17003 20893
rect 17221 20927 17279 20933
rect 17221 20893 17233 20927
rect 17267 20924 17279 20927
rect 17604 20924 17632 20952
rect 17267 20896 17632 20924
rect 18325 20927 18383 20933
rect 17267 20893 17279 20896
rect 17221 20887 17279 20893
rect 18325 20893 18337 20927
rect 18371 20924 18383 20927
rect 18877 20927 18935 20933
rect 18877 20924 18889 20927
rect 18371 20896 18889 20924
rect 18371 20893 18383 20896
rect 18325 20887 18383 20893
rect 18877 20893 18889 20896
rect 18923 20893 18935 20927
rect 18877 20887 18935 20893
rect 13955 20828 14228 20856
rect 16577 20859 16635 20865
rect 13955 20825 13967 20828
rect 13909 20819 13967 20825
rect 16577 20825 16589 20859
rect 16623 20825 16635 20859
rect 16960 20856 16988 20887
rect 18966 20884 18972 20936
rect 19024 20924 19030 20936
rect 19061 20927 19119 20933
rect 19061 20924 19073 20927
rect 19024 20896 19073 20924
rect 19024 20884 19030 20896
rect 19061 20893 19073 20896
rect 19107 20893 19119 20927
rect 19168 20924 19196 20955
rect 19702 20952 19708 20970
rect 19760 20952 19766 21004
rect 19797 20995 19855 21001
rect 19797 20961 19809 20995
rect 19843 20961 19855 20995
rect 19797 20955 19855 20961
rect 19426 20924 19432 20936
rect 19168 20896 19432 20924
rect 19061 20887 19119 20893
rect 19426 20884 19432 20896
rect 19484 20884 19490 20936
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20924 19579 20927
rect 19812 20924 19840 20955
rect 20070 20952 20076 21004
rect 20128 21001 20134 21004
rect 20128 20995 20157 21001
rect 20145 20961 20157 20995
rect 20128 20955 20157 20961
rect 20128 20952 20134 20955
rect 20254 20952 20260 21004
rect 20312 20952 20318 21004
rect 21818 20952 21824 21004
rect 21876 20952 21882 21004
rect 22020 21001 22048 21032
rect 22830 21020 22836 21032
rect 22888 21020 22894 21072
rect 22005 20995 22063 21001
rect 22005 20961 22017 20995
rect 22051 20961 22063 20995
rect 22005 20955 22063 20961
rect 23014 20952 23020 21004
rect 23072 20992 23078 21004
rect 23109 20995 23167 21001
rect 23109 20992 23121 20995
rect 23072 20964 23121 20992
rect 23072 20952 23078 20964
rect 23109 20961 23121 20964
rect 23155 20961 23167 20995
rect 23109 20955 23167 20961
rect 23201 20995 23259 21001
rect 23201 20961 23213 20995
rect 23247 20992 23259 20995
rect 23860 20992 23888 21088
rect 23247 20964 23888 20992
rect 23247 20961 23259 20964
rect 23201 20955 23259 20961
rect 19567 20896 19748 20924
rect 19812 20896 19849 20924
rect 19567 20893 19579 20896
rect 19521 20887 19579 20893
rect 18693 20859 18751 20865
rect 16960 20828 17264 20856
rect 16577 20819 16635 20825
rect 17236 20800 17264 20828
rect 18693 20825 18705 20859
rect 18739 20856 18751 20859
rect 19613 20859 19671 20865
rect 19613 20856 19625 20859
rect 18739 20828 19625 20856
rect 18739 20825 18751 20828
rect 18693 20819 18751 20825
rect 19613 20825 19625 20828
rect 19659 20825 19671 20859
rect 19720 20856 19748 20896
rect 19821 20856 19849 20896
rect 19720 20828 20944 20856
rect 19613 20819 19671 20825
rect 20916 20800 20944 20828
rect 22462 20816 22468 20868
rect 22520 20856 22526 20868
rect 24394 20856 24400 20868
rect 22520 20828 24400 20856
rect 22520 20816 22526 20828
rect 24394 20816 24400 20828
rect 24452 20816 24458 20868
rect 12406 20760 13860 20788
rect 14001 20791 14059 20797
rect 11609 20751 11667 20757
rect 14001 20757 14013 20791
rect 14047 20788 14059 20791
rect 14090 20788 14096 20800
rect 14047 20760 14096 20788
rect 14047 20757 14059 20760
rect 14001 20751 14059 20757
rect 14090 20748 14096 20760
rect 14148 20748 14154 20800
rect 14369 20791 14427 20797
rect 14369 20757 14381 20791
rect 14415 20788 14427 20791
rect 14734 20788 14740 20800
rect 14415 20760 14740 20788
rect 14415 20757 14427 20760
rect 14369 20751 14427 20757
rect 14734 20748 14740 20760
rect 14792 20748 14798 20800
rect 17218 20748 17224 20800
rect 17276 20748 17282 20800
rect 19242 20748 19248 20800
rect 19300 20788 19306 20800
rect 20070 20788 20076 20800
rect 19300 20760 20076 20788
rect 19300 20748 19306 20760
rect 20070 20748 20076 20760
rect 20128 20748 20134 20800
rect 20898 20748 20904 20800
rect 20956 20748 20962 20800
rect 21821 20791 21879 20797
rect 21821 20757 21833 20791
rect 21867 20788 21879 20791
rect 22186 20788 22192 20800
rect 21867 20760 22192 20788
rect 21867 20757 21879 20760
rect 21821 20751 21879 20757
rect 22186 20748 22192 20760
rect 22244 20748 22250 20800
rect 23382 20748 23388 20800
rect 23440 20748 23446 20800
rect 552 20698 28428 20720
rect 552 20646 3882 20698
rect 3934 20646 3946 20698
rect 3998 20646 4010 20698
rect 4062 20646 4074 20698
rect 4126 20646 4138 20698
rect 4190 20646 10851 20698
rect 10903 20646 10915 20698
rect 10967 20646 10979 20698
rect 11031 20646 11043 20698
rect 11095 20646 11107 20698
rect 11159 20646 17820 20698
rect 17872 20646 17884 20698
rect 17936 20646 17948 20698
rect 18000 20646 18012 20698
rect 18064 20646 18076 20698
rect 18128 20646 24789 20698
rect 24841 20646 24853 20698
rect 24905 20646 24917 20698
rect 24969 20646 24981 20698
rect 25033 20646 25045 20698
rect 25097 20646 28428 20698
rect 552 20624 28428 20646
rect 5810 20544 5816 20596
rect 5868 20544 5874 20596
rect 6822 20544 6828 20596
rect 6880 20584 6886 20596
rect 8757 20587 8815 20593
rect 8757 20584 8769 20587
rect 6880 20556 8769 20584
rect 6880 20544 6886 20556
rect 8757 20553 8769 20556
rect 8803 20584 8815 20587
rect 9401 20587 9459 20593
rect 9401 20584 9413 20587
rect 8803 20556 9413 20584
rect 8803 20553 8815 20556
rect 8757 20547 8815 20553
rect 9401 20553 9413 20556
rect 9447 20553 9459 20587
rect 9401 20547 9459 20553
rect 9493 20587 9551 20593
rect 9493 20553 9505 20587
rect 9539 20584 9551 20587
rect 9950 20584 9956 20596
rect 9539 20556 9956 20584
rect 9539 20553 9551 20556
rect 9493 20547 9551 20553
rect 9950 20544 9956 20556
rect 10008 20544 10014 20596
rect 11054 20544 11060 20596
rect 11112 20584 11118 20596
rect 11793 20587 11851 20593
rect 11793 20584 11805 20587
rect 11112 20556 11805 20584
rect 11112 20544 11118 20556
rect 11793 20553 11805 20556
rect 11839 20553 11851 20587
rect 11793 20547 11851 20553
rect 12802 20544 12808 20596
rect 12860 20544 12866 20596
rect 16298 20544 16304 20596
rect 16356 20544 16362 20596
rect 16390 20544 16396 20596
rect 16448 20584 16454 20596
rect 19334 20584 19340 20596
rect 16448 20556 19340 20584
rect 16448 20544 16454 20556
rect 19334 20544 19340 20556
rect 19392 20544 19398 20596
rect 19518 20544 19524 20596
rect 19576 20584 19582 20596
rect 20165 20587 20223 20593
rect 20165 20584 20177 20587
rect 19576 20556 20177 20584
rect 19576 20544 19582 20556
rect 20165 20553 20177 20556
rect 20211 20553 20223 20587
rect 20165 20547 20223 20553
rect 20898 20544 20904 20596
rect 20956 20544 20962 20596
rect 21174 20544 21180 20596
rect 21232 20544 21238 20596
rect 21818 20544 21824 20596
rect 21876 20544 21882 20596
rect 22186 20544 22192 20596
rect 22244 20544 22250 20596
rect 23382 20544 23388 20596
rect 23440 20544 23446 20596
rect 6730 20476 6736 20528
rect 6788 20476 6794 20528
rect 12710 20516 12716 20528
rect 9324 20488 12716 20516
rect 6086 20408 6092 20460
rect 6144 20448 6150 20460
rect 7190 20448 7196 20460
rect 6144 20420 7196 20448
rect 6144 20408 6150 20420
rect 7190 20408 7196 20420
rect 7248 20408 7254 20460
rect 7282 20408 7288 20460
rect 7340 20448 7346 20460
rect 8386 20448 8392 20460
rect 7340 20420 8392 20448
rect 7340 20408 7346 20420
rect 8386 20408 8392 20420
rect 8444 20408 8450 20460
rect 8478 20408 8484 20460
rect 8536 20408 8542 20460
rect 9324 20448 9352 20488
rect 12710 20476 12716 20488
rect 12768 20516 12774 20528
rect 12768 20488 15976 20516
rect 12768 20476 12774 20488
rect 9232 20420 9352 20448
rect 1765 20383 1823 20389
rect 1765 20349 1777 20383
rect 1811 20380 1823 20383
rect 1946 20380 1952 20392
rect 1811 20352 1952 20380
rect 1811 20349 1823 20352
rect 1765 20343 1823 20349
rect 1946 20340 1952 20352
rect 2004 20340 2010 20392
rect 5626 20340 5632 20392
rect 5684 20380 5690 20392
rect 5813 20383 5871 20389
rect 5813 20380 5825 20383
rect 5684 20352 5825 20380
rect 5684 20340 5690 20352
rect 5813 20349 5825 20352
rect 5859 20349 5871 20383
rect 5813 20343 5871 20349
rect 5994 20340 6000 20392
rect 6052 20340 6058 20392
rect 6914 20340 6920 20392
rect 6972 20340 6978 20392
rect 7098 20340 7104 20392
rect 7156 20340 7162 20392
rect 8496 20380 8524 20408
rect 9232 20389 9260 20420
rect 9582 20408 9588 20460
rect 9640 20408 9646 20460
rect 12618 20448 12624 20460
rect 11348 20420 12624 20448
rect 8573 20383 8631 20389
rect 8573 20380 8585 20383
rect 7208 20376 8348 20380
rect 8496 20376 8585 20380
rect 7208 20352 8585 20376
rect 5350 20272 5356 20324
rect 5408 20312 5414 20324
rect 5718 20312 5724 20324
rect 5408 20284 5724 20312
rect 5408 20272 5414 20284
rect 5718 20272 5724 20284
rect 5776 20312 5782 20324
rect 6730 20312 6736 20324
rect 5776 20284 6736 20312
rect 5776 20272 5782 20284
rect 6730 20272 6736 20284
rect 6788 20312 6794 20324
rect 7208 20312 7236 20352
rect 8320 20348 8524 20352
rect 8573 20349 8585 20352
rect 8619 20349 8631 20383
rect 8573 20343 8631 20349
rect 9033 20383 9091 20389
rect 9033 20349 9045 20383
rect 9079 20349 9091 20383
rect 9033 20343 9091 20349
rect 9217 20383 9275 20389
rect 9217 20349 9229 20383
rect 9263 20349 9275 20383
rect 9217 20343 9275 20349
rect 6788 20284 7236 20312
rect 7285 20315 7343 20321
rect 6788 20272 6794 20284
rect 7285 20281 7297 20315
rect 7331 20312 7343 20315
rect 9048 20312 9076 20343
rect 9306 20340 9312 20392
rect 9364 20340 9370 20392
rect 11149 20383 11207 20389
rect 11149 20349 11161 20383
rect 11195 20380 11207 20383
rect 11238 20380 11244 20392
rect 11195 20352 11244 20380
rect 11195 20349 11207 20352
rect 11149 20343 11207 20349
rect 11238 20340 11244 20352
rect 11296 20340 11302 20392
rect 11348 20312 11376 20420
rect 12618 20408 12624 20420
rect 12676 20408 12682 20460
rect 13817 20451 13875 20457
rect 13096 20420 13676 20448
rect 11974 20340 11980 20392
rect 12032 20340 12038 20392
rect 12345 20383 12403 20389
rect 12345 20349 12357 20383
rect 12391 20380 12403 20383
rect 12986 20380 12992 20392
rect 12391 20352 12992 20380
rect 12391 20349 12403 20352
rect 12345 20343 12403 20349
rect 12986 20340 12992 20352
rect 13044 20340 13050 20392
rect 13096 20389 13124 20420
rect 13648 20392 13676 20420
rect 13817 20417 13829 20451
rect 13863 20448 13875 20451
rect 13998 20448 14004 20460
rect 13863 20420 14004 20448
rect 13863 20417 13875 20420
rect 13817 20411 13875 20417
rect 13998 20408 14004 20420
rect 14056 20408 14062 20460
rect 14734 20408 14740 20460
rect 14792 20448 14798 20460
rect 15378 20448 15384 20460
rect 14792 20420 15384 20448
rect 14792 20408 14798 20420
rect 15378 20408 15384 20420
rect 15436 20408 15442 20460
rect 13081 20383 13139 20389
rect 13081 20349 13093 20383
rect 13127 20349 13139 20383
rect 13081 20343 13139 20349
rect 13170 20340 13176 20392
rect 13228 20380 13234 20392
rect 13541 20383 13599 20389
rect 13541 20380 13553 20383
rect 13228 20352 13553 20380
rect 13228 20340 13234 20352
rect 13541 20349 13553 20352
rect 13587 20349 13599 20383
rect 13541 20343 13599 20349
rect 13630 20340 13636 20392
rect 13688 20340 13694 20392
rect 7331 20284 11376 20312
rect 7331 20281 7343 20284
rect 7285 20275 7343 20281
rect 11422 20272 11428 20324
rect 11480 20312 11486 20324
rect 12069 20315 12127 20321
rect 12069 20312 12081 20315
rect 11480 20284 12081 20312
rect 11480 20272 11486 20284
rect 12069 20281 12081 20284
rect 12115 20281 12127 20315
rect 12069 20275 12127 20281
rect 1578 20204 1584 20256
rect 1636 20204 1642 20256
rect 4982 20204 4988 20256
rect 5040 20244 5046 20256
rect 6086 20244 6092 20256
rect 5040 20216 6092 20244
rect 5040 20204 5046 20216
rect 6086 20204 6092 20216
rect 6144 20244 6150 20256
rect 7006 20244 7012 20256
rect 6144 20216 7012 20244
rect 6144 20204 6150 20216
rect 7006 20204 7012 20216
rect 7064 20204 7070 20256
rect 7190 20204 7196 20256
rect 7248 20244 7254 20256
rect 8941 20247 8999 20253
rect 8941 20244 8953 20247
rect 7248 20216 8953 20244
rect 7248 20204 7254 20216
rect 8941 20213 8953 20216
rect 8987 20213 8999 20247
rect 8941 20207 8999 20213
rect 11330 20204 11336 20256
rect 11388 20204 11394 20256
rect 12084 20244 12112 20275
rect 12158 20272 12164 20324
rect 12216 20272 12222 20324
rect 12805 20315 12863 20321
rect 12805 20281 12817 20315
rect 12851 20312 12863 20315
rect 13817 20315 13875 20321
rect 13817 20312 13829 20315
rect 12851 20284 13829 20312
rect 12851 20281 12863 20284
rect 12805 20275 12863 20281
rect 13817 20281 13829 20284
rect 13863 20281 13875 20315
rect 15948 20312 15976 20488
rect 16758 20408 16764 20460
rect 16816 20408 16822 20460
rect 16942 20408 16948 20460
rect 17000 20448 17006 20460
rect 17126 20448 17132 20460
rect 17000 20420 17132 20448
rect 17000 20408 17006 20420
rect 17126 20408 17132 20420
rect 17184 20408 17190 20460
rect 19352 20448 19380 20544
rect 21192 20516 21220 20544
rect 20824 20488 21220 20516
rect 20824 20457 20852 20488
rect 20441 20451 20499 20457
rect 20441 20448 20453 20451
rect 19352 20420 20453 20448
rect 20441 20417 20453 20420
rect 20487 20417 20499 20451
rect 20441 20411 20499 20417
rect 20625 20451 20683 20457
rect 20625 20417 20637 20451
rect 20671 20448 20683 20451
rect 20809 20451 20867 20457
rect 20809 20448 20821 20451
rect 20671 20420 20821 20448
rect 20671 20417 20683 20420
rect 20625 20411 20683 20417
rect 20809 20417 20821 20420
rect 20855 20417 20867 20451
rect 21836 20448 21864 20544
rect 20809 20411 20867 20417
rect 20916 20420 21128 20448
rect 16574 20340 16580 20392
rect 16632 20380 16638 20392
rect 18693 20383 18751 20389
rect 18693 20380 18705 20383
rect 16632 20352 18705 20380
rect 16632 20340 16638 20352
rect 18693 20349 18705 20352
rect 18739 20349 18751 20383
rect 18693 20343 18751 20349
rect 20349 20383 20407 20389
rect 20349 20349 20361 20383
rect 20395 20349 20407 20383
rect 20349 20343 20407 20349
rect 18325 20315 18383 20321
rect 18325 20312 18337 20315
rect 15948 20284 18337 20312
rect 13817 20275 13875 20281
rect 18325 20281 18337 20284
rect 18371 20312 18383 20315
rect 18785 20315 18843 20321
rect 18785 20312 18797 20315
rect 18371 20284 18797 20312
rect 18371 20281 18383 20284
rect 18325 20275 18383 20281
rect 18785 20281 18797 20284
rect 18831 20312 18843 20315
rect 18966 20312 18972 20324
rect 18831 20284 18972 20312
rect 18831 20281 18843 20284
rect 18785 20275 18843 20281
rect 18966 20272 18972 20284
rect 19024 20272 19030 20324
rect 20364 20312 20392 20343
rect 20530 20340 20536 20392
rect 20588 20380 20594 20392
rect 20916 20380 20944 20420
rect 20588 20352 20944 20380
rect 20588 20340 20594 20352
rect 20990 20340 20996 20392
rect 21048 20340 21054 20392
rect 21100 20389 21128 20420
rect 21652 20420 21864 20448
rect 22373 20451 22431 20457
rect 21652 20389 21680 20420
rect 22373 20417 22385 20451
rect 22419 20448 22431 20451
rect 23400 20448 23428 20544
rect 22419 20420 23428 20448
rect 22419 20417 22431 20420
rect 22373 20411 22431 20417
rect 21085 20383 21143 20389
rect 21085 20349 21097 20383
rect 21131 20349 21143 20383
rect 21085 20343 21143 20349
rect 21637 20383 21695 20389
rect 21637 20349 21649 20383
rect 21683 20349 21695 20383
rect 21637 20343 21695 20349
rect 21726 20340 21732 20392
rect 21784 20340 21790 20392
rect 22094 20340 22100 20392
rect 22152 20340 22158 20392
rect 22462 20340 22468 20392
rect 22520 20340 22526 20392
rect 22833 20383 22891 20389
rect 22833 20349 22845 20383
rect 22879 20380 22891 20383
rect 23474 20380 23480 20392
rect 22879 20352 23480 20380
rect 22879 20349 22891 20352
rect 22833 20343 22891 20349
rect 23474 20340 23480 20352
rect 23532 20340 23538 20392
rect 21453 20315 21511 20321
rect 21453 20312 21465 20315
rect 20364 20284 21465 20312
rect 21453 20281 21465 20284
rect 21499 20281 21511 20315
rect 21453 20275 21511 20281
rect 12342 20244 12348 20256
rect 12084 20216 12348 20244
rect 12342 20204 12348 20216
rect 12400 20204 12406 20256
rect 12894 20204 12900 20256
rect 12952 20244 12958 20256
rect 12989 20247 13047 20253
rect 12989 20244 13001 20247
rect 12952 20216 13001 20244
rect 12952 20204 12958 20216
rect 12989 20213 13001 20216
rect 13035 20244 13047 20247
rect 13170 20244 13176 20256
rect 13035 20216 13176 20244
rect 13035 20213 13047 20216
rect 12989 20207 13047 20213
rect 13170 20204 13176 20216
rect 13228 20204 13234 20256
rect 14826 20204 14832 20256
rect 14884 20204 14890 20256
rect 16669 20247 16727 20253
rect 16669 20213 16681 20247
rect 16715 20244 16727 20247
rect 17218 20244 17224 20256
rect 16715 20216 17224 20244
rect 16715 20213 16727 20216
rect 16669 20207 16727 20213
rect 17218 20204 17224 20216
rect 17276 20204 17282 20256
rect 18049 20247 18107 20253
rect 18049 20213 18061 20247
rect 18095 20244 18107 20247
rect 18138 20244 18144 20256
rect 18095 20216 18144 20244
rect 18095 20213 18107 20216
rect 18049 20207 18107 20213
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 21468 20244 21496 20275
rect 21634 20244 21640 20256
rect 21468 20216 21640 20244
rect 21634 20204 21640 20216
rect 21692 20204 21698 20256
rect 21744 20244 21772 20340
rect 22373 20315 22431 20321
rect 22373 20281 22385 20315
rect 22419 20312 22431 20315
rect 22649 20315 22707 20321
rect 22649 20312 22661 20315
rect 22419 20284 22661 20312
rect 22419 20281 22431 20284
rect 22373 20275 22431 20281
rect 22649 20281 22661 20284
rect 22695 20281 22707 20315
rect 22649 20275 22707 20281
rect 22741 20315 22799 20321
rect 22741 20281 22753 20315
rect 22787 20281 22799 20315
rect 22741 20275 22799 20281
rect 22756 20244 22784 20275
rect 21744 20216 22784 20244
rect 22830 20204 22836 20256
rect 22888 20244 22894 20256
rect 23017 20247 23075 20253
rect 23017 20244 23029 20247
rect 22888 20216 23029 20244
rect 22888 20204 22894 20216
rect 23017 20213 23029 20216
rect 23063 20213 23075 20247
rect 23017 20207 23075 20213
rect 552 20154 28587 20176
rect 552 20102 7366 20154
rect 7418 20102 7430 20154
rect 7482 20102 7494 20154
rect 7546 20102 7558 20154
rect 7610 20102 7622 20154
rect 7674 20102 14335 20154
rect 14387 20102 14399 20154
rect 14451 20102 14463 20154
rect 14515 20102 14527 20154
rect 14579 20102 14591 20154
rect 14643 20102 21304 20154
rect 21356 20102 21368 20154
rect 21420 20102 21432 20154
rect 21484 20102 21496 20154
rect 21548 20102 21560 20154
rect 21612 20102 28273 20154
rect 28325 20102 28337 20154
rect 28389 20102 28401 20154
rect 28453 20102 28465 20154
rect 28517 20102 28529 20154
rect 28581 20102 28587 20154
rect 552 20080 28587 20102
rect 4341 20043 4399 20049
rect 3068 20012 4292 20040
rect 1578 19981 1584 19984
rect 1572 19972 1584 19981
rect 1539 19944 1584 19972
rect 1572 19935 1584 19944
rect 1578 19932 1584 19935
rect 1636 19932 1642 19984
rect 1118 19864 1124 19916
rect 1176 19904 1182 19916
rect 1305 19907 1363 19913
rect 1305 19904 1317 19907
rect 1176 19876 1317 19904
rect 1176 19864 1182 19876
rect 1305 19873 1317 19876
rect 1351 19873 1363 19907
rect 1305 19867 1363 19873
rect 2961 19771 3019 19777
rect 2961 19768 2973 19771
rect 2240 19740 2973 19768
rect 1486 19660 1492 19712
rect 1544 19700 1550 19712
rect 2240 19700 2268 19740
rect 2961 19737 2973 19740
rect 3007 19737 3019 19771
rect 2961 19731 3019 19737
rect 1544 19672 2268 19700
rect 2685 19703 2743 19709
rect 1544 19660 1550 19672
rect 2685 19669 2697 19703
rect 2731 19700 2743 19703
rect 2866 19700 2872 19712
rect 2731 19672 2872 19700
rect 2731 19669 2743 19672
rect 2685 19663 2743 19669
rect 2866 19660 2872 19672
rect 2924 19700 2930 19712
rect 3068 19700 3096 20012
rect 3129 19975 3187 19981
rect 3129 19941 3141 19975
rect 3175 19972 3187 19975
rect 3329 19975 3387 19981
rect 3175 19944 3280 19972
rect 3175 19941 3187 19944
rect 3129 19935 3187 19941
rect 3252 19904 3280 19944
rect 3329 19941 3341 19975
rect 3375 19972 3387 19975
rect 3602 19972 3608 19984
rect 3375 19944 3608 19972
rect 3375 19941 3387 19944
rect 3329 19935 3387 19941
rect 3602 19932 3608 19944
rect 3660 19932 3666 19984
rect 4264 19972 4292 20012
rect 4341 20009 4353 20043
rect 4387 20040 4399 20043
rect 4801 20043 4859 20049
rect 4801 20040 4813 20043
rect 4387 20012 4813 20040
rect 4387 20009 4399 20012
rect 4341 20003 4399 20009
rect 4801 20009 4813 20012
rect 4847 20009 4859 20043
rect 4801 20003 4859 20009
rect 6641 20043 6699 20049
rect 6641 20009 6653 20043
rect 6687 20040 6699 20043
rect 7006 20040 7012 20052
rect 6687 20012 7012 20040
rect 6687 20009 6699 20012
rect 6641 20003 6699 20009
rect 7006 20000 7012 20012
rect 7064 20000 7070 20052
rect 7101 20043 7159 20049
rect 7101 20009 7113 20043
rect 7147 20040 7159 20043
rect 7285 20043 7343 20049
rect 7285 20040 7297 20043
rect 7147 20012 7297 20040
rect 7147 20009 7159 20012
rect 7101 20003 7159 20009
rect 7285 20009 7297 20012
rect 7331 20009 7343 20043
rect 7285 20003 7343 20009
rect 7561 20043 7619 20049
rect 7561 20009 7573 20043
rect 7607 20009 7619 20043
rect 7561 20003 7619 20009
rect 8389 20043 8447 20049
rect 8389 20009 8401 20043
rect 8435 20040 8447 20043
rect 9030 20040 9036 20052
rect 8435 20012 9036 20040
rect 8435 20009 8447 20012
rect 8389 20003 8447 20009
rect 6457 19975 6515 19981
rect 6457 19972 6469 19975
rect 4264 19944 6469 19972
rect 6457 19941 6469 19944
rect 6503 19972 6515 19975
rect 6503 19944 7328 19972
rect 6503 19941 6515 19944
rect 6457 19935 6515 19941
rect 3252 19876 3832 19904
rect 3804 19780 3832 19876
rect 4798 19864 4804 19916
rect 4856 19904 4862 19916
rect 5169 19907 5227 19913
rect 5169 19904 5181 19907
rect 4856 19876 5181 19904
rect 4856 19864 4862 19876
rect 5169 19873 5181 19876
rect 5215 19904 5227 19907
rect 6089 19907 6147 19913
rect 5215 19876 5856 19904
rect 5215 19873 5227 19876
rect 5169 19867 5227 19873
rect 4982 19796 4988 19848
rect 5040 19796 5046 19848
rect 5074 19796 5080 19848
rect 5132 19796 5138 19848
rect 5261 19839 5319 19845
rect 5261 19805 5273 19839
rect 5307 19836 5319 19839
rect 5718 19836 5724 19848
rect 5307 19808 5724 19836
rect 5307 19805 5319 19808
rect 5261 19799 5319 19805
rect 5718 19796 5724 19808
rect 5776 19796 5782 19848
rect 5828 19836 5856 19876
rect 6089 19873 6101 19907
rect 6135 19904 6147 19907
rect 6178 19904 6184 19916
rect 6135 19876 6184 19904
rect 6135 19873 6147 19876
rect 6089 19867 6147 19873
rect 6178 19864 6184 19876
rect 6236 19864 6242 19916
rect 6730 19864 6736 19916
rect 6788 19864 6794 19916
rect 6914 19864 6920 19916
rect 6972 19904 6978 19916
rect 7193 19907 7251 19913
rect 7193 19904 7205 19907
rect 6972 19876 7205 19904
rect 6972 19864 6978 19876
rect 7193 19873 7205 19876
rect 7239 19873 7251 19907
rect 7300 19904 7328 19944
rect 7374 19932 7380 19984
rect 7432 19981 7438 19984
rect 7432 19975 7454 19981
rect 7442 19941 7454 19975
rect 7576 19972 7604 20003
rect 9030 20000 9036 20012
rect 9088 20040 9094 20052
rect 9306 20040 9312 20052
rect 9088 20012 9312 20040
rect 9088 20000 9094 20012
rect 9306 20000 9312 20012
rect 9364 20000 9370 20052
rect 11330 20000 11336 20052
rect 11388 20000 11394 20052
rect 11974 20000 11980 20052
rect 12032 20040 12038 20052
rect 12345 20043 12403 20049
rect 12345 20040 12357 20043
rect 12032 20012 12357 20040
rect 12032 20000 12038 20012
rect 12345 20009 12357 20012
rect 12391 20009 12403 20043
rect 12345 20003 12403 20009
rect 12986 20000 12992 20052
rect 13044 20040 13050 20052
rect 13262 20040 13268 20052
rect 13044 20012 13268 20040
rect 13044 20000 13050 20012
rect 13262 20000 13268 20012
rect 13320 20000 13326 20052
rect 13538 20000 13544 20052
rect 13596 20000 13602 20052
rect 13630 20000 13636 20052
rect 13688 20000 13694 20052
rect 13801 20043 13859 20049
rect 13801 20009 13813 20043
rect 13847 20040 13859 20043
rect 14734 20040 14740 20052
rect 13847 20012 14740 20040
rect 13847 20009 13859 20012
rect 13801 20003 13859 20009
rect 14734 20000 14740 20012
rect 14792 20040 14798 20052
rect 14918 20040 14924 20052
rect 14792 20012 14924 20040
rect 14792 20000 14798 20012
rect 14918 20000 14924 20012
rect 14976 20000 14982 20052
rect 15378 20000 15384 20052
rect 15436 20040 15442 20052
rect 15473 20043 15531 20049
rect 15473 20040 15485 20043
rect 15436 20012 15485 20040
rect 15436 20000 15442 20012
rect 15473 20009 15485 20012
rect 15519 20009 15531 20043
rect 15473 20003 15531 20009
rect 16390 20000 16396 20052
rect 16448 20000 16454 20052
rect 16669 20043 16727 20049
rect 16669 20009 16681 20043
rect 16715 20040 16727 20043
rect 16758 20040 16764 20052
rect 16715 20012 16764 20040
rect 16715 20009 16727 20012
rect 16669 20003 16727 20009
rect 16758 20000 16764 20012
rect 16816 20000 16822 20052
rect 17218 20000 17224 20052
rect 17276 20000 17282 20052
rect 20717 20043 20775 20049
rect 20717 20009 20729 20043
rect 20763 20040 20775 20043
rect 20990 20040 20996 20052
rect 20763 20012 20996 20040
rect 20763 20009 20775 20012
rect 20717 20003 20775 20009
rect 20990 20000 20996 20012
rect 21048 20000 21054 20052
rect 21453 20043 21511 20049
rect 21453 20009 21465 20043
rect 21499 20009 21511 20043
rect 21453 20003 21511 20009
rect 8570 19972 8576 19984
rect 7576 19944 8576 19972
rect 7432 19935 7454 19941
rect 7432 19932 7438 19935
rect 8570 19932 8576 19944
rect 8628 19932 8634 19984
rect 11232 19975 11290 19981
rect 11232 19941 11244 19975
rect 11278 19972 11290 19975
rect 11348 19972 11376 20000
rect 13648 19972 13676 20000
rect 14001 19975 14059 19981
rect 14001 19972 14013 19975
rect 11278 19944 11376 19972
rect 13096 19944 13676 19972
rect 13832 19944 14013 19972
rect 11278 19941 11290 19944
rect 11232 19935 11290 19941
rect 8021 19907 8079 19913
rect 8021 19904 8033 19907
rect 7300 19876 8033 19904
rect 7193 19867 7251 19873
rect 8021 19873 8033 19876
rect 8067 19904 8079 19907
rect 8110 19904 8116 19916
rect 8067 19876 8116 19904
rect 8067 19873 8079 19876
rect 8021 19867 8079 19873
rect 8110 19864 8116 19876
rect 8168 19864 8174 19916
rect 8205 19907 8263 19913
rect 8205 19873 8217 19907
rect 8251 19873 8263 19907
rect 8205 19867 8263 19873
rect 6825 19839 6883 19845
rect 6825 19836 6837 19839
rect 5828 19808 6837 19836
rect 6825 19805 6837 19808
rect 6871 19836 6883 19839
rect 7282 19836 7288 19848
rect 6871 19808 7288 19836
rect 6871 19805 6883 19808
rect 6825 19799 6883 19805
rect 7282 19796 7288 19808
rect 7340 19796 7346 19848
rect 7561 19839 7619 19845
rect 7561 19805 7573 19839
rect 7607 19836 7619 19839
rect 8220 19836 8248 19867
rect 9766 19864 9772 19916
rect 9824 19864 9830 19916
rect 9950 19864 9956 19916
rect 10008 19864 10014 19916
rect 10045 19907 10103 19913
rect 10045 19873 10057 19907
rect 10091 19904 10103 19907
rect 12802 19904 12808 19916
rect 10091 19876 12808 19904
rect 10091 19873 10103 19876
rect 10045 19867 10103 19873
rect 12802 19864 12808 19876
rect 12860 19864 12866 19916
rect 13096 19913 13124 19944
rect 13832 19916 13860 19944
rect 14001 19941 14013 19944
rect 14047 19972 14059 19975
rect 16114 19972 16120 19984
rect 14047 19944 16120 19972
rect 14047 19941 14059 19944
rect 14001 19935 14059 19941
rect 16114 19932 16120 19944
rect 16172 19932 16178 19984
rect 16408 19972 16436 20000
rect 21468 19972 21496 20003
rect 22094 20000 22100 20052
rect 22152 20000 22158 20052
rect 23014 20000 23020 20052
rect 23072 20000 23078 20052
rect 24302 20000 24308 20052
rect 24360 20000 24366 20052
rect 21910 19972 21916 19984
rect 16408 19944 16896 19972
rect 13081 19907 13139 19913
rect 13081 19873 13093 19907
rect 13127 19873 13139 19907
rect 13081 19867 13139 19873
rect 13170 19864 13176 19916
rect 13228 19864 13234 19916
rect 13814 19864 13820 19916
rect 13872 19864 13878 19916
rect 13906 19864 13912 19916
rect 13964 19904 13970 19916
rect 14093 19907 14151 19913
rect 14093 19904 14105 19907
rect 13964 19876 14105 19904
rect 13964 19864 13970 19876
rect 14093 19873 14105 19876
rect 14139 19873 14151 19907
rect 14093 19867 14151 19873
rect 14182 19864 14188 19916
rect 14240 19904 14246 19916
rect 14349 19907 14407 19913
rect 14349 19904 14361 19907
rect 14240 19876 14361 19904
rect 14240 19864 14246 19876
rect 14349 19873 14361 19876
rect 14395 19873 14407 19907
rect 14349 19867 14407 19873
rect 16209 19907 16267 19913
rect 16209 19873 16221 19907
rect 16255 19904 16267 19907
rect 16408 19904 16436 19944
rect 16255 19876 16436 19904
rect 16761 19907 16819 19913
rect 16255 19873 16267 19876
rect 16209 19867 16267 19873
rect 16761 19873 16773 19907
rect 16807 19873 16819 19907
rect 16761 19867 16819 19873
rect 7607 19808 8248 19836
rect 9784 19836 9812 19864
rect 10965 19839 11023 19845
rect 10965 19836 10977 19839
rect 9784 19808 10977 19836
rect 7607 19805 7619 19808
rect 7561 19799 7619 19805
rect 3786 19728 3792 19780
rect 3844 19768 3850 19780
rect 3973 19771 4031 19777
rect 3973 19768 3985 19771
rect 3844 19740 3985 19768
rect 3844 19728 3850 19740
rect 3973 19737 3985 19740
rect 4019 19737 4031 19771
rect 3973 19731 4031 19737
rect 4356 19740 4660 19768
rect 4356 19709 4384 19740
rect 3145 19703 3203 19709
rect 3145 19700 3157 19703
rect 2924 19672 3157 19700
rect 2924 19660 2930 19672
rect 3145 19669 3157 19672
rect 3191 19669 3203 19703
rect 3145 19663 3203 19669
rect 4341 19703 4399 19709
rect 4341 19669 4353 19703
rect 4387 19700 4399 19703
rect 4430 19700 4436 19712
rect 4387 19672 4436 19700
rect 4387 19669 4399 19672
rect 4341 19663 4399 19669
rect 4430 19660 4436 19672
rect 4488 19660 4494 19712
rect 4522 19660 4528 19712
rect 4580 19660 4586 19712
rect 4632 19700 4660 19740
rect 6656 19740 6868 19768
rect 6656 19712 6684 19740
rect 5534 19700 5540 19712
rect 4632 19672 5540 19700
rect 5534 19660 5540 19672
rect 5592 19660 5598 19712
rect 6454 19660 6460 19712
rect 6512 19660 6518 19712
rect 6638 19660 6644 19712
rect 6696 19660 6702 19712
rect 6840 19709 6868 19740
rect 8036 19712 8064 19808
rect 10965 19805 10977 19808
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 6825 19703 6883 19709
rect 6825 19669 6837 19703
rect 6871 19669 6883 19703
rect 6825 19663 6883 19669
rect 8018 19660 8024 19712
rect 8076 19660 8082 19712
rect 10137 19703 10195 19709
rect 10137 19669 10149 19703
rect 10183 19700 10195 19703
rect 10226 19700 10232 19712
rect 10183 19672 10232 19700
rect 10183 19669 10195 19672
rect 10137 19663 10195 19669
rect 10226 19660 10232 19672
rect 10284 19660 10290 19712
rect 10318 19660 10324 19712
rect 10376 19660 10382 19712
rect 10980 19700 11008 19799
rect 12894 19796 12900 19848
rect 12952 19836 12958 19848
rect 13265 19839 13323 19845
rect 13265 19836 13277 19839
rect 12952 19808 13277 19836
rect 12952 19796 12958 19808
rect 13265 19805 13277 19808
rect 13311 19805 13323 19839
rect 13265 19799 13323 19805
rect 13630 19796 13636 19848
rect 13688 19836 13694 19848
rect 16776 19836 16804 19867
rect 13688 19808 14136 19836
rect 13688 19796 13694 19808
rect 13446 19768 13452 19780
rect 12544 19740 13452 19768
rect 12544 19712 12572 19740
rect 13446 19728 13452 19740
rect 13504 19768 13510 19780
rect 13504 19740 13860 19768
rect 13504 19728 13510 19740
rect 11238 19700 11244 19712
rect 10980 19672 11244 19700
rect 11238 19660 11244 19672
rect 11296 19660 11302 19712
rect 12526 19660 12532 19712
rect 12584 19660 12590 19712
rect 12986 19660 12992 19712
rect 13044 19660 13050 19712
rect 13262 19660 13268 19712
rect 13320 19700 13326 19712
rect 13630 19700 13636 19712
rect 13320 19672 13636 19700
rect 13320 19660 13326 19672
rect 13630 19660 13636 19672
rect 13688 19660 13694 19712
rect 13832 19709 13860 19740
rect 13817 19703 13875 19709
rect 13817 19669 13829 19703
rect 13863 19669 13875 19703
rect 14108 19700 14136 19808
rect 16316 19808 16804 19836
rect 16316 19709 16344 19808
rect 16868 19709 16896 19944
rect 20916 19944 21496 19972
rect 21836 19944 21916 19972
rect 20916 19913 20944 19944
rect 18877 19907 18935 19913
rect 18877 19873 18889 19907
rect 18923 19904 18935 19907
rect 19521 19907 19579 19913
rect 19521 19904 19533 19907
rect 18923 19876 19533 19904
rect 18923 19873 18935 19876
rect 18877 19867 18935 19873
rect 19521 19873 19533 19876
rect 19567 19873 19579 19907
rect 19521 19867 19579 19873
rect 20901 19907 20959 19913
rect 20901 19873 20913 19907
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 21085 19907 21143 19913
rect 21085 19873 21097 19907
rect 21131 19873 21143 19907
rect 21085 19867 21143 19873
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 20070 19836 20076 19848
rect 19392 19808 20076 19836
rect 19392 19796 19398 19808
rect 20070 19796 20076 19808
rect 20128 19836 20134 19848
rect 20916 19836 20944 19867
rect 20128 19808 20944 19836
rect 20128 19796 20134 19808
rect 21100 19768 21128 19867
rect 21174 19864 21180 19916
rect 21232 19904 21238 19916
rect 21269 19907 21327 19913
rect 21269 19904 21281 19907
rect 21232 19876 21281 19904
rect 21232 19864 21238 19876
rect 21269 19873 21281 19876
rect 21315 19873 21327 19907
rect 21269 19867 21327 19873
rect 21545 19907 21603 19913
rect 21545 19873 21557 19907
rect 21591 19904 21603 19907
rect 21634 19904 21640 19916
rect 21591 19876 21640 19904
rect 21591 19873 21603 19876
rect 21545 19867 21603 19873
rect 21284 19836 21312 19867
rect 21634 19864 21640 19876
rect 21692 19904 21698 19916
rect 21729 19907 21787 19913
rect 21729 19904 21741 19907
rect 21692 19876 21741 19904
rect 21692 19864 21698 19876
rect 21729 19873 21741 19876
rect 21775 19873 21787 19907
rect 21729 19867 21787 19873
rect 21836 19836 21864 19944
rect 21910 19932 21916 19944
rect 21968 19932 21974 19984
rect 22278 19904 22284 19916
rect 21284 19808 21864 19836
rect 22066 19876 22284 19904
rect 22066 19768 22094 19876
rect 22278 19864 22284 19876
rect 22336 19904 22342 19916
rect 23032 19904 23060 20000
rect 23198 19913 23204 19916
rect 22336 19876 23060 19904
rect 22336 19864 22342 19876
rect 23192 19867 23204 19913
rect 23198 19864 23204 19867
rect 23256 19864 23262 19916
rect 22922 19796 22928 19848
rect 22980 19796 22986 19848
rect 21100 19740 22094 19768
rect 16301 19703 16359 19709
rect 16301 19700 16313 19703
rect 14108 19672 16313 19700
rect 13817 19663 13875 19669
rect 16301 19669 16313 19672
rect 16347 19669 16359 19703
rect 16301 19663 16359 19669
rect 16853 19703 16911 19709
rect 16853 19669 16865 19703
rect 16899 19669 16911 19703
rect 16853 19663 16911 19669
rect 18230 19660 18236 19712
rect 18288 19700 18294 19712
rect 18785 19703 18843 19709
rect 18785 19700 18797 19703
rect 18288 19672 18797 19700
rect 18288 19660 18294 19672
rect 18785 19669 18797 19672
rect 18831 19700 18843 19703
rect 18874 19700 18880 19712
rect 18831 19672 18880 19700
rect 18831 19669 18843 19672
rect 18785 19663 18843 19669
rect 18874 19660 18880 19672
rect 18932 19660 18938 19712
rect 21266 19660 21272 19712
rect 21324 19660 21330 19712
rect 552 19610 28428 19632
rect 552 19558 3882 19610
rect 3934 19558 3946 19610
rect 3998 19558 4010 19610
rect 4062 19558 4074 19610
rect 4126 19558 4138 19610
rect 4190 19558 10851 19610
rect 10903 19558 10915 19610
rect 10967 19558 10979 19610
rect 11031 19558 11043 19610
rect 11095 19558 11107 19610
rect 11159 19558 17820 19610
rect 17872 19558 17884 19610
rect 17936 19558 17948 19610
rect 18000 19558 18012 19610
rect 18064 19558 18076 19610
rect 18128 19558 24789 19610
rect 24841 19558 24853 19610
rect 24905 19558 24917 19610
rect 24969 19558 24981 19610
rect 25033 19558 25045 19610
rect 25097 19558 28428 19610
rect 552 19536 28428 19558
rect 1670 19456 1676 19508
rect 1728 19496 1734 19508
rect 1765 19499 1823 19505
rect 1765 19496 1777 19499
rect 1728 19468 1777 19496
rect 1728 19456 1734 19468
rect 1765 19465 1777 19468
rect 1811 19465 1823 19499
rect 1765 19459 1823 19465
rect 1946 19456 1952 19508
rect 2004 19456 2010 19508
rect 3694 19456 3700 19508
rect 3752 19496 3758 19508
rect 4430 19496 4436 19508
rect 3752 19468 4436 19496
rect 3752 19456 3758 19468
rect 4430 19456 4436 19468
rect 4488 19456 4494 19508
rect 5537 19499 5595 19505
rect 5537 19465 5549 19499
rect 5583 19496 5595 19499
rect 5718 19496 5724 19508
rect 5583 19468 5724 19496
rect 5583 19465 5595 19468
rect 5537 19459 5595 19465
rect 5718 19456 5724 19468
rect 5776 19456 5782 19508
rect 6089 19499 6147 19505
rect 6089 19465 6101 19499
rect 6135 19465 6147 19499
rect 6089 19459 6147 19465
rect 1397 19431 1455 19437
rect 1397 19397 1409 19431
rect 1443 19428 1455 19431
rect 1486 19428 1492 19440
rect 1443 19400 1492 19428
rect 1443 19397 1455 19400
rect 1397 19391 1455 19397
rect 1486 19388 1492 19400
rect 1544 19388 1550 19440
rect 2516 19332 3188 19360
rect 2409 19295 2467 19301
rect 2409 19261 2421 19295
rect 2455 19292 2467 19295
rect 2516 19292 2544 19332
rect 2455 19264 2544 19292
rect 2593 19295 2651 19301
rect 2455 19261 2467 19264
rect 2409 19255 2467 19261
rect 2593 19261 2605 19295
rect 2639 19292 2651 19295
rect 3160 19292 3188 19332
rect 3602 19320 3608 19372
rect 3660 19320 3666 19372
rect 3712 19369 3740 19456
rect 3697 19363 3755 19369
rect 3697 19329 3709 19363
rect 3743 19329 3755 19363
rect 3697 19323 3755 19329
rect 3421 19295 3479 19301
rect 2639 19264 3096 19292
rect 3160 19264 3372 19292
rect 2639 19261 2651 19264
rect 2593 19255 2651 19261
rect 1765 19227 1823 19233
rect 1765 19193 1777 19227
rect 1811 19224 1823 19227
rect 2685 19227 2743 19233
rect 2685 19224 2697 19227
rect 1811 19196 2697 19224
rect 1811 19193 1823 19196
rect 1765 19187 1823 19193
rect 2685 19193 2697 19196
rect 2731 19193 2743 19227
rect 2685 19187 2743 19193
rect 2866 19184 2872 19236
rect 2924 19184 2930 19236
rect 3068 19233 3096 19264
rect 3053 19227 3111 19233
rect 3053 19193 3065 19227
rect 3099 19224 3111 19227
rect 3237 19227 3295 19233
rect 3237 19224 3249 19227
rect 3099 19196 3249 19224
rect 3099 19193 3111 19196
rect 3053 19187 3111 19193
rect 3237 19193 3249 19196
rect 3283 19193 3295 19227
rect 3344 19224 3372 19264
rect 3421 19261 3433 19295
rect 3467 19292 3479 19295
rect 3786 19292 3792 19304
rect 3467 19264 3792 19292
rect 3467 19261 3479 19264
rect 3421 19255 3479 19261
rect 3786 19252 3792 19264
rect 3844 19292 3850 19304
rect 3881 19295 3939 19301
rect 3881 19292 3893 19295
rect 3844 19264 3893 19292
rect 3844 19252 3850 19264
rect 3881 19261 3893 19264
rect 3927 19261 3939 19295
rect 3881 19255 3939 19261
rect 3697 19227 3755 19233
rect 3697 19224 3709 19227
rect 3344 19196 3709 19224
rect 3237 19187 3295 19193
rect 3697 19193 3709 19196
rect 3743 19193 3755 19227
rect 3697 19187 3755 19193
rect 2130 19116 2136 19168
rect 2188 19156 2194 19168
rect 2501 19159 2559 19165
rect 2501 19156 2513 19159
rect 2188 19128 2513 19156
rect 2188 19116 2194 19128
rect 2501 19125 2513 19128
rect 2547 19125 2559 19159
rect 3896 19156 3924 19255
rect 3970 19252 3976 19304
rect 4028 19252 4034 19304
rect 4157 19295 4215 19301
rect 4157 19261 4169 19295
rect 4203 19292 4215 19295
rect 5442 19292 5448 19304
rect 4203 19264 5448 19292
rect 4203 19261 4215 19264
rect 4157 19255 4215 19261
rect 5442 19252 5448 19264
rect 5500 19252 5506 19304
rect 6104 19292 6132 19459
rect 6454 19456 6460 19508
rect 6512 19456 6518 19508
rect 6914 19456 6920 19508
rect 6972 19456 6978 19508
rect 8110 19456 8116 19508
rect 8168 19456 8174 19508
rect 8202 19456 8208 19508
rect 8260 19496 8266 19508
rect 16025 19499 16083 19505
rect 8260 19468 13768 19496
rect 8260 19456 8266 19468
rect 6472 19428 6500 19456
rect 7374 19428 7380 19440
rect 6472 19400 7380 19428
rect 7374 19388 7380 19400
rect 7432 19388 7438 19440
rect 8128 19428 8156 19456
rect 13740 19440 13768 19468
rect 16025 19465 16037 19499
rect 16071 19496 16083 19499
rect 16942 19496 16948 19508
rect 16071 19468 16948 19496
rect 16071 19465 16083 19468
rect 16025 19459 16083 19465
rect 16942 19456 16948 19468
rect 17000 19456 17006 19508
rect 20070 19456 20076 19508
rect 20128 19456 20134 19508
rect 20533 19499 20591 19505
rect 20533 19465 20545 19499
rect 20579 19496 20591 19499
rect 21266 19496 21272 19508
rect 20579 19468 21272 19496
rect 20579 19465 20591 19468
rect 20533 19459 20591 19465
rect 21266 19456 21272 19468
rect 21324 19456 21330 19508
rect 21821 19499 21879 19505
rect 21821 19465 21833 19499
rect 21867 19496 21879 19499
rect 22094 19496 22100 19508
rect 21867 19468 22100 19496
rect 21867 19465 21879 19468
rect 21821 19459 21879 19465
rect 22094 19456 22100 19468
rect 22152 19456 22158 19508
rect 23198 19456 23204 19508
rect 23256 19456 23262 19508
rect 9582 19428 9588 19440
rect 8128 19400 8800 19428
rect 6178 19320 6184 19372
rect 6236 19360 6242 19372
rect 8018 19360 8024 19372
rect 6236 19332 8024 19360
rect 6236 19320 6242 19332
rect 8018 19320 8024 19332
rect 8076 19320 8082 19372
rect 6641 19295 6699 19301
rect 6641 19292 6653 19295
rect 6104 19264 6653 19292
rect 6641 19261 6653 19264
rect 6687 19292 6699 19295
rect 6822 19292 6828 19304
rect 6687 19264 6828 19292
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 6917 19295 6975 19301
rect 6917 19261 6929 19295
rect 6963 19292 6975 19295
rect 8128 19292 8156 19400
rect 8665 19363 8723 19369
rect 8665 19329 8677 19363
rect 8711 19329 8723 19363
rect 8665 19323 8723 19329
rect 6963 19264 8156 19292
rect 6963 19261 6975 19264
rect 6917 19255 6975 19261
rect 4424 19227 4482 19233
rect 4424 19193 4436 19227
rect 4470 19224 4482 19227
rect 4890 19224 4896 19236
rect 4470 19196 4896 19224
rect 4470 19193 4482 19196
rect 4424 19187 4482 19193
rect 4890 19184 4896 19196
rect 4948 19184 4954 19236
rect 5074 19184 5080 19236
rect 5132 19224 5138 19236
rect 6273 19227 6331 19233
rect 6273 19224 6285 19227
rect 5132 19196 6285 19224
rect 5132 19184 5138 19196
rect 6273 19193 6285 19196
rect 6319 19224 6331 19227
rect 6733 19227 6791 19233
rect 6733 19224 6745 19227
rect 6319 19196 6745 19224
rect 6319 19193 6331 19196
rect 6273 19187 6331 19193
rect 6656 19168 6684 19196
rect 6733 19193 6745 19196
rect 6779 19193 6791 19227
rect 6733 19187 6791 19193
rect 8680 19168 8708 19323
rect 8772 19301 8800 19400
rect 9416 19400 9588 19428
rect 9416 19301 9444 19400
rect 9582 19388 9588 19400
rect 9640 19388 9646 19440
rect 9677 19431 9735 19437
rect 9677 19397 9689 19431
rect 9723 19428 9735 19431
rect 9950 19428 9956 19440
rect 9723 19400 9956 19428
rect 9723 19397 9735 19400
rect 9677 19391 9735 19397
rect 9950 19388 9956 19400
rect 10008 19388 10014 19440
rect 10042 19388 10048 19440
rect 10100 19388 10106 19440
rect 13081 19431 13139 19437
rect 13081 19397 13093 19431
rect 13127 19428 13139 19431
rect 13170 19428 13176 19440
rect 13127 19400 13176 19428
rect 13127 19397 13139 19400
rect 13081 19391 13139 19397
rect 13170 19388 13176 19400
rect 13228 19388 13234 19440
rect 13722 19388 13728 19440
rect 13780 19428 13786 19440
rect 14001 19431 14059 19437
rect 14001 19428 14013 19431
rect 13780 19400 14013 19428
rect 13780 19388 13786 19400
rect 14001 19397 14013 19400
rect 14047 19428 14059 19431
rect 17402 19428 17408 19440
rect 14047 19400 17408 19428
rect 14047 19397 14059 19400
rect 14001 19391 14059 19397
rect 17402 19388 17408 19400
rect 17460 19428 17466 19440
rect 17460 19400 18552 19428
rect 17460 19388 17466 19400
rect 18524 19372 18552 19400
rect 20714 19388 20720 19440
rect 20772 19388 20778 19440
rect 9493 19363 9551 19369
rect 9493 19329 9505 19363
rect 9539 19329 9551 19363
rect 9493 19323 9551 19329
rect 8757 19295 8815 19301
rect 8757 19261 8769 19295
rect 8803 19261 8815 19295
rect 8757 19255 8815 19261
rect 9401 19295 9459 19301
rect 9401 19261 9413 19295
rect 9447 19261 9459 19295
rect 9508 19292 9536 19323
rect 11238 19320 11244 19372
rect 11296 19360 11302 19372
rect 11296 19332 11744 19360
rect 11296 19320 11302 19332
rect 9766 19292 9772 19304
rect 9508 19264 9772 19292
rect 9401 19255 9459 19261
rect 9766 19252 9772 19264
rect 9824 19252 9830 19304
rect 9861 19295 9919 19301
rect 9861 19261 9873 19295
rect 9907 19292 9919 19295
rect 9950 19292 9956 19304
rect 9907 19264 9956 19292
rect 9907 19261 9919 19264
rect 9861 19255 9919 19261
rect 9950 19252 9956 19264
rect 10008 19252 10014 19304
rect 11716 19301 11744 19332
rect 12802 19320 12808 19372
rect 12860 19360 12866 19372
rect 13538 19360 13544 19372
rect 12860 19332 13544 19360
rect 12860 19320 12866 19332
rect 13538 19320 13544 19332
rect 13596 19320 13602 19372
rect 15749 19363 15807 19369
rect 15749 19329 15761 19363
rect 15795 19329 15807 19363
rect 15749 19323 15807 19329
rect 17880 19332 18460 19360
rect 10137 19295 10195 19301
rect 10137 19261 10149 19295
rect 10183 19292 10195 19295
rect 10321 19295 10379 19301
rect 10321 19292 10333 19295
rect 10183 19264 10333 19292
rect 10183 19261 10195 19264
rect 10137 19255 10195 19261
rect 10321 19261 10333 19264
rect 10367 19261 10379 19295
rect 10321 19255 10379 19261
rect 10413 19295 10471 19301
rect 10413 19261 10425 19295
rect 10459 19292 10471 19295
rect 11701 19295 11759 19301
rect 10459 19264 11008 19292
rect 10459 19261 10471 19264
rect 10413 19255 10471 19261
rect 10980 19168 11008 19264
rect 11701 19261 11713 19295
rect 11747 19261 11759 19295
rect 11701 19255 11759 19261
rect 15378 19252 15384 19304
rect 15436 19292 15442 19304
rect 15657 19295 15715 19301
rect 15657 19292 15669 19295
rect 15436 19264 15669 19292
rect 15436 19252 15442 19264
rect 15657 19261 15669 19264
rect 15703 19261 15715 19295
rect 15764 19292 15792 19323
rect 17402 19292 17408 19304
rect 15764 19264 17408 19292
rect 15657 19255 15715 19261
rect 17402 19252 17408 19264
rect 17460 19252 17466 19304
rect 17678 19252 17684 19304
rect 17736 19292 17742 19304
rect 17880 19292 17908 19332
rect 17736 19264 17908 19292
rect 17736 19252 17742 19264
rect 17954 19252 17960 19304
rect 18012 19252 18018 19304
rect 18046 19252 18052 19304
rect 18104 19252 18110 19304
rect 18230 19252 18236 19304
rect 18288 19252 18294 19304
rect 18322 19252 18328 19304
rect 18380 19252 18386 19304
rect 18432 19292 18460 19332
rect 18506 19320 18512 19372
rect 18564 19320 18570 19372
rect 20162 19320 20168 19372
rect 20220 19360 20226 19372
rect 20625 19363 20683 19369
rect 20625 19360 20637 19363
rect 20220 19332 20637 19360
rect 20220 19320 20226 19332
rect 20625 19329 20637 19332
rect 20671 19329 20683 19363
rect 22189 19363 22247 19369
rect 22189 19360 22201 19363
rect 20625 19323 20683 19329
rect 22020 19332 22201 19360
rect 18693 19295 18751 19301
rect 18693 19292 18705 19295
rect 18432 19264 18705 19292
rect 18693 19261 18705 19264
rect 18739 19261 18751 19295
rect 18693 19255 18751 19261
rect 18892 19264 19334 19292
rect 11974 19233 11980 19236
rect 11968 19187 11980 19233
rect 11974 19184 11980 19187
rect 12032 19184 12038 19236
rect 15010 19224 15016 19236
rect 13372 19196 15016 19224
rect 13372 19168 13400 19196
rect 15010 19184 15016 19196
rect 15068 19184 15074 19236
rect 15289 19227 15347 19233
rect 15289 19193 15301 19227
rect 15335 19224 15347 19227
rect 18892 19224 18920 19264
rect 15335 19196 18920 19224
rect 18960 19227 19018 19233
rect 15335 19193 15347 19196
rect 15289 19187 15347 19193
rect 18960 19193 18972 19227
rect 19006 19193 19018 19227
rect 19306 19224 19334 19264
rect 20990 19252 20996 19304
rect 21048 19252 21054 19304
rect 21542 19252 21548 19304
rect 21600 19252 21606 19304
rect 21790 19292 21956 19294
rect 22020 19292 22048 19332
rect 22189 19329 22201 19332
rect 22235 19329 22247 19363
rect 22189 19323 22247 19329
rect 21790 19266 22048 19292
rect 21560 19224 21588 19252
rect 19306 19196 21588 19224
rect 21790 19233 21818 19266
rect 21928 19264 22048 19266
rect 22094 19252 22100 19304
rect 22152 19252 22158 19304
rect 22278 19252 22284 19304
rect 22336 19252 22342 19304
rect 22554 19252 22560 19304
rect 22612 19252 22618 19304
rect 22741 19295 22799 19301
rect 22741 19261 22753 19295
rect 22787 19292 22799 19295
rect 22830 19292 22836 19304
rect 22787 19264 22836 19292
rect 22787 19261 22799 19264
rect 22741 19255 22799 19261
rect 22830 19252 22836 19264
rect 22888 19252 22894 19304
rect 22925 19295 22983 19301
rect 22925 19261 22937 19295
rect 22971 19292 22983 19295
rect 23385 19295 23443 19301
rect 23385 19292 23397 19295
rect 22971 19264 23397 19292
rect 22971 19261 22983 19264
rect 22925 19255 22983 19261
rect 23385 19261 23397 19264
rect 23431 19261 23443 19295
rect 23385 19255 23443 19261
rect 21790 19227 21863 19233
rect 21790 19196 21817 19227
rect 18960 19187 19018 19193
rect 21805 19193 21817 19196
rect 21851 19193 21863 19227
rect 21805 19187 21863 19193
rect 6086 19165 6092 19168
rect 5905 19159 5963 19165
rect 5905 19156 5917 19159
rect 3896 19128 5917 19156
rect 2501 19119 2559 19125
rect 5905 19125 5917 19128
rect 5951 19125 5963 19159
rect 5905 19119 5963 19125
rect 6073 19159 6092 19165
rect 6073 19125 6085 19159
rect 6073 19119 6092 19125
rect 6086 19116 6092 19119
rect 6144 19116 6150 19168
rect 6638 19116 6644 19168
rect 6696 19116 6702 19168
rect 8386 19116 8392 19168
rect 8444 19116 8450 19168
rect 8662 19116 8668 19168
rect 8720 19116 8726 19168
rect 9030 19116 9036 19168
rect 9088 19116 9094 19168
rect 10962 19116 10968 19168
rect 11020 19116 11026 19168
rect 13354 19116 13360 19168
rect 13412 19116 13418 19168
rect 13998 19116 14004 19168
rect 14056 19156 14062 19168
rect 16574 19156 16580 19168
rect 14056 19128 16580 19156
rect 14056 19116 14062 19128
rect 16574 19116 16580 19128
rect 16632 19116 16638 19168
rect 18509 19159 18567 19165
rect 18509 19125 18521 19159
rect 18555 19156 18567 19159
rect 18984 19156 19012 19187
rect 21910 19184 21916 19236
rect 21968 19224 21974 19236
rect 22005 19227 22063 19233
rect 22005 19224 22017 19227
rect 21968 19196 22017 19224
rect 21968 19184 21974 19196
rect 22005 19193 22017 19196
rect 22051 19193 22063 19227
rect 22005 19187 22063 19193
rect 18555 19128 19012 19156
rect 20257 19159 20315 19165
rect 18555 19125 18567 19128
rect 18509 19119 18567 19125
rect 20257 19125 20269 19159
rect 20303 19156 20315 19159
rect 20438 19156 20444 19168
rect 20303 19128 20444 19156
rect 20303 19125 20315 19128
rect 20257 19119 20315 19125
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 20901 19159 20959 19165
rect 20901 19125 20913 19159
rect 20947 19156 20959 19159
rect 21174 19156 21180 19168
rect 20947 19128 21180 19156
rect 20947 19125 20959 19128
rect 20901 19119 20959 19125
rect 21174 19116 21180 19128
rect 21232 19116 21238 19168
rect 21634 19116 21640 19168
rect 21692 19116 21698 19168
rect 552 19066 28587 19088
rect 552 19014 7366 19066
rect 7418 19014 7430 19066
rect 7482 19014 7494 19066
rect 7546 19014 7558 19066
rect 7610 19014 7622 19066
rect 7674 19014 14335 19066
rect 14387 19014 14399 19066
rect 14451 19014 14463 19066
rect 14515 19014 14527 19066
rect 14579 19014 14591 19066
rect 14643 19014 21304 19066
rect 21356 19014 21368 19066
rect 21420 19014 21432 19066
rect 21484 19014 21496 19066
rect 21548 19014 21560 19066
rect 21612 19014 28273 19066
rect 28325 19014 28337 19066
rect 28389 19014 28401 19066
rect 28453 19014 28465 19066
rect 28517 19014 28529 19066
rect 28581 19014 28587 19066
rect 552 18992 28587 19014
rect 3970 18912 3976 18964
rect 4028 18952 4034 18964
rect 4157 18955 4215 18961
rect 4157 18952 4169 18955
rect 4028 18924 4169 18952
rect 4028 18912 4034 18924
rect 4157 18921 4169 18924
rect 4203 18921 4215 18955
rect 4157 18915 4215 18921
rect 4522 18912 4528 18964
rect 4580 18912 4586 18964
rect 4890 18912 4896 18964
rect 4948 18912 4954 18964
rect 5442 18912 5448 18964
rect 5500 18952 5506 18964
rect 8754 18952 8760 18964
rect 5500 18924 8760 18952
rect 5500 18912 5506 18924
rect 8754 18912 8760 18924
rect 8812 18912 8818 18964
rect 11790 18912 11796 18964
rect 11848 18912 11854 18964
rect 11974 18912 11980 18964
rect 12032 18912 12038 18964
rect 12986 18912 12992 18964
rect 13044 18952 13050 18964
rect 13044 18924 13768 18952
rect 13044 18912 13050 18924
rect 3602 18776 3608 18828
rect 3660 18776 3666 18828
rect 4433 18819 4491 18825
rect 4433 18785 4445 18819
rect 4479 18785 4491 18819
rect 4540 18816 4568 18912
rect 8849 18887 8907 18893
rect 8849 18884 8861 18887
rect 8680 18856 8861 18884
rect 8680 18828 8708 18856
rect 8849 18853 8861 18856
rect 8895 18853 8907 18887
rect 8849 18847 8907 18853
rect 9030 18844 9036 18896
rect 9088 18844 9094 18896
rect 13170 18844 13176 18896
rect 13228 18844 13234 18896
rect 13354 18844 13360 18896
rect 13412 18844 13418 18896
rect 5077 18819 5135 18825
rect 5077 18816 5089 18819
rect 4540 18788 5089 18816
rect 4433 18779 4491 18785
rect 5077 18785 5089 18788
rect 5123 18785 5135 18819
rect 5077 18779 5135 18785
rect 4448 18680 4476 18779
rect 6730 18776 6736 18828
rect 6788 18776 6794 18828
rect 8662 18776 8668 18828
rect 8720 18776 8726 18828
rect 8757 18819 8815 18825
rect 8757 18785 8769 18819
rect 8803 18785 8815 18819
rect 8757 18779 8815 18785
rect 6825 18751 6883 18757
rect 6825 18717 6837 18751
rect 6871 18748 6883 18751
rect 7098 18748 7104 18760
rect 6871 18720 7104 18748
rect 6871 18717 6883 18720
rect 6825 18711 6883 18717
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 8772 18748 8800 18779
rect 9582 18776 9588 18828
rect 9640 18816 9646 18828
rect 10962 18816 10968 18828
rect 9640 18788 10968 18816
rect 9640 18776 9646 18788
rect 10962 18776 10968 18788
rect 11020 18776 11026 18828
rect 11609 18819 11667 18825
rect 11609 18785 11621 18819
rect 11655 18816 11667 18819
rect 11701 18819 11759 18825
rect 11701 18816 11713 18819
rect 11655 18788 11713 18816
rect 11655 18785 11667 18788
rect 11609 18779 11667 18785
rect 11701 18785 11713 18788
rect 11747 18785 11759 18819
rect 11701 18779 11759 18785
rect 11885 18819 11943 18825
rect 11885 18785 11897 18819
rect 11931 18785 11943 18819
rect 11885 18779 11943 18785
rect 11900 18748 11928 18779
rect 12158 18776 12164 18828
rect 12216 18776 12222 18828
rect 12986 18776 12992 18828
rect 13044 18816 13050 18828
rect 13372 18816 13400 18844
rect 13633 18819 13691 18825
rect 13633 18816 13645 18819
rect 13044 18788 13645 18816
rect 13044 18776 13050 18788
rect 13633 18785 13645 18788
rect 13679 18785 13691 18819
rect 13740 18816 13768 18924
rect 14182 18912 14188 18964
rect 14240 18952 14246 18964
rect 14277 18955 14335 18961
rect 14277 18952 14289 18955
rect 14240 18924 14289 18952
rect 14240 18912 14246 18924
rect 14277 18921 14289 18924
rect 14323 18921 14335 18955
rect 17954 18952 17960 18964
rect 14277 18915 14335 18921
rect 16776 18924 17960 18952
rect 13817 18819 13875 18825
rect 13817 18816 13829 18819
rect 13740 18788 13829 18816
rect 13633 18779 13691 18785
rect 13817 18785 13829 18788
rect 13863 18785 13875 18819
rect 13817 18779 13875 18785
rect 13909 18819 13967 18825
rect 13909 18785 13921 18819
rect 13955 18785 13967 18819
rect 13909 18779 13967 18785
rect 14001 18819 14059 18825
rect 14001 18785 14013 18819
rect 14047 18816 14059 18819
rect 14826 18816 14832 18828
rect 14047 18788 14832 18816
rect 14047 18785 14059 18788
rect 14001 18779 14059 18785
rect 13262 18748 13268 18760
rect 8772 18720 8984 18748
rect 11900 18720 13268 18748
rect 8956 18692 8984 18720
rect 13262 18708 13268 18720
rect 13320 18708 13326 18760
rect 13354 18708 13360 18760
rect 13412 18748 13418 18760
rect 13924 18748 13952 18779
rect 14826 18776 14832 18788
rect 14884 18776 14890 18828
rect 13412 18720 13952 18748
rect 13412 18708 13418 18720
rect 4706 18680 4712 18692
rect 4448 18652 4712 18680
rect 4706 18640 4712 18652
rect 4764 18680 4770 18692
rect 8846 18680 8852 18692
rect 4764 18652 8852 18680
rect 4764 18640 4770 18652
rect 8846 18640 8852 18652
rect 8904 18640 8910 18692
rect 8938 18640 8944 18692
rect 8996 18640 9002 18692
rect 13538 18640 13544 18692
rect 13596 18680 13602 18692
rect 16776 18680 16804 18924
rect 17954 18912 17960 18924
rect 18012 18912 18018 18964
rect 18046 18912 18052 18964
rect 18104 18952 18110 18964
rect 18699 18955 18757 18961
rect 18699 18952 18711 18955
rect 18104 18924 18711 18952
rect 18104 18912 18110 18924
rect 18699 18921 18711 18924
rect 18745 18921 18757 18955
rect 18699 18915 18757 18921
rect 18785 18955 18843 18961
rect 18785 18921 18797 18955
rect 18831 18952 18843 18955
rect 18874 18952 18880 18964
rect 18831 18924 18880 18952
rect 18831 18921 18843 18924
rect 18785 18915 18843 18921
rect 18874 18912 18880 18924
rect 18932 18912 18938 18964
rect 21634 18952 21640 18964
rect 18984 18924 21640 18952
rect 17402 18844 17408 18896
rect 17460 18844 17466 18896
rect 18322 18844 18328 18896
rect 18380 18884 18386 18896
rect 18601 18887 18659 18893
rect 18601 18884 18613 18887
rect 18380 18856 18613 18884
rect 18380 18844 18386 18856
rect 18601 18853 18613 18856
rect 18647 18884 18659 18887
rect 18984 18884 19012 18924
rect 21634 18912 21640 18924
rect 21692 18912 21698 18964
rect 18647 18856 19012 18884
rect 20349 18887 20407 18893
rect 18647 18853 18659 18856
rect 18601 18847 18659 18853
rect 20349 18853 20361 18887
rect 20395 18884 20407 18887
rect 20717 18887 20775 18893
rect 20717 18884 20729 18887
rect 20395 18856 20729 18884
rect 20395 18853 20407 18856
rect 20349 18847 20407 18853
rect 20717 18853 20729 18856
rect 20763 18853 20775 18887
rect 20717 18847 20775 18853
rect 20806 18844 20812 18896
rect 20864 18884 20870 18896
rect 20864 18856 21036 18884
rect 20864 18844 20870 18856
rect 16850 18776 16856 18828
rect 16908 18776 16914 18828
rect 17313 18819 17371 18825
rect 17313 18816 17325 18819
rect 17236 18788 17325 18816
rect 17236 18757 17264 18788
rect 17313 18785 17325 18788
rect 17359 18785 17371 18819
rect 17313 18779 17371 18785
rect 16945 18751 17003 18757
rect 16945 18717 16957 18751
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 17221 18751 17279 18757
rect 17221 18717 17233 18751
rect 17267 18717 17279 18751
rect 17420 18748 17448 18844
rect 17494 18776 17500 18828
rect 17552 18776 17558 18828
rect 17586 18776 17592 18828
rect 17644 18776 17650 18828
rect 18877 18819 18935 18825
rect 18877 18785 18889 18819
rect 18923 18816 18935 18819
rect 19242 18816 19248 18828
rect 18923 18788 19248 18816
rect 18923 18785 18935 18788
rect 18877 18779 18935 18785
rect 19242 18776 19248 18788
rect 19300 18776 19306 18828
rect 20257 18819 20315 18825
rect 20257 18785 20269 18819
rect 20303 18816 20315 18819
rect 20530 18816 20536 18828
rect 20303 18788 20536 18816
rect 20303 18785 20315 18788
rect 20257 18779 20315 18785
rect 20272 18748 20300 18779
rect 20530 18776 20536 18788
rect 20588 18816 20594 18828
rect 21008 18825 21036 18856
rect 23290 18844 23296 18896
rect 23348 18884 23354 18896
rect 23569 18887 23627 18893
rect 23569 18884 23581 18887
rect 23348 18856 23581 18884
rect 23348 18844 23354 18856
rect 23569 18853 23581 18856
rect 23615 18853 23627 18887
rect 23569 18847 23627 18853
rect 20901 18819 20959 18825
rect 20588 18788 20760 18816
rect 20588 18776 20594 18788
rect 20732 18760 20760 18788
rect 20901 18785 20913 18819
rect 20947 18785 20959 18819
rect 20901 18779 20959 18785
rect 20993 18819 21051 18825
rect 20993 18785 21005 18819
rect 21039 18785 21051 18819
rect 20993 18779 21051 18785
rect 22005 18819 22063 18825
rect 22005 18785 22017 18819
rect 22051 18816 22063 18819
rect 23750 18816 23756 18828
rect 22051 18788 23756 18816
rect 22051 18785 22063 18788
rect 22005 18779 22063 18785
rect 17420 18720 20300 18748
rect 17221 18711 17279 18717
rect 13596 18652 16804 18680
rect 16960 18680 16988 18711
rect 20438 18708 20444 18760
rect 20496 18708 20502 18760
rect 20714 18708 20720 18760
rect 20772 18708 20778 18760
rect 20916 18748 20944 18779
rect 23750 18776 23756 18788
rect 23808 18816 23814 18828
rect 23845 18819 23903 18825
rect 23845 18816 23857 18819
rect 23808 18788 23857 18816
rect 23808 18776 23814 18788
rect 23845 18785 23857 18788
rect 23891 18785 23903 18819
rect 23845 18779 23903 18785
rect 21910 18748 21916 18760
rect 20916 18720 21916 18748
rect 21910 18708 21916 18720
rect 21968 18708 21974 18760
rect 20530 18680 20536 18692
rect 16960 18652 20536 18680
rect 13596 18640 13602 18652
rect 20530 18640 20536 18652
rect 20588 18640 20594 18692
rect 4525 18615 4583 18621
rect 4525 18581 4537 18615
rect 4571 18612 4583 18615
rect 4890 18612 4896 18624
rect 4571 18584 4896 18612
rect 4571 18581 4583 18584
rect 4525 18575 4583 18581
rect 4890 18572 4896 18584
rect 4948 18612 4954 18624
rect 5442 18612 5448 18624
rect 4948 18584 5448 18612
rect 4948 18572 4954 18584
rect 5442 18572 5448 18584
rect 5500 18572 5506 18624
rect 7006 18572 7012 18624
rect 7064 18572 7070 18624
rect 8754 18572 8760 18624
rect 8812 18612 8818 18624
rect 9033 18615 9091 18621
rect 9033 18612 9045 18615
rect 8812 18584 9045 18612
rect 8812 18572 8818 18584
rect 9033 18581 9045 18584
rect 9079 18581 9091 18615
rect 9033 18575 9091 18581
rect 12618 18572 12624 18624
rect 12676 18612 12682 18624
rect 13265 18615 13323 18621
rect 13265 18612 13277 18615
rect 12676 18584 13277 18612
rect 12676 18572 12682 18584
rect 13265 18581 13277 18584
rect 13311 18612 13323 18615
rect 13814 18612 13820 18624
rect 13311 18584 13820 18612
rect 13311 18581 13323 18584
rect 13265 18575 13323 18581
rect 13814 18572 13820 18584
rect 13872 18572 13878 18624
rect 17313 18615 17371 18621
rect 17313 18581 17325 18615
rect 17359 18612 17371 18615
rect 17402 18612 17408 18624
rect 17359 18584 17408 18612
rect 17359 18581 17371 18584
rect 17313 18575 17371 18581
rect 17402 18572 17408 18584
rect 17460 18572 17466 18624
rect 19886 18572 19892 18624
rect 19944 18572 19950 18624
rect 22186 18572 22192 18624
rect 22244 18612 22250 18624
rect 22554 18612 22560 18624
rect 22244 18584 22560 18612
rect 22244 18572 22250 18584
rect 22554 18572 22560 18584
rect 22612 18572 22618 18624
rect 552 18522 28428 18544
rect 552 18470 3882 18522
rect 3934 18470 3946 18522
rect 3998 18470 4010 18522
rect 4062 18470 4074 18522
rect 4126 18470 4138 18522
rect 4190 18470 10851 18522
rect 10903 18470 10915 18522
rect 10967 18470 10979 18522
rect 11031 18470 11043 18522
rect 11095 18470 11107 18522
rect 11159 18470 17820 18522
rect 17872 18470 17884 18522
rect 17936 18470 17948 18522
rect 18000 18470 18012 18522
rect 18064 18470 18076 18522
rect 18128 18470 24789 18522
rect 24841 18470 24853 18522
rect 24905 18470 24917 18522
rect 24969 18470 24981 18522
rect 25033 18470 25045 18522
rect 25097 18470 28428 18522
rect 552 18448 28428 18470
rect 2961 18411 3019 18417
rect 2961 18377 2973 18411
rect 3007 18408 3019 18411
rect 3602 18408 3608 18420
rect 3007 18380 3608 18408
rect 3007 18377 3019 18380
rect 2961 18371 3019 18377
rect 3602 18368 3608 18380
rect 3660 18368 3666 18420
rect 5902 18408 5908 18420
rect 4356 18380 5908 18408
rect 1578 18164 1584 18216
rect 1636 18164 1642 18216
rect 1848 18207 1906 18213
rect 1848 18173 1860 18207
rect 1894 18204 1906 18207
rect 2130 18204 2136 18216
rect 1894 18176 2136 18204
rect 1894 18173 1906 18176
rect 1848 18167 1906 18173
rect 2130 18164 2136 18176
rect 2188 18164 2194 18216
rect 4356 18213 4384 18380
rect 5902 18368 5908 18380
rect 5960 18368 5966 18420
rect 8662 18368 8668 18420
rect 8720 18408 8726 18420
rect 8720 18380 8984 18408
rect 8720 18368 8726 18380
rect 5353 18343 5411 18349
rect 5353 18309 5365 18343
rect 5399 18309 5411 18343
rect 5353 18303 5411 18309
rect 7285 18343 7343 18349
rect 7285 18309 7297 18343
rect 7331 18340 7343 18343
rect 7331 18312 8800 18340
rect 7331 18309 7343 18312
rect 7285 18303 7343 18309
rect 4430 18232 4436 18284
rect 4488 18232 4494 18284
rect 4614 18232 4620 18284
rect 4672 18272 4678 18284
rect 4893 18275 4951 18281
rect 4893 18272 4905 18275
rect 4672 18244 4905 18272
rect 4672 18232 4678 18244
rect 4893 18241 4905 18244
rect 4939 18241 4951 18275
rect 4893 18235 4951 18241
rect 4341 18207 4399 18213
rect 4341 18173 4353 18207
rect 4387 18173 4399 18207
rect 4341 18167 4399 18173
rect 4985 18207 5043 18213
rect 4985 18173 4997 18207
rect 5031 18204 5043 18207
rect 5074 18204 5080 18216
rect 5031 18176 5080 18204
rect 5031 18173 5043 18176
rect 4985 18167 5043 18173
rect 5074 18164 5080 18176
rect 5132 18164 5138 18216
rect 5368 18204 5396 18303
rect 5905 18275 5963 18281
rect 5905 18241 5917 18275
rect 5951 18272 5963 18275
rect 7126 18275 7184 18281
rect 7126 18272 7138 18275
rect 5951 18244 7138 18272
rect 5951 18241 5963 18244
rect 5905 18235 5963 18241
rect 7126 18241 7138 18244
rect 7172 18241 7184 18275
rect 7929 18275 7987 18281
rect 7929 18272 7941 18275
rect 7126 18235 7184 18241
rect 7576 18244 7941 18272
rect 6270 18204 6276 18216
rect 5368 18176 6276 18204
rect 6270 18164 6276 18176
rect 6328 18164 6334 18216
rect 6546 18164 6552 18216
rect 6604 18204 6610 18216
rect 6641 18207 6699 18213
rect 6641 18204 6653 18207
rect 6604 18176 6653 18204
rect 6604 18164 6610 18176
rect 6641 18173 6653 18176
rect 6687 18173 6699 18207
rect 6641 18167 6699 18173
rect 6917 18207 6975 18213
rect 6917 18173 6929 18207
rect 6963 18204 6975 18207
rect 7006 18204 7012 18216
rect 6963 18176 7012 18204
rect 6963 18173 6975 18176
rect 6917 18167 6975 18173
rect 7006 18164 7012 18176
rect 7064 18164 7070 18216
rect 5810 18136 5816 18148
rect 4724 18108 5816 18136
rect 4724 18077 4752 18108
rect 5810 18096 5816 18108
rect 5868 18136 5874 18148
rect 6181 18139 6239 18145
rect 6181 18136 6193 18139
rect 5868 18108 6193 18136
rect 5868 18096 5874 18108
rect 6181 18105 6193 18108
rect 6227 18105 6239 18139
rect 6181 18099 6239 18105
rect 6457 18139 6515 18145
rect 6457 18105 6469 18139
rect 6503 18136 6515 18139
rect 7576 18136 7604 18244
rect 7929 18241 7941 18244
rect 7975 18272 7987 18275
rect 8386 18272 8392 18284
rect 7975 18244 8392 18272
rect 7975 18241 7987 18244
rect 7929 18235 7987 18241
rect 8386 18232 8392 18244
rect 8444 18232 8450 18284
rect 8772 18281 8800 18312
rect 8956 18281 8984 18380
rect 9030 18368 9036 18420
rect 9088 18368 9094 18420
rect 11514 18368 11520 18420
rect 11572 18408 11578 18420
rect 12069 18411 12127 18417
rect 12069 18408 12081 18411
rect 11572 18380 12081 18408
rect 11572 18368 11578 18380
rect 12069 18377 12081 18380
rect 12115 18377 12127 18411
rect 12069 18371 12127 18377
rect 8757 18275 8815 18281
rect 8757 18241 8769 18275
rect 8803 18241 8815 18275
rect 8757 18235 8815 18241
rect 8941 18275 8999 18281
rect 8941 18241 8953 18275
rect 8987 18241 8999 18275
rect 9048 18272 9076 18368
rect 12084 18272 12112 18371
rect 12158 18368 12164 18420
rect 12216 18408 12222 18420
rect 12253 18411 12311 18417
rect 12253 18408 12265 18411
rect 12216 18380 12265 18408
rect 12216 18368 12222 18380
rect 12253 18377 12265 18380
rect 12299 18377 12311 18411
rect 12253 18371 12311 18377
rect 13170 18368 13176 18420
rect 13228 18417 13234 18420
rect 13228 18411 13253 18417
rect 13241 18377 13253 18411
rect 13228 18371 13253 18377
rect 13228 18368 13234 18371
rect 13354 18368 13360 18420
rect 13412 18368 13418 18420
rect 13906 18368 13912 18420
rect 13964 18408 13970 18420
rect 14829 18411 14887 18417
rect 14829 18408 14841 18411
rect 13964 18380 14841 18408
rect 13964 18368 13970 18380
rect 14829 18377 14841 18380
rect 14875 18408 14887 18411
rect 17405 18411 17463 18417
rect 14875 18380 16804 18408
rect 14875 18377 14887 18380
rect 14829 18371 14887 18377
rect 16776 18284 16804 18380
rect 17405 18377 17417 18411
rect 17451 18408 17463 18411
rect 17586 18408 17592 18420
rect 17451 18380 17592 18408
rect 17451 18377 17463 18380
rect 17405 18371 17463 18377
rect 17586 18368 17592 18380
rect 17644 18368 17650 18420
rect 19886 18368 19892 18420
rect 19944 18368 19950 18420
rect 16853 18343 16911 18349
rect 16853 18309 16865 18343
rect 16899 18340 16911 18343
rect 17494 18340 17500 18352
rect 16899 18312 17500 18340
rect 16899 18309 16911 18312
rect 16853 18303 16911 18309
rect 17494 18300 17500 18312
rect 17552 18300 17558 18352
rect 13998 18272 14004 18284
rect 9048 18244 9352 18272
rect 12084 18244 14004 18272
rect 8941 18235 8999 18241
rect 7837 18207 7895 18213
rect 7837 18173 7849 18207
rect 7883 18204 7895 18207
rect 7883 18176 8708 18204
rect 7883 18173 7895 18176
rect 7837 18167 7895 18173
rect 6503 18108 7604 18136
rect 8680 18136 8708 18176
rect 8846 18164 8852 18216
rect 8904 18164 8910 18216
rect 9324 18213 9352 18244
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 16758 18232 16764 18284
rect 16816 18232 16822 18284
rect 17052 18244 17540 18272
rect 17052 18216 17080 18244
rect 9033 18207 9091 18213
rect 9033 18173 9045 18207
rect 9079 18173 9091 18207
rect 9033 18167 9091 18173
rect 9309 18207 9367 18213
rect 9309 18173 9321 18207
rect 9355 18173 9367 18207
rect 9309 18167 9367 18173
rect 9048 18136 9076 18167
rect 9582 18164 9588 18216
rect 9640 18164 9646 18216
rect 9674 18164 9680 18216
rect 9732 18164 9738 18216
rect 11701 18207 11759 18213
rect 11701 18173 11713 18207
rect 11747 18204 11759 18207
rect 12434 18204 12440 18216
rect 11747 18176 12440 18204
rect 11747 18173 11759 18176
rect 11701 18167 11759 18173
rect 12434 18164 12440 18176
rect 12492 18204 12498 18216
rect 13541 18207 13599 18213
rect 12492 18176 13124 18204
rect 12492 18164 12498 18176
rect 9493 18139 9551 18145
rect 9493 18136 9505 18139
rect 8680 18108 9076 18136
rect 9232 18108 9505 18136
rect 6503 18105 6515 18108
rect 6457 18099 6515 18105
rect 8956 18080 8984 18108
rect 4709 18071 4767 18077
rect 4709 18037 4721 18071
rect 4755 18037 4767 18071
rect 4709 18031 4767 18037
rect 5994 18028 6000 18080
rect 6052 18068 6058 18080
rect 6089 18071 6147 18077
rect 6089 18068 6101 18071
rect 6052 18040 6101 18068
rect 6052 18028 6058 18040
rect 6089 18037 6101 18040
rect 6135 18037 6147 18071
rect 6089 18031 6147 18037
rect 7006 18028 7012 18080
rect 7064 18028 7070 18080
rect 8205 18071 8263 18077
rect 8205 18037 8217 18071
rect 8251 18068 8263 18071
rect 8478 18068 8484 18080
rect 8251 18040 8484 18068
rect 8251 18037 8263 18040
rect 8205 18031 8263 18037
rect 8478 18028 8484 18040
rect 8536 18028 8542 18080
rect 8938 18028 8944 18080
rect 8996 18028 9002 18080
rect 9232 18077 9260 18108
rect 9493 18105 9505 18108
rect 9539 18105 9551 18139
rect 9493 18099 9551 18105
rect 12529 18139 12587 18145
rect 12529 18105 12541 18139
rect 12575 18136 12587 18139
rect 12618 18136 12624 18148
rect 12575 18108 12624 18136
rect 12575 18105 12587 18108
rect 12529 18099 12587 18105
rect 12618 18096 12624 18108
rect 12676 18096 12682 18148
rect 12710 18096 12716 18148
rect 12768 18096 12774 18148
rect 12894 18096 12900 18148
rect 12952 18136 12958 18148
rect 12989 18139 13047 18145
rect 12989 18136 13001 18139
rect 12952 18108 13001 18136
rect 12952 18096 12958 18108
rect 12989 18105 13001 18108
rect 13035 18105 13047 18139
rect 13096 18136 13124 18176
rect 13541 18173 13553 18207
rect 13587 18204 13599 18207
rect 13722 18204 13728 18216
rect 13587 18176 13728 18204
rect 13587 18173 13599 18176
rect 13541 18167 13599 18173
rect 13722 18164 13728 18176
rect 13780 18164 13786 18216
rect 17034 18164 17040 18216
rect 17092 18164 17098 18216
rect 17512 18213 17540 18244
rect 17221 18207 17279 18213
rect 17221 18173 17233 18207
rect 17267 18204 17279 18207
rect 17313 18207 17371 18213
rect 17313 18204 17325 18207
rect 17267 18176 17325 18204
rect 17267 18173 17279 18176
rect 17221 18167 17279 18173
rect 17313 18173 17325 18176
rect 17359 18173 17371 18207
rect 17313 18167 17371 18173
rect 17497 18207 17555 18213
rect 17497 18173 17509 18207
rect 17543 18173 17555 18207
rect 17497 18167 17555 18173
rect 13189 18139 13247 18145
rect 13189 18136 13201 18139
rect 13096 18108 13201 18136
rect 12989 18099 13047 18105
rect 13189 18105 13201 18108
rect 13235 18105 13247 18139
rect 13189 18099 13247 18105
rect 9217 18071 9275 18077
rect 9217 18037 9229 18071
rect 9263 18037 9275 18071
rect 9217 18031 9275 18037
rect 9858 18028 9864 18080
rect 9916 18028 9922 18080
rect 12069 18071 12127 18077
rect 12069 18037 12081 18071
rect 12115 18068 12127 18071
rect 12345 18071 12403 18077
rect 12345 18068 12357 18071
rect 12115 18040 12357 18068
rect 12115 18037 12127 18040
rect 12069 18031 12127 18037
rect 12345 18037 12357 18040
rect 12391 18037 12403 18071
rect 13004 18068 13032 18099
rect 16482 18096 16488 18148
rect 16540 18145 16546 18148
rect 16540 18099 16552 18145
rect 17328 18136 17356 18167
rect 18138 18164 18144 18216
rect 18196 18204 18202 18216
rect 19521 18207 19579 18213
rect 19521 18204 19533 18207
rect 18196 18176 19533 18204
rect 18196 18164 18202 18176
rect 19521 18173 19533 18176
rect 19567 18173 19579 18207
rect 19521 18167 19579 18173
rect 19705 18207 19763 18213
rect 19705 18173 19717 18207
rect 19751 18204 19763 18207
rect 19904 18204 19932 18368
rect 19751 18176 19932 18204
rect 19751 18173 19763 18176
rect 19705 18167 19763 18173
rect 18322 18136 18328 18148
rect 17328 18108 18328 18136
rect 16540 18096 16546 18099
rect 18322 18096 18328 18108
rect 18380 18096 18386 18148
rect 14826 18068 14832 18080
rect 13004 18040 14832 18068
rect 12345 18031 12403 18037
rect 14826 18028 14832 18040
rect 14884 18068 14890 18080
rect 15378 18068 15384 18080
rect 14884 18040 15384 18068
rect 14884 18028 14890 18040
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 19610 18028 19616 18080
rect 19668 18028 19674 18080
rect 552 17978 28587 18000
rect 552 17926 7366 17978
rect 7418 17926 7430 17978
rect 7482 17926 7494 17978
rect 7546 17926 7558 17978
rect 7610 17926 7622 17978
rect 7674 17926 14335 17978
rect 14387 17926 14399 17978
rect 14451 17926 14463 17978
rect 14515 17926 14527 17978
rect 14579 17926 14591 17978
rect 14643 17926 21304 17978
rect 21356 17926 21368 17978
rect 21420 17926 21432 17978
rect 21484 17926 21496 17978
rect 21548 17926 21560 17978
rect 21612 17926 28273 17978
rect 28325 17926 28337 17978
rect 28389 17926 28401 17978
rect 28453 17926 28465 17978
rect 28517 17926 28529 17978
rect 28581 17926 28587 17978
rect 552 17904 28587 17926
rect 7006 17824 7012 17876
rect 7064 17864 7070 17876
rect 7193 17867 7251 17873
rect 7193 17864 7205 17867
rect 7064 17836 7205 17864
rect 7064 17824 7070 17836
rect 7193 17833 7205 17836
rect 7239 17833 7251 17867
rect 7193 17827 7251 17833
rect 8941 17867 8999 17873
rect 8941 17833 8953 17867
rect 8987 17864 8999 17867
rect 9674 17864 9680 17876
rect 8987 17836 9680 17864
rect 8987 17833 8999 17836
rect 8941 17827 8999 17833
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 10965 17867 11023 17873
rect 10965 17833 10977 17867
rect 11011 17833 11023 17867
rect 10965 17827 11023 17833
rect 10536 17799 10594 17805
rect 10536 17765 10548 17799
rect 10582 17796 10594 17799
rect 10980 17796 11008 17827
rect 13354 17824 13360 17876
rect 13412 17864 13418 17876
rect 13722 17864 13728 17876
rect 13412 17836 13728 17864
rect 13412 17824 13418 17836
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 14093 17867 14151 17873
rect 14093 17833 14105 17867
rect 14139 17864 14151 17867
rect 14369 17867 14427 17873
rect 14369 17864 14381 17867
rect 14139 17836 14381 17864
rect 14139 17833 14151 17836
rect 14093 17827 14151 17833
rect 14369 17833 14381 17836
rect 14415 17833 14427 17867
rect 18690 17864 18696 17876
rect 14369 17827 14427 17833
rect 14752 17836 18696 17864
rect 10582 17768 11008 17796
rect 10582 17765 10594 17768
rect 10536 17759 10594 17765
rect 13262 17756 13268 17808
rect 13320 17796 13326 17808
rect 14752 17796 14780 17836
rect 13320 17768 14780 17796
rect 13320 17756 13326 17768
rect 3228 17731 3286 17737
rect 3228 17697 3240 17731
rect 3274 17728 3286 17731
rect 3694 17728 3700 17740
rect 3274 17700 3700 17728
rect 3274 17697 3286 17700
rect 3228 17691 3286 17697
rect 3694 17688 3700 17700
rect 3752 17688 3758 17740
rect 5810 17688 5816 17740
rect 5868 17728 5874 17740
rect 5905 17731 5963 17737
rect 5905 17728 5917 17731
rect 5868 17700 5917 17728
rect 5868 17688 5874 17700
rect 5905 17697 5917 17700
rect 5951 17697 5963 17731
rect 5905 17691 5963 17697
rect 5997 17731 6055 17737
rect 5997 17697 6009 17731
rect 6043 17728 6055 17731
rect 6086 17728 6092 17740
rect 6043 17700 6092 17728
rect 6043 17697 6055 17700
rect 5997 17691 6055 17697
rect 6086 17688 6092 17700
rect 6144 17688 6150 17740
rect 6365 17731 6423 17737
rect 6365 17697 6377 17731
rect 6411 17728 6423 17731
rect 6546 17728 6552 17740
rect 6411 17700 6552 17728
rect 6411 17697 6423 17700
rect 6365 17691 6423 17697
rect 6546 17688 6552 17700
rect 6604 17688 6610 17740
rect 7282 17688 7288 17740
rect 7340 17688 7346 17740
rect 8294 17688 8300 17740
rect 8352 17688 8358 17740
rect 8478 17688 8484 17740
rect 8536 17728 8542 17740
rect 8757 17731 8815 17737
rect 8757 17728 8769 17731
rect 8536 17700 8769 17728
rect 8536 17688 8542 17700
rect 8757 17697 8769 17700
rect 8803 17697 8815 17731
rect 8757 17691 8815 17697
rect 10042 17688 10048 17740
rect 10100 17728 10106 17740
rect 11149 17731 11207 17737
rect 11149 17728 11161 17731
rect 10100 17700 11161 17728
rect 10100 17688 10106 17700
rect 11149 17697 11161 17700
rect 11195 17697 11207 17731
rect 11149 17691 11207 17697
rect 11701 17731 11759 17737
rect 11701 17697 11713 17731
rect 11747 17697 11759 17731
rect 11701 17691 11759 17697
rect 11977 17731 12035 17737
rect 11977 17697 11989 17731
rect 12023 17697 12035 17731
rect 11977 17691 12035 17697
rect 12161 17731 12219 17737
rect 12161 17697 12173 17731
rect 12207 17728 12219 17731
rect 12345 17731 12403 17737
rect 12345 17728 12357 17731
rect 12207 17700 12357 17728
rect 12207 17697 12219 17700
rect 12161 17691 12219 17697
rect 12345 17697 12357 17700
rect 12391 17697 12403 17731
rect 12345 17691 12403 17697
rect 1578 17620 1584 17672
rect 1636 17660 1642 17672
rect 2961 17663 3019 17669
rect 2961 17660 2973 17663
rect 1636 17632 2973 17660
rect 1636 17620 1642 17632
rect 2961 17629 2973 17632
rect 3007 17629 3019 17663
rect 2961 17623 3019 17629
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17629 8631 17663
rect 8573 17623 8631 17629
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17660 10839 17663
rect 11238 17660 11244 17672
rect 10827 17632 11244 17660
rect 10827 17629 10839 17632
rect 10781 17623 10839 17629
rect 6549 17595 6607 17601
rect 6549 17561 6561 17595
rect 6595 17592 6607 17595
rect 8588 17592 8616 17623
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 6595 17564 8616 17592
rect 6595 17561 6607 17564
rect 6549 17555 6607 17561
rect 8846 17552 8852 17604
rect 8904 17592 8910 17604
rect 9401 17595 9459 17601
rect 9401 17592 9413 17595
rect 8904 17564 9413 17592
rect 8904 17552 8910 17564
rect 9401 17561 9413 17564
rect 9447 17592 9459 17595
rect 9582 17592 9588 17604
rect 9447 17564 9588 17592
rect 9447 17561 9459 17564
rect 9401 17555 9459 17561
rect 9582 17552 9588 17564
rect 9640 17552 9646 17604
rect 11716 17592 11744 17691
rect 11992 17660 12020 17691
rect 12618 17688 12624 17740
rect 12676 17728 12682 17740
rect 13354 17728 13360 17740
rect 12676 17700 13360 17728
rect 12676 17688 12682 17700
rect 13354 17688 13360 17700
rect 13412 17688 13418 17740
rect 13449 17731 13507 17737
rect 13449 17697 13461 17731
rect 13495 17728 13507 17731
rect 13495 17700 13676 17728
rect 13495 17697 13507 17700
rect 13449 17691 13507 17697
rect 13648 17672 13676 17700
rect 13722 17688 13728 17740
rect 13780 17688 13786 17740
rect 14737 17732 14795 17737
rect 14660 17731 14795 17732
rect 14660 17728 14749 17731
rect 13832 17704 14749 17728
rect 13832 17700 14688 17704
rect 12434 17660 12440 17672
rect 11992 17632 12440 17660
rect 12434 17620 12440 17632
rect 12492 17620 12498 17672
rect 12989 17663 13047 17669
rect 12989 17629 13001 17663
rect 13035 17660 13047 17663
rect 13170 17660 13176 17672
rect 13035 17632 13176 17660
rect 13035 17629 13047 17632
rect 12989 17623 13047 17629
rect 13170 17620 13176 17632
rect 13228 17620 13234 17672
rect 13265 17663 13323 17669
rect 13265 17629 13277 17663
rect 13311 17660 13323 17663
rect 13311 17632 13400 17660
rect 13311 17629 13323 17632
rect 13265 17623 13323 17629
rect 13081 17595 13139 17601
rect 13081 17592 13093 17595
rect 11716 17564 13093 17592
rect 13081 17561 13093 17564
rect 13127 17561 13139 17595
rect 13081 17555 13139 17561
rect 4341 17527 4399 17533
rect 4341 17493 4353 17527
rect 4387 17524 4399 17527
rect 4614 17524 4620 17536
rect 4387 17496 4620 17524
rect 4387 17493 4399 17496
rect 4341 17487 4399 17493
rect 4614 17484 4620 17496
rect 4672 17484 4678 17536
rect 6270 17484 6276 17536
rect 6328 17484 6334 17536
rect 8754 17484 8760 17536
rect 8812 17484 8818 17536
rect 11514 17484 11520 17536
rect 11572 17484 11578 17536
rect 12710 17484 12716 17536
rect 12768 17524 12774 17536
rect 13372 17524 13400 17632
rect 13538 17620 13544 17672
rect 13596 17620 13602 17672
rect 13630 17620 13636 17672
rect 13688 17660 13694 17672
rect 13832 17660 13860 17700
rect 14737 17697 14749 17704
rect 14783 17697 14795 17731
rect 14737 17691 14795 17697
rect 13688 17632 13860 17660
rect 13688 17620 13694 17632
rect 14550 17620 14556 17672
rect 14608 17620 14614 17672
rect 14642 17620 14648 17672
rect 14700 17620 14706 17672
rect 14752 17660 14780 17691
rect 14826 17688 14832 17740
rect 14884 17688 14890 17740
rect 15010 17688 15016 17740
rect 15068 17688 15074 17740
rect 15102 17688 15108 17740
rect 15160 17728 15166 17740
rect 16117 17731 16175 17737
rect 16117 17728 16129 17731
rect 15160 17700 16129 17728
rect 15160 17688 15166 17700
rect 16117 17697 16129 17700
rect 16163 17697 16175 17731
rect 16500 17728 16528 17836
rect 18690 17824 18696 17836
rect 18748 17864 18754 17876
rect 19061 17867 19119 17873
rect 19061 17864 19073 17867
rect 18748 17836 19073 17864
rect 18748 17824 18754 17836
rect 19061 17833 19073 17836
rect 19107 17833 19119 17867
rect 19061 17827 19119 17833
rect 19610 17824 19616 17876
rect 19668 17864 19674 17876
rect 19668 17836 19748 17864
rect 19668 17824 19674 17836
rect 19720 17796 19748 17836
rect 20714 17824 20720 17876
rect 20772 17864 20778 17876
rect 20993 17867 21051 17873
rect 20993 17864 21005 17867
rect 20772 17836 21005 17864
rect 20772 17824 20778 17836
rect 20993 17833 21005 17836
rect 21039 17833 21051 17867
rect 20993 17827 21051 17833
rect 19858 17799 19916 17805
rect 19858 17796 19870 17799
rect 17696 17768 19656 17796
rect 19720 17768 19870 17796
rect 17696 17740 17724 17768
rect 16669 17731 16727 17737
rect 16669 17728 16681 17731
rect 16500 17700 16681 17728
rect 16117 17691 16175 17697
rect 16669 17697 16681 17700
rect 16715 17697 16727 17731
rect 16669 17691 16727 17697
rect 16758 17688 16764 17740
rect 16816 17728 16822 17740
rect 17678 17728 17684 17740
rect 16816 17700 17684 17728
rect 16816 17688 16822 17700
rect 17678 17688 17684 17700
rect 17736 17688 17742 17740
rect 19628 17737 19656 17768
rect 19858 17765 19870 17768
rect 19904 17765 19916 17799
rect 19858 17759 19916 17765
rect 17937 17731 17995 17737
rect 17937 17728 17949 17731
rect 17788 17700 17949 17728
rect 15654 17660 15660 17672
rect 14752 17632 15660 17660
rect 15654 17620 15660 17632
rect 15712 17620 15718 17672
rect 16482 17620 16488 17672
rect 16540 17620 16546 17672
rect 17034 17620 17040 17672
rect 17092 17660 17098 17672
rect 17788 17660 17816 17700
rect 17937 17697 17949 17700
rect 17983 17697 17995 17731
rect 17937 17691 17995 17697
rect 19613 17731 19671 17737
rect 19613 17697 19625 17731
rect 19659 17697 19671 17731
rect 19613 17691 19671 17697
rect 17092 17632 17816 17660
rect 17092 17620 17098 17632
rect 14277 17595 14335 17601
rect 13832 17564 14228 17592
rect 13832 17524 13860 17564
rect 12768 17496 13860 17524
rect 12768 17484 12774 17496
rect 13998 17484 14004 17536
rect 14056 17524 14062 17536
rect 14093 17527 14151 17533
rect 14093 17524 14105 17527
rect 14056 17496 14105 17524
rect 14056 17484 14062 17496
rect 14093 17493 14105 17496
rect 14139 17493 14151 17527
rect 14200 17524 14228 17564
rect 14277 17561 14289 17595
rect 14323 17592 14335 17595
rect 14458 17592 14464 17604
rect 14323 17564 14464 17592
rect 14323 17561 14335 17564
rect 14277 17555 14335 17561
rect 14458 17552 14464 17564
rect 14516 17552 14522 17604
rect 15197 17595 15255 17601
rect 15197 17561 15209 17595
rect 15243 17592 15255 17595
rect 16500 17592 16528 17620
rect 15243 17564 16528 17592
rect 15243 17561 15255 17564
rect 15197 17555 15255 17561
rect 14550 17524 14556 17536
rect 14200 17496 14556 17524
rect 14093 17487 14151 17493
rect 14550 17484 14556 17496
rect 14608 17484 14614 17536
rect 14642 17484 14648 17536
rect 14700 17524 14706 17536
rect 16942 17524 16948 17536
rect 14700 17496 16948 17524
rect 14700 17484 14706 17496
rect 16942 17484 16948 17496
rect 17000 17484 17006 17536
rect 552 17434 28428 17456
rect 552 17382 3882 17434
rect 3934 17382 3946 17434
rect 3998 17382 4010 17434
rect 4062 17382 4074 17434
rect 4126 17382 4138 17434
rect 4190 17382 10851 17434
rect 10903 17382 10915 17434
rect 10967 17382 10979 17434
rect 11031 17382 11043 17434
rect 11095 17382 11107 17434
rect 11159 17382 17820 17434
rect 17872 17382 17884 17434
rect 17936 17382 17948 17434
rect 18000 17382 18012 17434
rect 18064 17382 18076 17434
rect 18128 17382 24789 17434
rect 24841 17382 24853 17434
rect 24905 17382 24917 17434
rect 24969 17382 24981 17434
rect 25033 17382 25045 17434
rect 25097 17382 28428 17434
rect 552 17360 28428 17382
rect 3694 17280 3700 17332
rect 3752 17280 3758 17332
rect 8938 17280 8944 17332
rect 8996 17280 9002 17332
rect 9858 17280 9864 17332
rect 9916 17280 9922 17332
rect 10042 17280 10048 17332
rect 10100 17280 10106 17332
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 12529 17323 12587 17329
rect 12529 17320 12541 17323
rect 12492 17292 12541 17320
rect 12492 17280 12498 17292
rect 12529 17289 12541 17292
rect 12575 17289 12587 17323
rect 12529 17283 12587 17289
rect 12894 17280 12900 17332
rect 12952 17320 12958 17332
rect 13173 17323 13231 17329
rect 13173 17320 13185 17323
rect 12952 17292 13185 17320
rect 12952 17280 12958 17292
rect 13173 17289 13185 17292
rect 13219 17289 13231 17323
rect 13173 17283 13231 17289
rect 13357 17323 13415 17329
rect 13357 17289 13369 17323
rect 13403 17320 13415 17323
rect 13446 17320 13452 17332
rect 13403 17292 13452 17320
rect 13403 17289 13415 17292
rect 13357 17283 13415 17289
rect 13188 17252 13216 17283
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 13998 17280 14004 17332
rect 14056 17320 14062 17332
rect 15286 17320 15292 17332
rect 14056 17292 15292 17320
rect 14056 17280 14062 17292
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 16117 17323 16175 17329
rect 16117 17289 16129 17323
rect 16163 17289 16175 17323
rect 16117 17283 16175 17289
rect 16132 17252 16160 17283
rect 17034 17280 17040 17332
rect 17092 17280 17098 17332
rect 19334 17252 19340 17264
rect 13188 17224 13952 17252
rect 16132 17224 16804 17252
rect 12897 17187 12955 17193
rect 12897 17153 12909 17187
rect 12943 17184 12955 17187
rect 13354 17184 13360 17196
rect 12943 17156 13360 17184
rect 12943 17153 12955 17156
rect 12897 17147 12955 17153
rect 13354 17144 13360 17156
rect 13412 17144 13418 17196
rect 3326 17076 3332 17128
rect 3384 17076 3390 17128
rect 3418 17076 3424 17128
rect 3476 17076 3482 17128
rect 3605 17119 3663 17125
rect 3605 17085 3617 17119
rect 3651 17116 3663 17119
rect 3881 17119 3939 17125
rect 3881 17116 3893 17119
rect 3651 17088 3893 17116
rect 3651 17085 3663 17088
rect 3605 17079 3663 17085
rect 3881 17085 3893 17088
rect 3927 17085 3939 17119
rect 3881 17079 3939 17085
rect 12710 17076 12716 17128
rect 12768 17076 12774 17128
rect 13924 17116 13952 17224
rect 14093 17187 14151 17193
rect 14093 17153 14105 17187
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 14369 17187 14427 17193
rect 14369 17153 14381 17187
rect 14415 17153 14427 17187
rect 14369 17147 14427 17153
rect 15289 17187 15347 17193
rect 15289 17153 15301 17187
rect 15335 17184 15347 17187
rect 16577 17187 16635 17193
rect 16577 17184 16589 17187
rect 15335 17156 15608 17184
rect 15335 17153 15347 17156
rect 15289 17147 15347 17153
rect 14001 17119 14059 17125
rect 14001 17116 14013 17119
rect 13924 17088 14013 17116
rect 14001 17085 14013 17088
rect 14047 17085 14059 17119
rect 14001 17079 14059 17085
rect 6730 17008 6736 17060
rect 6788 17048 6794 17060
rect 8389 17051 8447 17057
rect 8389 17048 8401 17051
rect 6788 17020 8401 17048
rect 6788 17008 6794 17020
rect 8389 17017 8401 17020
rect 8435 17017 8447 17051
rect 8389 17011 8447 17017
rect 9677 17051 9735 17057
rect 9677 17017 9689 17051
rect 9723 17048 9735 17051
rect 10410 17048 10416 17060
rect 9723 17020 10416 17048
rect 9723 17017 9735 17020
rect 9677 17011 9735 17017
rect 10410 17008 10416 17020
rect 10468 17008 10474 17060
rect 12989 17051 13047 17057
rect 12989 17017 13001 17051
rect 13035 17048 13047 17051
rect 13035 17020 14044 17048
rect 13035 17017 13047 17020
rect 12989 17011 13047 17017
rect 14016 16992 14044 17020
rect 6546 16940 6552 16992
rect 6604 16980 6610 16992
rect 8570 16980 8576 16992
rect 6604 16952 8576 16980
rect 6604 16940 6610 16952
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 8662 16940 8668 16992
rect 8720 16940 8726 16992
rect 8757 16983 8815 16989
rect 8757 16949 8769 16983
rect 8803 16980 8815 16983
rect 8938 16980 8944 16992
rect 8803 16952 8944 16980
rect 8803 16949 8815 16952
rect 8757 16943 8815 16949
rect 8938 16940 8944 16952
rect 8996 16940 9002 16992
rect 9766 16940 9772 16992
rect 9824 16980 9830 16992
rect 9877 16983 9935 16989
rect 9877 16980 9889 16983
rect 9824 16952 9889 16980
rect 9824 16940 9830 16952
rect 9877 16949 9889 16952
rect 9923 16949 9935 16983
rect 9877 16943 9935 16949
rect 12526 16940 12532 16992
rect 12584 16980 12590 16992
rect 13170 16980 13176 16992
rect 13228 16989 13234 16992
rect 13228 16983 13257 16989
rect 12584 16952 13176 16980
rect 12584 16940 12590 16952
rect 13170 16940 13176 16952
rect 13245 16980 13257 16983
rect 13630 16980 13636 16992
rect 13245 16952 13636 16980
rect 13245 16949 13257 16952
rect 13228 16943 13257 16949
rect 13228 16940 13234 16943
rect 13630 16940 13636 16952
rect 13688 16940 13694 16992
rect 13998 16940 14004 16992
rect 14056 16940 14062 16992
rect 14108 16980 14136 17147
rect 14384 17048 14412 17147
rect 15194 17076 15200 17128
rect 15252 17076 15258 17128
rect 15381 17119 15439 17125
rect 15381 17085 15393 17119
rect 15427 17085 15439 17119
rect 15381 17079 15439 17085
rect 15396 17048 15424 17079
rect 15470 17076 15476 17128
rect 15528 17076 15534 17128
rect 15580 17125 15608 17156
rect 15764 17156 16589 17184
rect 15764 17125 15792 17156
rect 16577 17153 16589 17156
rect 16623 17153 16635 17187
rect 16577 17147 16635 17153
rect 16666 17144 16672 17196
rect 16724 17144 16730 17196
rect 15566 17119 15624 17125
rect 15566 17085 15578 17119
rect 15612 17085 15624 17119
rect 15566 17079 15624 17085
rect 15749 17119 15807 17125
rect 15749 17085 15761 17119
rect 15795 17085 15807 17119
rect 15749 17079 15807 17085
rect 15930 17076 15936 17128
rect 15988 17125 15994 17128
rect 15988 17116 15996 17125
rect 15988 17088 16033 17116
rect 15988 17079 15996 17088
rect 15988 17076 15994 17079
rect 14384 17020 15424 17048
rect 15010 16980 15016 16992
rect 14108 16952 15016 16980
rect 15010 16940 15016 16952
rect 15068 16940 15074 16992
rect 15396 16980 15424 17020
rect 15838 17008 15844 17060
rect 15896 17008 15902 17060
rect 16206 17008 16212 17060
rect 16264 17008 16270 17060
rect 16390 17048 16396 17060
rect 16316 17020 16396 17048
rect 16316 16980 16344 17020
rect 16390 17008 16396 17020
rect 16448 17008 16454 17060
rect 16684 17048 16712 17144
rect 16776 17116 16804 17224
rect 17512 17224 19340 17252
rect 16850 17144 16856 17196
rect 16908 17184 16914 17196
rect 17512 17184 17540 17224
rect 19334 17212 19340 17224
rect 19392 17252 19398 17264
rect 23290 17252 23296 17264
rect 19392 17224 23296 17252
rect 19392 17212 19398 17224
rect 23290 17212 23296 17224
rect 23348 17212 23354 17264
rect 17773 17187 17831 17193
rect 17773 17184 17785 17187
rect 16908 17156 17540 17184
rect 16908 17144 16914 17156
rect 17313 17119 17371 17125
rect 17313 17116 17325 17119
rect 16776 17088 17325 17116
rect 17313 17085 17325 17088
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 17402 17076 17408 17128
rect 17460 17076 17466 17128
rect 17512 17125 17540 17156
rect 17696 17156 17785 17184
rect 17696 17125 17724 17156
rect 17773 17153 17785 17156
rect 17819 17153 17831 17187
rect 18138 17184 18144 17196
rect 17773 17147 17831 17153
rect 17880 17156 18144 17184
rect 17497 17119 17555 17125
rect 17497 17085 17509 17119
rect 17543 17085 17555 17119
rect 17497 17079 17555 17085
rect 17681 17119 17739 17125
rect 17681 17085 17693 17119
rect 17727 17085 17739 17119
rect 17681 17079 17739 17085
rect 17880 17048 17908 17156
rect 18138 17144 18144 17156
rect 18196 17144 18202 17196
rect 18233 17187 18291 17193
rect 18233 17153 18245 17187
rect 18279 17184 18291 17187
rect 18690 17184 18696 17196
rect 18279 17156 18696 17184
rect 18279 17153 18291 17156
rect 18233 17147 18291 17153
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 18966 17144 18972 17196
rect 19024 17144 19030 17196
rect 17954 17076 17960 17128
rect 18012 17076 18018 17128
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17085 18107 17119
rect 18049 17079 18107 17085
rect 16684 17020 17908 17048
rect 15396 16952 16344 16980
rect 17494 16940 17500 16992
rect 17552 16980 17558 16992
rect 18064 16980 18092 17079
rect 18598 17076 18604 17128
rect 18656 17116 18662 17128
rect 19061 17119 19119 17125
rect 19061 17116 19073 17119
rect 18656 17088 19073 17116
rect 18656 17076 18662 17088
rect 19061 17085 19073 17088
rect 19107 17085 19119 17119
rect 19061 17079 19119 17085
rect 20346 17076 20352 17128
rect 20404 17076 20410 17128
rect 17552 16952 18092 16980
rect 17552 16940 17558 16952
rect 18598 16940 18604 16992
rect 18656 16980 18662 16992
rect 18693 16983 18751 16989
rect 18693 16980 18705 16983
rect 18656 16952 18705 16980
rect 18656 16940 18662 16952
rect 18693 16949 18705 16952
rect 18739 16949 18751 16983
rect 18693 16943 18751 16949
rect 20162 16940 20168 16992
rect 20220 16980 20226 16992
rect 20441 16983 20499 16989
rect 20441 16980 20453 16983
rect 20220 16952 20453 16980
rect 20220 16940 20226 16952
rect 20441 16949 20453 16952
rect 20487 16949 20499 16983
rect 20441 16943 20499 16949
rect 552 16890 28587 16912
rect 552 16838 7366 16890
rect 7418 16838 7430 16890
rect 7482 16838 7494 16890
rect 7546 16838 7558 16890
rect 7610 16838 7622 16890
rect 7674 16838 14335 16890
rect 14387 16838 14399 16890
rect 14451 16838 14463 16890
rect 14515 16838 14527 16890
rect 14579 16838 14591 16890
rect 14643 16838 21304 16890
rect 21356 16838 21368 16890
rect 21420 16838 21432 16890
rect 21484 16838 21496 16890
rect 21548 16838 21560 16890
rect 21612 16838 28273 16890
rect 28325 16838 28337 16890
rect 28389 16838 28401 16890
rect 28453 16838 28465 16890
rect 28517 16838 28529 16890
rect 28581 16838 28587 16890
rect 552 16816 28587 16838
rect 3418 16736 3424 16788
rect 3476 16776 3482 16788
rect 4157 16779 4215 16785
rect 4157 16776 4169 16779
rect 3476 16748 4169 16776
rect 3476 16736 3482 16748
rect 4157 16745 4169 16748
rect 4203 16745 4215 16779
rect 4157 16739 4215 16745
rect 4798 16736 4804 16788
rect 4856 16776 4862 16788
rect 6822 16776 6828 16788
rect 4856 16748 5304 16776
rect 4856 16736 4862 16748
rect 4433 16711 4491 16717
rect 4433 16677 4445 16711
rect 4479 16708 4491 16711
rect 4614 16708 4620 16720
rect 4479 16680 4620 16708
rect 4479 16677 4491 16680
rect 4433 16671 4491 16677
rect 4614 16668 4620 16680
rect 4672 16708 4678 16720
rect 4672 16680 5212 16708
rect 4672 16668 4678 16680
rect 5184 16652 5212 16680
rect 2130 16600 2136 16652
rect 2188 16600 2194 16652
rect 4341 16643 4399 16649
rect 4341 16609 4353 16643
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 4356 16572 4384 16603
rect 4522 16600 4528 16652
rect 4580 16600 4586 16652
rect 4706 16600 4712 16652
rect 4764 16600 4770 16652
rect 5166 16600 5172 16652
rect 5224 16600 5230 16652
rect 5276 16649 5304 16748
rect 6380 16748 6828 16776
rect 6270 16668 6276 16720
rect 6328 16668 6334 16720
rect 6380 16717 6408 16748
rect 6822 16736 6828 16748
rect 6880 16776 6886 16788
rect 7929 16779 7987 16785
rect 6880 16748 7788 16776
rect 6880 16736 6886 16748
rect 6365 16711 6423 16717
rect 6365 16677 6377 16711
rect 6411 16677 6423 16711
rect 7282 16708 7288 16720
rect 6365 16671 6423 16677
rect 6564 16680 7288 16708
rect 6477 16665 6535 16671
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16609 5319 16643
rect 6089 16643 6147 16649
rect 6089 16640 6101 16643
rect 5261 16603 5319 16609
rect 5552 16612 6101 16640
rect 4356 16544 4752 16572
rect 4724 16448 4752 16544
rect 5276 16504 5304 16603
rect 5350 16532 5356 16584
rect 5408 16532 5414 16584
rect 5552 16504 5580 16612
rect 6089 16609 6101 16612
rect 6135 16640 6147 16643
rect 6178 16640 6184 16652
rect 6135 16612 6184 16640
rect 6135 16609 6147 16612
rect 6089 16603 6147 16609
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 6477 16631 6489 16665
rect 6523 16662 6535 16665
rect 6564 16662 6592 16680
rect 7282 16668 7288 16680
rect 7340 16708 7346 16720
rect 7340 16680 7604 16708
rect 7340 16668 7346 16680
rect 6523 16634 6592 16662
rect 6641 16643 6699 16649
rect 6523 16631 6535 16634
rect 6477 16625 6535 16631
rect 6641 16609 6653 16643
rect 6687 16609 6699 16643
rect 6641 16603 6699 16609
rect 5994 16572 6000 16584
rect 5644 16544 6000 16572
rect 5644 16513 5672 16544
rect 5994 16532 6000 16544
rect 6052 16532 6058 16584
rect 6546 16532 6552 16584
rect 6604 16572 6610 16584
rect 6656 16572 6684 16603
rect 6730 16600 6736 16652
rect 6788 16600 6794 16652
rect 6914 16600 6920 16652
rect 6972 16600 6978 16652
rect 7101 16643 7159 16649
rect 7101 16609 7113 16643
rect 7147 16640 7159 16643
rect 7193 16643 7251 16649
rect 7193 16640 7205 16643
rect 7147 16612 7205 16640
rect 7147 16609 7159 16612
rect 7101 16603 7159 16609
rect 7193 16609 7205 16612
rect 7239 16609 7251 16643
rect 7193 16603 7251 16609
rect 7374 16600 7380 16652
rect 7432 16600 7438 16652
rect 7576 16581 7604 16680
rect 7760 16649 7788 16748
rect 7929 16745 7941 16779
rect 7975 16776 7987 16779
rect 8294 16776 8300 16788
rect 7975 16748 8300 16776
rect 7975 16745 7987 16748
rect 7929 16739 7987 16745
rect 8294 16736 8300 16748
rect 8352 16736 8358 16788
rect 8404 16748 9076 16776
rect 8018 16668 8024 16720
rect 8076 16708 8082 16720
rect 8404 16708 8432 16748
rect 8076 16680 8432 16708
rect 8076 16668 8082 16680
rect 8944 16652 8996 16658
rect 7745 16643 7803 16649
rect 7745 16609 7757 16643
rect 7791 16609 7803 16643
rect 7745 16603 7803 16609
rect 9048 16649 9076 16748
rect 9766 16736 9772 16788
rect 9824 16736 9830 16788
rect 10318 16736 10324 16788
rect 10376 16736 10382 16788
rect 11514 16736 11520 16788
rect 11572 16736 11578 16788
rect 12526 16736 12532 16788
rect 12584 16736 12590 16788
rect 13078 16736 13084 16788
rect 13136 16776 13142 16788
rect 15381 16779 15439 16785
rect 13136 16748 15148 16776
rect 13136 16736 13142 16748
rect 9674 16668 9680 16720
rect 9732 16668 9738 16720
rect 9033 16643 9091 16649
rect 9033 16609 9045 16643
rect 9079 16609 9091 16643
rect 9033 16603 9091 16609
rect 9582 16600 9588 16652
rect 9640 16600 9646 16652
rect 9692 16640 9720 16668
rect 9769 16643 9827 16649
rect 9769 16640 9781 16643
rect 9692 16612 9781 16640
rect 9769 16609 9781 16612
rect 9815 16609 9827 16643
rect 9769 16603 9827 16609
rect 10137 16643 10195 16649
rect 10137 16609 10149 16643
rect 10183 16640 10195 16643
rect 10336 16640 10364 16736
rect 11416 16711 11474 16717
rect 11416 16677 11428 16711
rect 11462 16708 11474 16711
rect 11532 16708 11560 16736
rect 13096 16708 13124 16736
rect 11462 16680 11560 16708
rect 12820 16680 13124 16708
rect 11462 16677 11474 16680
rect 11416 16671 11474 16677
rect 10183 16612 10364 16640
rect 11149 16643 11207 16649
rect 10183 16609 10195 16612
rect 10137 16603 10195 16609
rect 11149 16609 11161 16643
rect 11195 16640 11207 16643
rect 11238 16640 11244 16652
rect 11195 16612 11244 16640
rect 11195 16609 11207 16612
rect 11149 16603 11207 16609
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 12820 16649 12848 16680
rect 14918 16668 14924 16720
rect 14976 16668 14982 16720
rect 15010 16668 15016 16720
rect 15068 16668 15074 16720
rect 12805 16643 12863 16649
rect 12805 16609 12817 16643
rect 12851 16609 12863 16643
rect 14936 16640 14964 16668
rect 12805 16603 12863 16609
rect 13096 16612 14964 16640
rect 15120 16638 15148 16748
rect 15381 16745 15393 16779
rect 15427 16776 15439 16779
rect 15470 16776 15476 16788
rect 15427 16748 15476 16776
rect 15427 16745 15439 16748
rect 15381 16739 15439 16745
rect 15470 16736 15476 16748
rect 15528 16736 15534 16788
rect 17494 16736 17500 16788
rect 17552 16736 17558 16788
rect 17589 16779 17647 16785
rect 17589 16745 17601 16779
rect 17635 16776 17647 16779
rect 17954 16776 17960 16788
rect 17635 16748 17960 16776
rect 17635 16745 17647 16748
rect 17589 16739 17647 16745
rect 17954 16736 17960 16748
rect 18012 16736 18018 16788
rect 18690 16736 18696 16788
rect 18748 16776 18754 16788
rect 18748 16748 18828 16776
rect 18748 16736 18754 16748
rect 15194 16668 15200 16720
rect 15252 16717 15258 16720
rect 15252 16711 15287 16717
rect 15275 16708 15287 16711
rect 15562 16708 15568 16720
rect 15275 16680 15568 16708
rect 15275 16677 15287 16680
rect 15252 16671 15287 16677
rect 15252 16668 15258 16671
rect 15562 16668 15568 16680
rect 15620 16708 15626 16720
rect 16206 16708 16212 16720
rect 15620 16680 16212 16708
rect 15620 16668 15626 16680
rect 16206 16668 16212 16680
rect 16264 16668 16270 16720
rect 16574 16668 16580 16720
rect 16632 16708 16638 16720
rect 18800 16717 18828 16748
rect 17773 16711 17831 16717
rect 17773 16708 17785 16711
rect 16632 16680 17785 16708
rect 16632 16668 16638 16680
rect 17773 16677 17785 16680
rect 17819 16677 17831 16711
rect 17773 16671 17831 16677
rect 18585 16711 18643 16717
rect 18585 16677 18597 16711
rect 18631 16708 18643 16711
rect 18785 16711 18843 16717
rect 18631 16680 18736 16708
rect 18631 16677 18643 16680
rect 18585 16671 18643 16677
rect 18708 16652 18736 16680
rect 18785 16677 18797 16711
rect 18831 16677 18843 16711
rect 18785 16671 18843 16677
rect 15749 16643 15807 16649
rect 15749 16640 15761 16643
rect 15212 16638 15761 16640
rect 15120 16612 15761 16638
rect 8944 16594 8996 16600
rect 13096 16581 13124 16612
rect 15120 16610 15240 16612
rect 15749 16609 15761 16612
rect 15795 16640 15807 16643
rect 15838 16640 15844 16652
rect 15795 16612 15844 16640
rect 15795 16609 15807 16612
rect 15749 16603 15807 16609
rect 15838 16600 15844 16612
rect 15896 16600 15902 16652
rect 15930 16600 15936 16652
rect 15988 16600 15994 16652
rect 16390 16600 16396 16652
rect 16448 16640 16454 16652
rect 16853 16643 16911 16649
rect 16853 16640 16865 16643
rect 16448 16612 16865 16640
rect 16448 16600 16454 16612
rect 16853 16609 16865 16612
rect 16899 16609 16911 16643
rect 16853 16603 16911 16609
rect 17338 16643 17396 16649
rect 17338 16609 17350 16643
rect 17384 16640 17396 16643
rect 18141 16643 18199 16649
rect 17384 16612 18092 16640
rect 17384 16609 17396 16612
rect 17338 16603 17396 16609
rect 7469 16575 7527 16581
rect 7469 16572 7481 16575
rect 6604 16544 6684 16572
rect 6748 16544 7481 16572
rect 6604 16532 6610 16544
rect 5276 16476 5580 16504
rect 5629 16507 5687 16513
rect 5629 16473 5641 16507
rect 5675 16473 5687 16507
rect 5629 16467 5687 16473
rect 6086 16464 6092 16516
rect 6144 16464 6150 16516
rect 6362 16464 6368 16516
rect 6420 16504 6426 16516
rect 6748 16504 6776 16544
rect 7469 16541 7481 16544
rect 7515 16541 7527 16575
rect 7469 16535 7527 16541
rect 7561 16575 7619 16581
rect 7561 16541 7573 16575
rect 7607 16572 7619 16575
rect 8021 16575 8079 16581
rect 8021 16572 8033 16575
rect 7607 16544 8033 16572
rect 7607 16541 7619 16544
rect 7561 16535 7619 16541
rect 8021 16541 8033 16544
rect 8067 16541 8079 16575
rect 8021 16535 8079 16541
rect 13081 16575 13139 16581
rect 13081 16541 13093 16575
rect 13127 16541 13139 16575
rect 13081 16535 13139 16541
rect 13446 16532 13452 16584
rect 13504 16532 13510 16584
rect 15286 16532 15292 16584
rect 15344 16572 15350 16584
rect 15948 16572 15976 16600
rect 15344 16544 15976 16572
rect 17129 16575 17187 16581
rect 15344 16532 15350 16544
rect 17129 16541 17141 16575
rect 17175 16541 17187 16575
rect 17129 16535 17187 16541
rect 6420 16476 6776 16504
rect 6420 16464 6426 16476
rect 7098 16464 7104 16516
rect 7156 16504 7162 16516
rect 8662 16504 8668 16516
rect 7156 16476 8668 16504
rect 7156 16464 7162 16476
rect 8662 16464 8668 16476
rect 8720 16464 8726 16516
rect 12897 16507 12955 16513
rect 12897 16473 12909 16507
rect 12943 16504 12955 16507
rect 13464 16504 13492 16532
rect 16574 16504 16580 16516
rect 12943 16476 13492 16504
rect 15212 16476 16580 16504
rect 12943 16473 12955 16476
rect 12897 16467 12955 16473
rect 1762 16396 1768 16448
rect 1820 16436 1826 16448
rect 1949 16439 2007 16445
rect 1949 16436 1961 16439
rect 1820 16408 1961 16436
rect 1820 16396 1826 16408
rect 1949 16405 1961 16408
rect 1995 16405 2007 16439
rect 1949 16399 2007 16405
rect 4706 16396 4712 16448
rect 4764 16396 4770 16448
rect 10321 16439 10379 16445
rect 10321 16405 10333 16439
rect 10367 16436 10379 16439
rect 10686 16436 10692 16448
rect 10367 16408 10692 16436
rect 10367 16405 10379 16408
rect 10321 16399 10379 16405
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 12986 16396 12992 16448
rect 13044 16396 13050 16448
rect 13078 16396 13084 16448
rect 13136 16436 13142 16448
rect 13354 16436 13360 16448
rect 13136 16408 13360 16436
rect 13136 16396 13142 16408
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 15212 16445 15240 16476
rect 16574 16464 16580 16476
rect 16632 16464 16638 16516
rect 17144 16504 17172 16535
rect 17218 16532 17224 16584
rect 17276 16532 17282 16584
rect 17494 16532 17500 16584
rect 17552 16572 17558 16584
rect 18064 16572 18092 16612
rect 18141 16609 18153 16643
rect 18187 16640 18199 16643
rect 18690 16640 18696 16652
rect 18187 16612 18696 16640
rect 18187 16609 18199 16612
rect 18141 16603 18199 16609
rect 18690 16600 18696 16612
rect 18748 16600 18754 16652
rect 19886 16600 19892 16652
rect 19944 16640 19950 16652
rect 19981 16643 20039 16649
rect 19981 16640 19993 16643
rect 19944 16612 19993 16640
rect 19944 16600 19950 16612
rect 19981 16609 19993 16612
rect 20027 16609 20039 16643
rect 19981 16603 20039 16609
rect 20162 16600 20168 16652
rect 20220 16600 20226 16652
rect 17552 16544 17980 16572
rect 18064 16544 18644 16572
rect 17552 16532 17558 16544
rect 17310 16504 17316 16516
rect 17144 16476 17316 16504
rect 17310 16464 17316 16476
rect 17368 16464 17374 16516
rect 15197 16439 15255 16445
rect 15197 16405 15209 16439
rect 15243 16405 15255 16439
rect 15197 16399 15255 16405
rect 15930 16396 15936 16448
rect 15988 16396 15994 16448
rect 17586 16396 17592 16448
rect 17644 16436 17650 16448
rect 17773 16439 17831 16445
rect 17773 16436 17785 16439
rect 17644 16408 17785 16436
rect 17644 16396 17650 16408
rect 17773 16405 17785 16408
rect 17819 16405 17831 16439
rect 17952 16436 17980 16544
rect 18616 16448 18644 16544
rect 19426 16532 19432 16584
rect 19484 16572 19490 16584
rect 20180 16572 20208 16600
rect 19484 16544 20208 16572
rect 19484 16532 19490 16544
rect 18417 16439 18475 16445
rect 18417 16436 18429 16439
rect 17952 16408 18429 16436
rect 17773 16399 17831 16405
rect 18417 16405 18429 16408
rect 18463 16405 18475 16439
rect 18417 16399 18475 16405
rect 18598 16396 18604 16448
rect 18656 16396 18662 16448
rect 20070 16396 20076 16448
rect 20128 16396 20134 16448
rect 552 16346 28428 16368
rect 552 16294 3882 16346
rect 3934 16294 3946 16346
rect 3998 16294 4010 16346
rect 4062 16294 4074 16346
rect 4126 16294 4138 16346
rect 4190 16294 10851 16346
rect 10903 16294 10915 16346
rect 10967 16294 10979 16346
rect 11031 16294 11043 16346
rect 11095 16294 11107 16346
rect 11159 16294 17820 16346
rect 17872 16294 17884 16346
rect 17936 16294 17948 16346
rect 18000 16294 18012 16346
rect 18064 16294 18076 16346
rect 18128 16294 24789 16346
rect 24841 16294 24853 16346
rect 24905 16294 24917 16346
rect 24969 16294 24981 16346
rect 25033 16294 25045 16346
rect 25097 16294 28428 16346
rect 552 16272 28428 16294
rect 3697 16235 3755 16241
rect 3697 16201 3709 16235
rect 3743 16232 3755 16235
rect 4522 16232 4528 16244
rect 3743 16204 4528 16232
rect 3743 16201 3755 16204
rect 3697 16195 3755 16201
rect 4522 16192 4528 16204
rect 4580 16192 4586 16244
rect 6730 16192 6736 16244
rect 6788 16192 6794 16244
rect 6822 16192 6828 16244
rect 6880 16192 6886 16244
rect 6914 16192 6920 16244
rect 6972 16192 6978 16244
rect 7285 16235 7343 16241
rect 7285 16201 7297 16235
rect 7331 16232 7343 16235
rect 7374 16232 7380 16244
rect 7331 16204 7380 16232
rect 7331 16201 7343 16204
rect 7285 16195 7343 16201
rect 7374 16192 7380 16204
rect 7432 16192 7438 16244
rect 9401 16235 9459 16241
rect 9401 16201 9413 16235
rect 9447 16232 9459 16235
rect 9582 16232 9588 16244
rect 9447 16204 9588 16232
rect 9447 16201 9459 16204
rect 9401 16195 9459 16201
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 15286 16192 15292 16244
rect 15344 16192 15350 16244
rect 16761 16235 16819 16241
rect 16761 16201 16773 16235
rect 16807 16201 16819 16235
rect 16761 16195 16819 16201
rect 2869 16167 2927 16173
rect 2869 16133 2881 16167
rect 2915 16164 2927 16167
rect 4430 16164 4436 16176
rect 2915 16136 4436 16164
rect 2915 16133 2927 16136
rect 2869 16127 2927 16133
rect 4430 16124 4436 16136
rect 4488 16124 4494 16176
rect 3234 16056 3240 16108
rect 3292 16096 3298 16108
rect 3329 16099 3387 16105
rect 3329 16096 3341 16099
rect 3292 16068 3341 16096
rect 3292 16056 3298 16068
rect 3329 16065 3341 16068
rect 3375 16065 3387 16099
rect 4448 16096 4476 16124
rect 4448 16068 4568 16096
rect 3329 16059 3387 16065
rect 1489 16031 1547 16037
rect 1489 15997 1501 16031
rect 1535 16028 1547 16031
rect 1578 16028 1584 16040
rect 1535 16000 1584 16028
rect 1535 15997 1547 16000
rect 1489 15991 1547 15997
rect 1578 15988 1584 16000
rect 1636 15988 1642 16040
rect 1762 16037 1768 16040
rect 1756 16028 1768 16037
rect 1723 16000 1768 16028
rect 1756 15991 1768 16000
rect 1762 15988 1768 15991
rect 1820 15988 1826 16040
rect 3421 16031 3479 16037
rect 3421 15997 3433 16031
rect 3467 16028 3479 16031
rect 3786 16028 3792 16040
rect 3467 16000 3792 16028
rect 3467 15997 3479 16000
rect 3421 15991 3479 15997
rect 3786 15988 3792 16000
rect 3844 15988 3850 16040
rect 4540 16037 4568 16068
rect 4433 16031 4491 16037
rect 4433 15997 4445 16031
rect 4479 15997 4491 16031
rect 4433 15991 4491 15997
rect 4525 16031 4583 16037
rect 4525 15997 4537 16031
rect 4571 15997 4583 16031
rect 4525 15991 4583 15997
rect 4246 15852 4252 15904
rect 4304 15852 4310 15904
rect 4448 15892 4476 15991
rect 4798 15988 4804 16040
rect 4856 15988 4862 16040
rect 5350 15988 5356 16040
rect 5408 15988 5414 16040
rect 6362 15988 6368 16040
rect 6420 16028 6426 16040
rect 6641 16031 6699 16037
rect 6641 16028 6653 16031
rect 6420 16000 6653 16028
rect 6420 15988 6426 16000
rect 6641 15997 6653 16000
rect 6687 16028 6699 16031
rect 6748 16028 6776 16192
rect 6687 16000 6776 16028
rect 6932 16028 6960 16192
rect 8662 16124 8668 16176
rect 8720 16164 8726 16176
rect 14369 16167 14427 16173
rect 8720 16136 9260 16164
rect 8720 16124 8726 16136
rect 8588 16068 9168 16096
rect 8588 16040 8616 16068
rect 7193 16031 7251 16037
rect 7193 16028 7205 16031
rect 6932 16000 7205 16028
rect 6687 15997 6699 16000
rect 6641 15991 6699 15997
rect 7193 15997 7205 16000
rect 7239 15997 7251 16031
rect 7377 16031 7435 16037
rect 7377 16028 7389 16031
rect 7193 15991 7251 15997
rect 7300 16000 7389 16028
rect 4614 15920 4620 15972
rect 4672 15920 4678 15972
rect 5368 15960 5396 15988
rect 5718 15960 5724 15972
rect 5368 15932 5724 15960
rect 5718 15920 5724 15932
rect 5776 15960 5782 15972
rect 6086 15960 6092 15972
rect 5776 15932 6092 15960
rect 5776 15920 5782 15932
rect 6086 15920 6092 15932
rect 6144 15960 6150 15972
rect 6546 15960 6552 15972
rect 6144 15932 6552 15960
rect 6144 15920 6150 15932
rect 6546 15920 6552 15932
rect 6604 15960 6610 15972
rect 6733 15963 6791 15969
rect 6733 15960 6745 15963
rect 6604 15932 6745 15960
rect 6604 15920 6610 15932
rect 6733 15929 6745 15932
rect 6779 15929 6791 15963
rect 6733 15923 6791 15929
rect 6917 15963 6975 15969
rect 6917 15929 6929 15963
rect 6963 15960 6975 15963
rect 7098 15960 7104 15972
rect 6963 15932 7104 15960
rect 6963 15929 6975 15932
rect 6917 15923 6975 15929
rect 7098 15920 7104 15932
rect 7156 15920 7162 15972
rect 7300 15904 7328 16000
rect 7377 15997 7389 16000
rect 7423 15997 7435 16031
rect 7377 15991 7435 15997
rect 8570 15988 8576 16040
rect 8628 15988 8634 16040
rect 8849 16031 8907 16037
rect 8849 15997 8861 16031
rect 8895 15997 8907 16031
rect 8849 15991 8907 15997
rect 8754 15920 8760 15972
rect 8812 15960 8818 15972
rect 8864 15960 8892 15991
rect 8938 15988 8944 16040
rect 8996 15988 9002 16040
rect 9140 16037 9168 16068
rect 9232 16037 9260 16136
rect 14369 16133 14381 16167
rect 14415 16164 14427 16167
rect 14415 16136 15700 16164
rect 14415 16133 14427 16136
rect 14369 16127 14427 16133
rect 11793 16099 11851 16105
rect 11793 16065 11805 16099
rect 11839 16096 11851 16099
rect 11882 16096 11888 16108
rect 11839 16068 11888 16096
rect 11839 16065 11851 16068
rect 11793 16059 11851 16065
rect 11882 16056 11888 16068
rect 11940 16056 11946 16108
rect 14093 16099 14151 16105
rect 14093 16065 14105 16099
rect 14139 16096 14151 16099
rect 14826 16096 14832 16108
rect 14139 16068 14832 16096
rect 14139 16065 14151 16068
rect 14093 16059 14151 16065
rect 14826 16056 14832 16068
rect 14884 16096 14890 16108
rect 14884 16068 15240 16096
rect 14884 16056 14890 16068
rect 9125 16031 9183 16037
rect 9125 15997 9137 16031
rect 9171 15997 9183 16031
rect 9125 15991 9183 15997
rect 9217 16031 9275 16037
rect 9217 15997 9229 16031
rect 9263 15997 9275 16031
rect 9217 15991 9275 15997
rect 10686 15988 10692 16040
rect 10744 16028 10750 16040
rect 10974 16031 11032 16037
rect 10974 16028 10986 16031
rect 10744 16000 10986 16028
rect 10744 15988 10750 16000
rect 10974 15997 10986 16000
rect 11020 15997 11032 16031
rect 10974 15991 11032 15997
rect 11238 15988 11244 16040
rect 11296 15988 11302 16040
rect 11606 15988 11612 16040
rect 11664 15988 11670 16040
rect 12897 16031 12955 16037
rect 12897 15997 12909 16031
rect 12943 15997 12955 16031
rect 12897 15991 12955 15997
rect 8812 15932 8892 15960
rect 12912 15960 12940 15991
rect 12986 15988 12992 16040
rect 13044 16028 13050 16040
rect 13081 16031 13139 16037
rect 13081 16028 13093 16031
rect 13044 16000 13093 16028
rect 13044 15988 13050 16000
rect 13081 15997 13093 16000
rect 13127 15997 13139 16031
rect 13081 15991 13139 15997
rect 13170 15988 13176 16040
rect 13228 15988 13234 16040
rect 13262 15988 13268 16040
rect 13320 16028 13326 16040
rect 13725 16031 13783 16037
rect 13725 16028 13737 16031
rect 13320 16000 13737 16028
rect 13320 15988 13326 16000
rect 13725 15997 13737 16000
rect 13771 15997 13783 16031
rect 13725 15991 13783 15997
rect 13998 15988 14004 16040
rect 14056 15988 14062 16040
rect 15212 16037 15240 16068
rect 15105 16031 15163 16037
rect 15105 16028 15117 16031
rect 15028 16000 15117 16028
rect 13538 15960 13544 15972
rect 12912 15932 13544 15960
rect 8812 15920 8818 15932
rect 13096 15904 13124 15932
rect 13538 15920 13544 15932
rect 13596 15920 13602 15972
rect 15028 15904 15056 16000
rect 15105 15997 15117 16000
rect 15151 15997 15163 16031
rect 15105 15991 15163 15997
rect 15197 16031 15255 16037
rect 15197 15997 15209 16031
rect 15243 15997 15255 16031
rect 15473 16031 15531 16037
rect 15473 16028 15485 16031
rect 15197 15991 15255 15997
rect 15396 16000 15485 16028
rect 15396 15969 15424 16000
rect 15473 15997 15485 16000
rect 15519 16028 15531 16031
rect 15562 16028 15568 16040
rect 15519 16000 15568 16028
rect 15519 15997 15531 16000
rect 15473 15991 15531 15997
rect 15562 15988 15568 16000
rect 15620 15988 15626 16040
rect 15672 16028 15700 16136
rect 15746 16124 15752 16176
rect 15804 16124 15810 16176
rect 16776 16164 16804 16195
rect 17402 16192 17408 16244
rect 17460 16232 17466 16244
rect 17497 16235 17555 16241
rect 17497 16232 17509 16235
rect 17460 16204 17509 16232
rect 17460 16192 17466 16204
rect 17497 16201 17509 16204
rect 17543 16201 17555 16235
rect 17497 16195 17555 16201
rect 17604 16204 17727 16232
rect 17604 16164 17632 16204
rect 16776 16136 17632 16164
rect 17699 16096 17727 16204
rect 17954 16192 17960 16244
rect 18012 16192 18018 16244
rect 18782 16192 18788 16244
rect 18840 16232 18846 16244
rect 19981 16235 20039 16241
rect 19981 16232 19993 16235
rect 18840 16204 19993 16232
rect 18840 16192 18846 16204
rect 19981 16201 19993 16204
rect 20027 16232 20039 16235
rect 20027 16204 21956 16232
rect 20027 16201 20039 16204
rect 19981 16195 20039 16201
rect 20530 16124 20536 16176
rect 20588 16124 20594 16176
rect 21928 16105 21956 16204
rect 21913 16099 21971 16105
rect 17699 16068 17816 16096
rect 15749 16031 15807 16037
rect 15749 16028 15761 16031
rect 15672 16000 15761 16028
rect 15749 15997 15761 16000
rect 15795 16028 15807 16031
rect 16574 16028 16580 16040
rect 15795 16000 16580 16028
rect 15795 15997 15807 16000
rect 15749 15991 15807 15997
rect 16574 15988 16580 16000
rect 16632 15988 16638 16040
rect 17034 15988 17040 16040
rect 17092 15988 17098 16040
rect 17126 15988 17132 16040
rect 17184 15988 17190 16040
rect 17221 16031 17279 16037
rect 17221 15997 17233 16031
rect 17267 15997 17279 16031
rect 17381 16031 17439 16037
rect 17381 16028 17393 16031
rect 17221 15991 17279 15997
rect 17353 15997 17393 16028
rect 17427 16022 17439 16031
rect 17494 16022 17500 16040
rect 17427 15997 17500 16022
rect 17353 15994 17500 15997
rect 17381 15991 17439 15994
rect 15381 15963 15439 15969
rect 15381 15929 15393 15963
rect 15427 15929 15439 15963
rect 15381 15923 15439 15929
rect 4706 15892 4712 15904
rect 4448 15864 4712 15892
rect 4706 15852 4712 15864
rect 4764 15852 4770 15904
rect 7282 15852 7288 15904
rect 7340 15852 7346 15904
rect 9858 15852 9864 15904
rect 9916 15852 9922 15904
rect 11422 15852 11428 15904
rect 11480 15852 11486 15904
rect 12713 15895 12771 15901
rect 12713 15861 12725 15895
rect 12759 15892 12771 15895
rect 12802 15892 12808 15904
rect 12759 15864 12808 15892
rect 12759 15861 12771 15864
rect 12713 15855 12771 15861
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 13078 15852 13084 15904
rect 13136 15852 13142 15904
rect 13630 15852 13636 15904
rect 13688 15852 13694 15904
rect 15010 15852 15016 15904
rect 15068 15892 15074 15904
rect 15565 15895 15623 15901
rect 15565 15892 15577 15895
rect 15068 15864 15577 15892
rect 15068 15852 15074 15864
rect 15565 15861 15577 15864
rect 15611 15861 15623 15895
rect 17236 15892 17264 15991
rect 17494 15988 17500 15994
rect 17552 15988 17558 16040
rect 17663 16031 17721 16037
rect 17663 15997 17675 16031
rect 17709 16028 17721 16031
rect 17709 15997 17724 16028
rect 17663 15991 17724 15997
rect 17586 15892 17592 15904
rect 17236 15864 17592 15892
rect 15565 15855 15623 15861
rect 17586 15852 17592 15864
rect 17644 15852 17650 15904
rect 17696 15892 17724 15991
rect 17788 15960 17816 16068
rect 21913 16065 21925 16099
rect 21959 16096 21971 16099
rect 22094 16096 22100 16108
rect 21959 16068 22100 16096
rect 21959 16065 21971 16068
rect 21913 16059 21971 16065
rect 22094 16056 22100 16068
rect 22152 16096 22158 16108
rect 22922 16096 22928 16108
rect 22152 16068 22928 16096
rect 22152 16056 22158 16068
rect 22922 16056 22928 16068
rect 22980 16056 22986 16108
rect 17862 15988 17868 16040
rect 17920 15988 17926 16040
rect 18506 15988 18512 16040
rect 18564 16028 18570 16040
rect 18693 16031 18751 16037
rect 18693 16028 18705 16031
rect 18564 16000 18705 16028
rect 18564 15988 18570 16000
rect 18693 15997 18705 16000
rect 18739 15997 18751 16031
rect 18693 15991 18751 15997
rect 18141 15963 18199 15969
rect 18141 15960 18153 15963
rect 17788 15932 18153 15960
rect 18141 15929 18153 15932
rect 18187 15929 18199 15963
rect 18141 15923 18199 15929
rect 20162 15920 20168 15972
rect 20220 15960 20226 15972
rect 21646 15963 21704 15969
rect 21646 15960 21658 15963
rect 20220 15932 21658 15960
rect 20220 15920 20226 15932
rect 21646 15929 21658 15932
rect 21692 15929 21704 15963
rect 21646 15923 21704 15929
rect 17770 15892 17776 15904
rect 17696 15864 17776 15892
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 552 15802 28587 15824
rect 552 15750 7366 15802
rect 7418 15750 7430 15802
rect 7482 15750 7494 15802
rect 7546 15750 7558 15802
rect 7610 15750 7622 15802
rect 7674 15750 14335 15802
rect 14387 15750 14399 15802
rect 14451 15750 14463 15802
rect 14515 15750 14527 15802
rect 14579 15750 14591 15802
rect 14643 15750 21304 15802
rect 21356 15750 21368 15802
rect 21420 15750 21432 15802
rect 21484 15750 21496 15802
rect 21548 15750 21560 15802
rect 21612 15750 28273 15802
rect 28325 15750 28337 15802
rect 28389 15750 28401 15802
rect 28453 15750 28465 15802
rect 28517 15750 28529 15802
rect 28581 15750 28587 15802
rect 552 15728 28587 15750
rect 2130 15648 2136 15700
rect 2188 15648 2194 15700
rect 4246 15688 4252 15700
rect 2746 15660 4252 15688
rect 2317 15555 2375 15561
rect 2317 15521 2329 15555
rect 2363 15552 2375 15555
rect 2746 15552 2774 15660
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 6454 15648 6460 15700
rect 6512 15688 6518 15700
rect 6641 15691 6699 15697
rect 6641 15688 6653 15691
rect 6512 15660 6653 15688
rect 6512 15648 6518 15660
rect 6641 15657 6653 15660
rect 6687 15657 6699 15691
rect 6641 15651 6699 15657
rect 13170 15648 13176 15700
rect 13228 15688 13234 15700
rect 13265 15691 13323 15697
rect 13265 15688 13277 15691
rect 13228 15660 13277 15688
rect 13228 15648 13234 15660
rect 13265 15657 13277 15660
rect 13311 15657 13323 15691
rect 13265 15651 13323 15657
rect 13630 15648 13636 15700
rect 13688 15648 13694 15700
rect 17310 15648 17316 15700
rect 17368 15648 17374 15700
rect 17589 15691 17647 15697
rect 17589 15657 17601 15691
rect 17635 15688 17647 15691
rect 17954 15688 17960 15700
rect 17635 15660 17960 15688
rect 17635 15657 17647 15660
rect 17589 15651 17647 15657
rect 17954 15648 17960 15660
rect 18012 15648 18018 15700
rect 20070 15648 20076 15700
rect 20128 15648 20134 15700
rect 20162 15648 20168 15700
rect 20220 15648 20226 15700
rect 20530 15648 20536 15700
rect 20588 15648 20594 15700
rect 6181 15623 6239 15629
rect 6181 15589 6193 15623
rect 6227 15620 6239 15623
rect 6227 15592 6592 15620
rect 6227 15589 6239 15592
rect 6181 15583 6239 15589
rect 2363 15524 2774 15552
rect 2363 15521 2375 15524
rect 2317 15515 2375 15521
rect 4522 15512 4528 15564
rect 4580 15552 4586 15564
rect 5077 15555 5135 15561
rect 5077 15552 5089 15555
rect 4580 15524 5089 15552
rect 4580 15512 4586 15524
rect 5077 15521 5089 15524
rect 5123 15552 5135 15555
rect 5442 15552 5448 15564
rect 5123 15524 5448 15552
rect 5123 15521 5135 15524
rect 5077 15515 5135 15521
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 6086 15561 6092 15564
rect 6079 15555 6092 15561
rect 6079 15552 6091 15555
rect 6047 15524 6091 15552
rect 6079 15521 6091 15524
rect 6079 15515 6092 15521
rect 6086 15512 6092 15515
rect 6144 15512 6150 15564
rect 6273 15555 6331 15561
rect 6273 15521 6285 15555
rect 6319 15552 6331 15555
rect 6362 15552 6368 15564
rect 6319 15524 6368 15552
rect 6319 15521 6331 15524
rect 6273 15515 6331 15521
rect 2406 15444 2412 15496
rect 2464 15484 2470 15496
rect 2501 15487 2559 15493
rect 2501 15484 2513 15487
rect 2464 15456 2513 15484
rect 2464 15444 2470 15456
rect 2501 15453 2513 15456
rect 2547 15484 2559 15487
rect 2547 15456 2774 15484
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 2746 15348 2774 15456
rect 5166 15444 5172 15496
rect 5224 15484 5230 15496
rect 6288 15484 6316 15515
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 6564 15561 6592 15592
rect 6549 15555 6607 15561
rect 6549 15521 6561 15555
rect 6595 15521 6607 15555
rect 6549 15515 6607 15521
rect 6733 15555 6791 15561
rect 6733 15521 6745 15555
rect 6779 15552 6791 15555
rect 7466 15552 7472 15564
rect 6779 15524 7472 15552
rect 6779 15521 6791 15524
rect 6733 15515 6791 15521
rect 7466 15512 7472 15524
rect 7524 15552 7530 15564
rect 9033 15555 9091 15561
rect 9033 15552 9045 15555
rect 7524 15524 9045 15552
rect 7524 15512 7530 15524
rect 9033 15521 9045 15524
rect 9079 15521 9091 15555
rect 9033 15515 9091 15521
rect 13446 15512 13452 15564
rect 13504 15512 13510 15564
rect 13541 15555 13599 15561
rect 13541 15521 13553 15555
rect 13587 15552 13599 15555
rect 13648 15552 13676 15648
rect 17328 15620 17356 15648
rect 20088 15620 20116 15648
rect 17328 15592 17448 15620
rect 13587 15524 13676 15552
rect 16945 15555 17003 15561
rect 13587 15521 13599 15524
rect 13541 15515 13599 15521
rect 16945 15521 16957 15555
rect 16991 15521 17003 15555
rect 16945 15515 17003 15521
rect 5224 15456 6316 15484
rect 5224 15444 5230 15456
rect 8570 15444 8576 15496
rect 8628 15444 8634 15496
rect 8662 15444 8668 15496
rect 8720 15484 8726 15496
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8720 15456 8953 15484
rect 8720 15444 8726 15456
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 13265 15487 13323 15493
rect 13265 15453 13277 15487
rect 13311 15484 13323 15487
rect 14182 15484 14188 15496
rect 13311 15456 14188 15484
rect 13311 15453 13323 15456
rect 13265 15447 13323 15453
rect 14182 15444 14188 15456
rect 14240 15444 14246 15496
rect 3786 15376 3792 15428
rect 3844 15416 3850 15428
rect 4709 15419 4767 15425
rect 4709 15416 4721 15419
rect 3844 15388 4721 15416
rect 3844 15376 3850 15388
rect 4709 15385 4721 15388
rect 4755 15385 4767 15419
rect 4709 15379 4767 15385
rect 9674 15376 9680 15428
rect 9732 15416 9738 15428
rect 10686 15416 10692 15428
rect 9732 15388 10692 15416
rect 9732 15376 9738 15388
rect 10686 15376 10692 15388
rect 10744 15376 10750 15428
rect 16960 15416 16988 15515
rect 17034 15512 17040 15564
rect 17092 15552 17098 15564
rect 17092 15524 17137 15552
rect 17092 15512 17098 15524
rect 17218 15512 17224 15564
rect 17276 15512 17282 15564
rect 17420 15561 17448 15592
rect 19720 15592 20116 15620
rect 20548 15620 20576 15648
rect 20548 15592 20944 15620
rect 17313 15555 17371 15561
rect 17313 15521 17325 15555
rect 17359 15521 17371 15555
rect 17313 15515 17371 15521
rect 17410 15555 17468 15561
rect 17410 15521 17422 15555
rect 17456 15521 17468 15555
rect 17957 15555 18015 15561
rect 17957 15552 17969 15555
rect 17410 15515 17468 15521
rect 17512 15524 17969 15552
rect 17328 15484 17356 15515
rect 17512 15484 17540 15524
rect 17957 15521 17969 15524
rect 18003 15552 18015 15555
rect 18003 15524 19012 15552
rect 18003 15521 18015 15524
rect 17957 15515 18015 15521
rect 17328 15456 17540 15484
rect 17681 15487 17739 15493
rect 17681 15453 17693 15487
rect 17727 15484 17739 15487
rect 18138 15484 18144 15496
rect 17727 15456 18144 15484
rect 17727 15453 17739 15456
rect 17681 15447 17739 15453
rect 18138 15444 18144 15456
rect 18196 15444 18202 15496
rect 18690 15444 18696 15496
rect 18748 15444 18754 15496
rect 18984 15493 19012 15524
rect 19058 15512 19064 15564
rect 19116 15512 19122 15564
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 19720 15561 19748 15592
rect 19521 15555 19579 15561
rect 19521 15552 19533 15555
rect 19392 15524 19533 15552
rect 19392 15512 19398 15524
rect 19521 15521 19533 15524
rect 19567 15521 19579 15555
rect 19521 15515 19579 15521
rect 19705 15555 19763 15561
rect 19705 15521 19717 15555
rect 19751 15521 19763 15555
rect 19705 15515 19763 15521
rect 19797 15555 19855 15561
rect 19797 15521 19809 15555
rect 19843 15521 19855 15555
rect 19797 15515 19855 15521
rect 18969 15487 19027 15493
rect 18969 15453 18981 15487
rect 19015 15484 19027 15487
rect 19015 15456 19104 15484
rect 19015 15453 19027 15456
rect 18969 15447 19027 15453
rect 17773 15419 17831 15425
rect 17773 15416 17785 15419
rect 16960 15388 17785 15416
rect 17773 15385 17785 15388
rect 17819 15385 17831 15419
rect 17773 15379 17831 15385
rect 19076 15360 19104 15456
rect 19812 15416 19840 15515
rect 19886 15512 19892 15564
rect 19944 15512 19950 15564
rect 19978 15512 19984 15564
rect 20036 15552 20042 15564
rect 20257 15555 20315 15561
rect 20257 15552 20269 15555
rect 20036 15524 20269 15552
rect 20036 15512 20042 15524
rect 20257 15521 20269 15524
rect 20303 15521 20315 15555
rect 20257 15515 20315 15521
rect 20622 15512 20628 15564
rect 20680 15512 20686 15564
rect 20916 15561 20944 15592
rect 20990 15580 20996 15632
rect 21048 15620 21054 15632
rect 22462 15620 22468 15632
rect 21048 15592 22468 15620
rect 21048 15580 21054 15592
rect 22462 15580 22468 15592
rect 22520 15580 22526 15632
rect 20901 15555 20959 15561
rect 20901 15521 20913 15555
rect 20947 15521 20959 15555
rect 20901 15515 20959 15521
rect 21266 15512 21272 15564
rect 21324 15512 21330 15564
rect 22750 15555 22808 15561
rect 22750 15552 22762 15555
rect 21468 15524 22762 15552
rect 19904 15484 19932 15512
rect 20441 15487 20499 15493
rect 20441 15484 20453 15487
rect 19904 15456 20453 15484
rect 20441 15453 20453 15456
rect 20487 15484 20499 15487
rect 20993 15487 21051 15493
rect 20993 15484 21005 15487
rect 20487 15456 21005 15484
rect 20487 15453 20499 15456
rect 20441 15447 20499 15453
rect 20993 15453 21005 15456
rect 21039 15453 21051 15487
rect 20993 15447 21051 15453
rect 21468 15425 21496 15524
rect 22750 15521 22762 15524
rect 22796 15521 22808 15555
rect 22750 15515 22808 15521
rect 22922 15512 22928 15564
rect 22980 15552 22986 15564
rect 23017 15555 23075 15561
rect 23017 15552 23029 15555
rect 22980 15524 23029 15552
rect 22980 15512 22986 15524
rect 23017 15521 23029 15524
rect 23063 15521 23075 15555
rect 23017 15515 23075 15521
rect 21453 15419 21511 15425
rect 19812 15388 20300 15416
rect 20272 15360 20300 15388
rect 21453 15385 21465 15419
rect 21499 15385 21511 15419
rect 21453 15379 21511 15385
rect 3326 15348 3332 15360
rect 2746 15320 3332 15348
rect 3326 15308 3332 15320
rect 3384 15348 3390 15360
rect 5810 15348 5816 15360
rect 3384 15320 5816 15348
rect 3384 15308 3390 15320
rect 5810 15308 5816 15320
rect 5868 15308 5874 15360
rect 9217 15351 9275 15357
rect 9217 15317 9229 15351
rect 9263 15348 9275 15351
rect 11974 15348 11980 15360
rect 9263 15320 11980 15348
rect 9263 15317 9275 15320
rect 9217 15311 9275 15317
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 17310 15308 17316 15360
rect 17368 15348 17374 15360
rect 17865 15351 17923 15357
rect 17865 15348 17877 15351
rect 17368 15320 17877 15348
rect 17368 15308 17374 15320
rect 17865 15317 17877 15320
rect 17911 15317 17923 15351
rect 17865 15311 17923 15317
rect 19058 15308 19064 15360
rect 19116 15308 19122 15360
rect 20254 15308 20260 15360
rect 20312 15308 20318 15360
rect 20346 15308 20352 15360
rect 20404 15308 20410 15360
rect 21634 15308 21640 15360
rect 21692 15308 21698 15360
rect 552 15258 28428 15280
rect 552 15206 3882 15258
rect 3934 15206 3946 15258
rect 3998 15206 4010 15258
rect 4062 15206 4074 15258
rect 4126 15206 4138 15258
rect 4190 15206 10851 15258
rect 10903 15206 10915 15258
rect 10967 15206 10979 15258
rect 11031 15206 11043 15258
rect 11095 15206 11107 15258
rect 11159 15206 17820 15258
rect 17872 15206 17884 15258
rect 17936 15206 17948 15258
rect 18000 15206 18012 15258
rect 18064 15206 18076 15258
rect 18128 15206 24789 15258
rect 24841 15206 24853 15258
rect 24905 15206 24917 15258
rect 24969 15206 24981 15258
rect 25033 15206 25045 15258
rect 25097 15206 28428 15258
rect 552 15184 28428 15206
rect 4430 15144 4436 15156
rect 2056 15116 4436 15144
rect 2056 15017 2084 15116
rect 2976 15085 3004 15116
rect 4430 15104 4436 15116
rect 4488 15104 4494 15156
rect 7466 15104 7472 15156
rect 7524 15104 7530 15156
rect 8570 15104 8576 15156
rect 8628 15144 8634 15156
rect 8665 15147 8723 15153
rect 8665 15144 8677 15147
rect 8628 15116 8677 15144
rect 8628 15104 8634 15116
rect 8665 15113 8677 15116
rect 8711 15144 8723 15147
rect 8849 15147 8907 15153
rect 8849 15144 8861 15147
rect 8711 15116 8861 15144
rect 8711 15113 8723 15116
rect 8665 15107 8723 15113
rect 8849 15113 8861 15116
rect 8895 15113 8907 15147
rect 8849 15107 8907 15113
rect 10428 15116 11551 15144
rect 2409 15079 2467 15085
rect 2409 15045 2421 15079
rect 2455 15045 2467 15079
rect 2409 15039 2467 15045
rect 2961 15079 3019 15085
rect 2961 15045 2973 15079
rect 3007 15045 3019 15079
rect 2961 15039 3019 15045
rect 3053 15079 3111 15085
rect 3053 15045 3065 15079
rect 3099 15076 3111 15079
rect 3142 15076 3148 15088
rect 3099 15048 3148 15076
rect 3099 15045 3111 15048
rect 3053 15039 3111 15045
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 14977 2099 15011
rect 2041 14971 2099 14977
rect 2424 14940 2452 15039
rect 3142 15036 3148 15048
rect 3200 15076 3206 15088
rect 3200 15048 3464 15076
rect 3200 15036 3206 15048
rect 2501 15011 2559 15017
rect 2501 14977 2513 15011
rect 2547 15008 2559 15011
rect 2547 14980 3280 15008
rect 2547 14977 2559 14980
rect 2501 14971 2559 14977
rect 2593 14943 2651 14949
rect 2593 14940 2605 14943
rect 2424 14912 2605 14940
rect 2593 14909 2605 14912
rect 2639 14940 2651 14943
rect 3050 14940 3056 14952
rect 2639 14912 3056 14940
rect 2639 14909 2651 14912
rect 2593 14903 2651 14909
rect 3050 14900 3056 14912
rect 3108 14900 3114 14952
rect 3252 14949 3280 14980
rect 3436 14949 3464 15048
rect 3605 15011 3663 15017
rect 3605 14977 3617 15011
rect 3651 15008 3663 15011
rect 4157 15011 4215 15017
rect 4157 15008 4169 15011
rect 3651 14980 4169 15008
rect 3651 14977 3663 14980
rect 3605 14971 3663 14977
rect 4157 14977 4169 14980
rect 4203 14977 4215 15011
rect 4448 15008 4476 15104
rect 7285 15079 7343 15085
rect 7285 15045 7297 15079
rect 7331 15045 7343 15079
rect 7285 15039 7343 15045
rect 9217 15079 9275 15085
rect 9217 15045 9229 15079
rect 9263 15076 9275 15079
rect 10428 15076 10456 15116
rect 9263 15048 10456 15076
rect 9263 15045 9275 15048
rect 9217 15039 9275 15045
rect 4448 14980 4844 15008
rect 4157 14971 4215 14977
rect 3237 14943 3295 14949
rect 3237 14909 3249 14943
rect 3283 14909 3295 14943
rect 3237 14903 3295 14909
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14909 3479 14943
rect 3421 14903 3479 14909
rect 3694 14900 3700 14952
rect 3752 14900 3758 14952
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14909 3847 14943
rect 3789 14903 3847 14909
rect 3329 14875 3387 14881
rect 3329 14841 3341 14875
rect 3375 14872 3387 14875
rect 3804 14872 3832 14903
rect 3878 14900 3884 14952
rect 3936 14900 3942 14952
rect 4341 14943 4399 14949
rect 4341 14909 4353 14943
rect 4387 14940 4399 14943
rect 4522 14940 4528 14952
rect 4387 14912 4528 14940
rect 4387 14909 4399 14912
rect 4341 14903 4399 14909
rect 4522 14900 4528 14912
rect 4580 14900 4586 14952
rect 4816 14949 4844 14980
rect 4617 14943 4675 14949
rect 4617 14909 4629 14943
rect 4663 14909 4675 14943
rect 4617 14903 4675 14909
rect 4801 14943 4859 14949
rect 4801 14909 4813 14943
rect 4847 14909 4859 14943
rect 4801 14903 4859 14909
rect 3375 14844 3832 14872
rect 4632 14872 4660 14903
rect 5166 14900 5172 14952
rect 5224 14900 5230 14952
rect 5902 14900 5908 14952
rect 5960 14900 5966 14952
rect 7300 14940 7328 15039
rect 8938 15008 8944 15020
rect 8496 14980 8944 15008
rect 8496 14949 8524 14980
rect 8938 14968 8944 14980
rect 8996 15008 9002 15020
rect 8996 14980 9628 15008
rect 8996 14968 9002 14980
rect 9600 14952 9628 14980
rect 9766 14968 9772 15020
rect 9824 14968 9830 15020
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 15008 10103 15011
rect 10091 14980 10180 15008
rect 10091 14977 10103 14980
rect 10045 14971 10103 14977
rect 7837 14943 7895 14949
rect 7837 14940 7849 14943
rect 7300 14912 7849 14940
rect 7837 14909 7849 14912
rect 7883 14940 7895 14943
rect 7929 14943 7987 14949
rect 7929 14940 7941 14943
rect 7883 14912 7941 14940
rect 7883 14909 7895 14912
rect 7837 14903 7895 14909
rect 7929 14909 7941 14912
rect 7975 14909 7987 14943
rect 7929 14903 7987 14909
rect 8481 14943 8539 14949
rect 8481 14909 8493 14943
rect 8527 14909 8539 14943
rect 8481 14903 8539 14909
rect 8665 14943 8723 14949
rect 8665 14909 8677 14943
rect 8711 14909 8723 14943
rect 8665 14903 8723 14909
rect 8757 14943 8815 14949
rect 8757 14909 8769 14943
rect 8803 14940 8815 14943
rect 9033 14943 9091 14949
rect 8803 14912 8984 14940
rect 8803 14909 8815 14912
rect 8757 14903 8815 14909
rect 5184 14872 5212 14900
rect 4632 14844 5212 14872
rect 6172 14875 6230 14881
rect 3375 14841 3387 14844
rect 3329 14835 3387 14841
rect 3436 14816 3464 14844
rect 6172 14841 6184 14875
rect 6218 14872 6230 14875
rect 6270 14872 6276 14884
rect 6218 14844 6276 14872
rect 6218 14841 6230 14844
rect 6172 14835 6230 14841
rect 6270 14832 6276 14844
rect 6328 14832 6334 14884
rect 6362 14832 6368 14884
rect 6420 14872 6426 14884
rect 7653 14875 7711 14881
rect 7653 14872 7665 14875
rect 6420 14844 7665 14872
rect 6420 14832 6426 14844
rect 7653 14841 7665 14844
rect 7699 14841 7711 14875
rect 8680 14872 8708 14903
rect 8680 14844 8800 14872
rect 7653 14835 7711 14841
rect 8772 14816 8800 14844
rect 8956 14816 8984 14912
rect 9033 14909 9045 14943
rect 9079 14909 9091 14943
rect 9033 14903 9091 14909
rect 9048 14872 9076 14903
rect 9582 14900 9588 14952
rect 9640 14900 9646 14952
rect 9677 14943 9735 14949
rect 9677 14909 9689 14943
rect 9723 14940 9735 14943
rect 9950 14940 9956 14952
rect 9723 14912 9956 14940
rect 9723 14909 9735 14912
rect 9677 14903 9735 14909
rect 9950 14900 9956 14912
rect 10008 14900 10014 14952
rect 10152 14872 10180 14980
rect 10229 14943 10287 14949
rect 10229 14909 10241 14943
rect 10275 14940 10287 14943
rect 10428 14940 10456 15048
rect 10505 15079 10563 15085
rect 10505 15045 10517 15079
rect 10551 15045 10563 15079
rect 10505 15039 10563 15045
rect 10520 15008 10548 15039
rect 10686 15036 10692 15088
rect 10744 15076 10750 15088
rect 10744 15048 10916 15076
rect 10744 15036 10750 15048
rect 10781 15011 10839 15017
rect 10781 15008 10793 15011
rect 10520 14980 10793 15008
rect 10781 14977 10793 14980
rect 10827 14977 10839 15011
rect 10888 15008 10916 15048
rect 11241 15011 11299 15017
rect 11241 15008 11253 15011
rect 10888 14980 11253 15008
rect 10781 14971 10839 14977
rect 11241 14977 11253 14980
rect 11287 15008 11299 15011
rect 11330 15008 11336 15020
rect 11287 14980 11336 15008
rect 11287 14977 11299 14980
rect 11241 14971 11299 14977
rect 11330 14968 11336 14980
rect 11388 14968 11394 15020
rect 11523 15008 11551 15116
rect 12066 15104 12072 15156
rect 12124 15104 12130 15156
rect 19978 15104 19984 15156
rect 20036 15104 20042 15156
rect 21266 15104 21272 15156
rect 21324 15144 21330 15156
rect 21637 15147 21695 15153
rect 21637 15144 21649 15147
rect 21324 15116 21649 15144
rect 21324 15104 21330 15116
rect 21637 15113 21649 15116
rect 21683 15113 21695 15147
rect 21637 15107 21695 15113
rect 13906 15036 13912 15088
rect 13964 15076 13970 15088
rect 16025 15079 16083 15085
rect 13964 15048 15976 15076
rect 13964 15036 13970 15048
rect 11609 15011 11667 15017
rect 11609 15008 11621 15011
rect 11523 14980 11621 15008
rect 11609 14977 11621 14980
rect 11655 14977 11667 15011
rect 11609 14971 11667 14977
rect 11790 14968 11796 15020
rect 11848 14968 11854 15020
rect 14277 15011 14335 15017
rect 14277 15008 14289 15011
rect 12544 14980 14289 15008
rect 12245 14953 12303 14959
rect 10275 14912 10456 14940
rect 10873 14943 10931 14949
rect 10275 14909 10287 14912
rect 10229 14903 10287 14909
rect 10873 14909 10885 14943
rect 10919 14909 10931 14943
rect 10873 14903 10931 14909
rect 11149 14943 11207 14949
rect 11149 14909 11161 14943
rect 11195 14909 11207 14943
rect 11149 14903 11207 14909
rect 11518 14943 11576 14949
rect 11518 14909 11530 14943
rect 11564 14940 11576 14943
rect 11564 14912 11652 14940
rect 11564 14909 11576 14912
rect 11518 14903 11576 14909
rect 10505 14875 10563 14881
rect 10505 14872 10517 14875
rect 9048 14844 9720 14872
rect 10152 14844 10517 14872
rect 9692 14816 9720 14844
rect 10505 14841 10517 14844
rect 10551 14872 10563 14875
rect 10551 14844 10732 14872
rect 10551 14841 10563 14844
rect 10505 14835 10563 14841
rect 10704 14816 10732 14844
rect 3418 14764 3424 14816
rect 3476 14764 3482 14816
rect 4065 14807 4123 14813
rect 4065 14773 4077 14807
rect 4111 14804 4123 14807
rect 6086 14804 6092 14816
rect 4111 14776 6092 14804
rect 4111 14773 4123 14776
rect 4065 14767 4123 14773
rect 6086 14764 6092 14776
rect 6144 14764 6150 14816
rect 7742 14764 7748 14816
rect 7800 14804 7806 14816
rect 8113 14807 8171 14813
rect 8113 14804 8125 14807
rect 7800 14776 8125 14804
rect 7800 14764 7806 14776
rect 8113 14773 8125 14776
rect 8159 14773 8171 14807
rect 8113 14767 8171 14773
rect 8754 14764 8760 14816
rect 8812 14764 8818 14816
rect 8938 14764 8944 14816
rect 8996 14764 9002 14816
rect 9674 14764 9680 14816
rect 9732 14764 9738 14816
rect 10318 14764 10324 14816
rect 10376 14764 10382 14816
rect 10594 14764 10600 14816
rect 10652 14764 10658 14816
rect 10686 14764 10692 14816
rect 10744 14764 10750 14816
rect 10888 14804 10916 14903
rect 11164 14872 11192 14903
rect 11164 14844 11560 14872
rect 11532 14816 11560 14844
rect 11333 14807 11391 14813
rect 11333 14804 11345 14807
rect 10888 14776 11345 14804
rect 11333 14773 11345 14776
rect 11379 14773 11391 14807
rect 11333 14767 11391 14773
rect 11514 14764 11520 14816
rect 11572 14764 11578 14816
rect 11624 14804 11652 14912
rect 11698 14900 11704 14952
rect 11756 14900 11762 14952
rect 11974 14900 11980 14952
rect 12032 14940 12038 14952
rect 12245 14940 12257 14953
rect 12032 14919 12257 14940
rect 12291 14919 12303 14953
rect 12032 14913 12303 14919
rect 12032 14912 12296 14913
rect 12032 14900 12038 14912
rect 12342 14900 12348 14952
rect 12400 14900 12406 14952
rect 12544 14949 12572 14980
rect 14277 14977 14289 14980
rect 14323 14977 14335 15011
rect 15565 15011 15623 15017
rect 15565 15008 15577 15011
rect 14277 14971 14335 14977
rect 14568 14980 15577 15008
rect 12529 14943 12587 14949
rect 12529 14909 12541 14943
rect 12575 14909 12587 14943
rect 12529 14903 12587 14909
rect 12621 14943 12679 14949
rect 12621 14909 12633 14943
rect 12667 14940 12679 14943
rect 12667 14912 14044 14940
rect 12667 14909 12679 14912
rect 12621 14903 12679 14909
rect 13814 14832 13820 14884
rect 13872 14832 13878 14884
rect 14016 14816 14044 14912
rect 14090 14900 14096 14952
rect 14148 14940 14154 14952
rect 14568 14949 14596 14980
rect 15565 14977 15577 14980
rect 15611 14977 15623 15011
rect 15565 14971 15623 14977
rect 14553 14943 14611 14949
rect 14553 14940 14565 14943
rect 14148 14912 14565 14940
rect 14148 14900 14154 14912
rect 14553 14909 14565 14912
rect 14599 14909 14611 14943
rect 14553 14903 14611 14909
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14909 14703 14943
rect 14645 14903 14703 14909
rect 14737 14943 14795 14949
rect 14737 14909 14749 14943
rect 14783 14940 14795 14943
rect 14826 14940 14832 14952
rect 14783 14912 14832 14940
rect 14783 14909 14795 14912
rect 14737 14903 14795 14909
rect 14660 14872 14688 14903
rect 14826 14900 14832 14912
rect 14884 14900 14890 14952
rect 14921 14943 14979 14949
rect 14921 14909 14933 14943
rect 14967 14940 14979 14943
rect 15010 14940 15016 14952
rect 14967 14912 15016 14940
rect 14967 14909 14979 14912
rect 14921 14903 14979 14909
rect 15010 14900 15016 14912
rect 15068 14900 15074 14952
rect 15654 14900 15660 14952
rect 15712 14900 15718 14952
rect 15948 14940 15976 15048
rect 16025 15045 16037 15079
rect 16071 15076 16083 15079
rect 17218 15076 17224 15088
rect 16071 15048 17224 15076
rect 16071 15045 16083 15048
rect 16025 15039 16083 15045
rect 17218 15036 17224 15048
rect 17276 15036 17282 15088
rect 18782 15076 18788 15088
rect 18248 15048 18788 15076
rect 18248 14949 18276 15048
rect 18782 15036 18788 15048
rect 18840 15076 18846 15088
rect 18840 15048 19012 15076
rect 18840 15036 18846 15048
rect 18322 14968 18328 15020
rect 18380 15008 18386 15020
rect 18877 15011 18935 15017
rect 18877 15008 18889 15011
rect 18380 14980 18889 15008
rect 18380 14968 18386 14980
rect 18877 14977 18889 14980
rect 18923 14977 18935 15011
rect 18877 14971 18935 14977
rect 18233 14943 18291 14949
rect 18233 14940 18245 14943
rect 15948 14912 18245 14940
rect 18233 14909 18245 14912
rect 18279 14909 18291 14943
rect 18233 14903 18291 14909
rect 16114 14872 16120 14884
rect 14660 14844 16120 14872
rect 16114 14832 16120 14844
rect 16172 14872 16178 14884
rect 17034 14872 17040 14884
rect 16172 14844 17040 14872
rect 16172 14832 16178 14844
rect 17034 14832 17040 14844
rect 17092 14832 17098 14884
rect 18892 14872 18920 14971
rect 18984 14949 19012 15048
rect 20254 15036 20260 15088
rect 20312 15076 20318 15088
rect 21545 15079 21603 15085
rect 20312 15048 21404 15076
rect 20312 15036 20318 15048
rect 19797 15011 19855 15017
rect 19797 14977 19809 15011
rect 19843 15008 19855 15011
rect 20533 15011 20591 15017
rect 20533 15008 20545 15011
rect 19843 14980 20545 15008
rect 19843 14977 19855 14980
rect 19797 14971 19855 14977
rect 20533 14977 20545 14980
rect 20579 15008 20591 15011
rect 20622 15008 20628 15020
rect 20579 14980 20628 15008
rect 20579 14977 20591 14980
rect 20533 14971 20591 14977
rect 20622 14968 20628 14980
rect 20680 14968 20686 15020
rect 20732 14980 21312 15008
rect 18969 14943 19027 14949
rect 18969 14909 18981 14943
rect 19015 14940 19027 14943
rect 19889 14943 19947 14949
rect 19889 14940 19901 14943
rect 19015 14912 19901 14940
rect 19015 14909 19027 14912
rect 18969 14903 19027 14909
rect 19889 14909 19901 14912
rect 19935 14909 19947 14943
rect 19889 14903 19947 14909
rect 20073 14943 20131 14949
rect 20073 14909 20085 14943
rect 20119 14909 20131 14943
rect 20073 14903 20131 14909
rect 20088 14872 20116 14903
rect 20438 14900 20444 14952
rect 20496 14900 20502 14952
rect 20732 14940 20760 14980
rect 20548 14912 20760 14940
rect 20548 14872 20576 14912
rect 20990 14900 20996 14952
rect 21048 14900 21054 14952
rect 21177 14943 21235 14949
rect 21177 14940 21189 14943
rect 21100 14912 21189 14940
rect 18892 14844 20576 14872
rect 20622 14832 20628 14884
rect 20680 14872 20686 14884
rect 21008 14872 21036 14900
rect 20680 14844 21036 14872
rect 20680 14832 20686 14844
rect 11698 14804 11704 14816
rect 11624 14776 11704 14804
rect 11698 14764 11704 14776
rect 11756 14764 11762 14816
rect 13906 14764 13912 14816
rect 13964 14764 13970 14816
rect 13998 14764 14004 14816
rect 14056 14764 14062 14816
rect 14182 14764 14188 14816
rect 14240 14804 14246 14816
rect 18322 14804 18328 14816
rect 14240 14776 18328 14804
rect 14240 14764 14246 14776
rect 18322 14764 18328 14776
rect 18380 14764 18386 14816
rect 20809 14807 20867 14813
rect 20809 14773 20821 14807
rect 20855 14804 20867 14807
rect 21100 14804 21128 14912
rect 21177 14909 21189 14912
rect 21223 14909 21235 14943
rect 21177 14903 21235 14909
rect 21284 14881 21312 14980
rect 21376 14949 21404 15048
rect 21545 15045 21557 15079
rect 21591 15045 21603 15079
rect 21545 15039 21603 15045
rect 21361 14943 21419 14949
rect 21361 14909 21373 14943
rect 21407 14909 21419 14943
rect 21560 14940 21588 15039
rect 21821 14943 21879 14949
rect 21821 14940 21833 14943
rect 21560 14912 21833 14940
rect 21361 14903 21419 14909
rect 21821 14909 21833 14912
rect 21867 14909 21879 14943
rect 21821 14903 21879 14909
rect 21910 14900 21916 14952
rect 21968 14940 21974 14952
rect 22186 14940 22192 14952
rect 21968 14912 22192 14940
rect 21968 14900 21974 14912
rect 22186 14900 22192 14912
rect 22244 14900 22250 14952
rect 21269 14875 21327 14881
rect 21269 14841 21281 14875
rect 21315 14872 21327 14875
rect 21634 14872 21640 14884
rect 21315 14844 21640 14872
rect 21315 14841 21327 14844
rect 21269 14835 21327 14841
rect 21634 14832 21640 14844
rect 21692 14832 21698 14884
rect 20855 14776 21128 14804
rect 20855 14773 20867 14776
rect 20809 14767 20867 14773
rect 552 14714 28587 14736
rect 552 14662 7366 14714
rect 7418 14662 7430 14714
rect 7482 14662 7494 14714
rect 7546 14662 7558 14714
rect 7610 14662 7622 14714
rect 7674 14662 14335 14714
rect 14387 14662 14399 14714
rect 14451 14662 14463 14714
rect 14515 14662 14527 14714
rect 14579 14662 14591 14714
rect 14643 14662 21304 14714
rect 21356 14662 21368 14714
rect 21420 14662 21432 14714
rect 21484 14662 21496 14714
rect 21548 14662 21560 14714
rect 21612 14662 28273 14714
rect 28325 14662 28337 14714
rect 28389 14662 28401 14714
rect 28453 14662 28465 14714
rect 28517 14662 28529 14714
rect 28581 14662 28587 14714
rect 552 14640 28587 14662
rect 3142 14560 3148 14612
rect 3200 14560 3206 14612
rect 3418 14560 3424 14612
rect 3476 14560 3482 14612
rect 6270 14560 6276 14612
rect 6328 14560 6334 14612
rect 9858 14560 9864 14612
rect 9916 14560 9922 14612
rect 10594 14560 10600 14612
rect 10652 14560 10658 14612
rect 11330 14560 11336 14612
rect 11388 14600 11394 14612
rect 12342 14600 12348 14612
rect 11388 14572 12348 14600
rect 11388 14560 11394 14572
rect 12342 14560 12348 14572
rect 12400 14600 12406 14612
rect 12437 14603 12495 14609
rect 12437 14600 12449 14603
rect 12400 14572 12449 14600
rect 12400 14560 12406 14572
rect 12437 14569 12449 14572
rect 12483 14569 12495 14603
rect 12437 14563 12495 14569
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 13909 14603 13967 14609
rect 13909 14600 13921 14603
rect 13872 14572 13921 14600
rect 13872 14560 13878 14572
rect 13909 14569 13921 14572
rect 13955 14569 13967 14603
rect 13909 14563 13967 14569
rect 13998 14560 14004 14612
rect 14056 14600 14062 14612
rect 14277 14603 14335 14609
rect 14277 14600 14289 14603
rect 14056 14572 14289 14600
rect 14056 14560 14062 14572
rect 14277 14569 14289 14572
rect 14323 14569 14335 14603
rect 14277 14563 14335 14569
rect 15562 14560 15568 14612
rect 15620 14560 15626 14612
rect 16114 14560 16120 14612
rect 16172 14560 16178 14612
rect 17310 14560 17316 14612
rect 17368 14560 17374 14612
rect 3160 14473 3188 14560
rect 3436 14473 3464 14560
rect 5442 14492 5448 14544
rect 5500 14532 5506 14544
rect 9876 14532 9904 14560
rect 5500 14504 9904 14532
rect 5500 14492 5506 14504
rect 3145 14467 3203 14473
rect 3145 14433 3157 14467
rect 3191 14433 3203 14467
rect 3145 14427 3203 14433
rect 3329 14467 3387 14473
rect 3329 14433 3341 14467
rect 3375 14433 3387 14467
rect 3329 14427 3387 14433
rect 3421 14467 3479 14473
rect 3421 14433 3433 14467
rect 3467 14433 3479 14467
rect 3421 14427 3479 14433
rect 3234 14396 3240 14408
rect 3160 14368 3240 14396
rect 3160 14337 3188 14368
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 3145 14331 3203 14337
rect 3145 14297 3157 14331
rect 3191 14297 3203 14331
rect 3344 14328 3372 14427
rect 3436 14396 3464 14427
rect 3786 14424 3792 14476
rect 3844 14424 3850 14476
rect 5994 14424 6000 14476
rect 6052 14424 6058 14476
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14464 6239 14467
rect 6457 14467 6515 14473
rect 6457 14464 6469 14467
rect 6227 14436 6469 14464
rect 6227 14433 6239 14436
rect 6181 14427 6239 14433
rect 6457 14433 6469 14436
rect 6503 14433 6515 14467
rect 6457 14427 6515 14433
rect 7742 14424 7748 14476
rect 7800 14464 7806 14476
rect 8481 14467 8539 14473
rect 8481 14464 8493 14467
rect 7800 14436 8493 14464
rect 7800 14424 7806 14436
rect 8481 14433 8493 14436
rect 8527 14433 8539 14467
rect 8481 14427 8539 14433
rect 8662 14424 8668 14476
rect 8720 14424 8726 14476
rect 10612 14473 10640 14560
rect 10686 14492 10692 14544
rect 10744 14532 10750 14544
rect 11698 14532 11704 14544
rect 10744 14504 11704 14532
rect 10744 14492 10750 14504
rect 11698 14492 11704 14504
rect 11756 14492 11762 14544
rect 12802 14541 12808 14544
rect 12796 14495 12808 14541
rect 12860 14532 12866 14544
rect 15105 14535 15163 14541
rect 15105 14532 15117 14535
rect 12860 14504 12896 14532
rect 14108 14504 15117 14532
rect 12802 14492 12808 14495
rect 12860 14492 12866 14504
rect 14108 14476 14136 14504
rect 15105 14501 15117 14504
rect 15151 14532 15163 14535
rect 15717 14535 15775 14541
rect 15717 14532 15729 14535
rect 15151 14504 15729 14532
rect 15151 14501 15163 14504
rect 15105 14495 15163 14501
rect 15717 14501 15729 14504
rect 15763 14501 15775 14535
rect 15717 14495 15775 14501
rect 15933 14535 15991 14541
rect 15933 14501 15945 14535
rect 15979 14532 15991 14535
rect 18877 14535 18935 14541
rect 15979 14504 17080 14532
rect 15979 14501 15991 14504
rect 15933 14495 15991 14501
rect 11330 14473 11336 14476
rect 10600 14467 10658 14473
rect 10600 14433 10612 14467
rect 10646 14433 10658 14467
rect 10600 14427 10658 14433
rect 11324 14427 11336 14473
rect 11330 14424 11336 14427
rect 11388 14424 11394 14476
rect 14090 14424 14096 14476
rect 14148 14424 14154 14476
rect 14277 14467 14335 14473
rect 14277 14433 14289 14467
rect 14323 14464 14335 14467
rect 14734 14464 14740 14476
rect 14323 14436 14740 14464
rect 14323 14433 14335 14436
rect 14277 14427 14335 14433
rect 14734 14424 14740 14436
rect 14792 14424 14798 14476
rect 16500 14473 16528 14504
rect 14921 14467 14979 14473
rect 14921 14433 14933 14467
rect 14967 14433 14979 14467
rect 14921 14427 14979 14433
rect 16301 14467 16359 14473
rect 16301 14433 16313 14467
rect 16347 14464 16359 14467
rect 16485 14467 16543 14473
rect 16347 14436 16381 14464
rect 16347 14433 16359 14436
rect 16301 14427 16359 14433
rect 16485 14433 16497 14467
rect 16531 14433 16543 14467
rect 16485 14427 16543 14433
rect 3697 14399 3755 14405
rect 3697 14396 3709 14399
rect 3436 14368 3709 14396
rect 3697 14365 3709 14368
rect 3743 14365 3755 14399
rect 3697 14359 3755 14365
rect 3804 14328 3832 14424
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14396 4215 14399
rect 4614 14396 4620 14408
rect 4203 14368 4620 14396
rect 4203 14365 4215 14368
rect 4157 14359 4215 14365
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 5810 14356 5816 14408
rect 5868 14356 5874 14408
rect 8110 14356 8116 14408
rect 8168 14396 8174 14408
rect 8680 14396 8708 14424
rect 8168 14368 8708 14396
rect 8168 14356 8174 14368
rect 8938 14356 8944 14408
rect 8996 14396 9002 14408
rect 9950 14396 9956 14408
rect 8996 14368 9956 14396
rect 8996 14356 9002 14368
rect 9950 14356 9956 14368
rect 10008 14356 10014 14408
rect 10413 14399 10471 14405
rect 10413 14365 10425 14399
rect 10459 14396 10471 14399
rect 11057 14399 11115 14405
rect 10459 14368 10548 14396
rect 10459 14365 10471 14368
rect 10413 14359 10471 14365
rect 3344 14300 3832 14328
rect 3145 14291 3203 14297
rect 5828 14260 5856 14356
rect 8665 14331 8723 14337
rect 8665 14297 8677 14331
rect 8711 14328 8723 14331
rect 9674 14328 9680 14340
rect 8711 14300 9680 14328
rect 8711 14297 8723 14300
rect 8665 14291 8723 14297
rect 9674 14288 9680 14300
rect 9732 14328 9738 14340
rect 10134 14328 10140 14340
rect 9732 14300 10140 14328
rect 9732 14288 9738 14300
rect 10134 14288 10140 14300
rect 10192 14288 10198 14340
rect 10520 14272 10548 14368
rect 11057 14365 11069 14399
rect 11103 14365 11115 14399
rect 12529 14399 12587 14405
rect 12529 14396 12541 14399
rect 11057 14359 11115 14365
rect 12406 14368 12541 14396
rect 10502 14260 10508 14272
rect 5828 14232 10508 14260
rect 10502 14220 10508 14232
rect 10560 14220 10566 14272
rect 10686 14220 10692 14272
rect 10744 14260 10750 14272
rect 10781 14263 10839 14269
rect 10781 14260 10793 14263
rect 10744 14232 10793 14260
rect 10744 14220 10750 14232
rect 10781 14229 10793 14232
rect 10827 14229 10839 14263
rect 11072 14260 11100 14359
rect 11238 14260 11244 14272
rect 11072 14232 11244 14260
rect 10781 14223 10839 14229
rect 11238 14220 11244 14232
rect 11296 14260 11302 14272
rect 12406 14260 12434 14368
rect 12529 14365 12541 14368
rect 12575 14365 12587 14399
rect 12529 14359 12587 14365
rect 13998 14356 14004 14408
rect 14056 14356 14062 14408
rect 14936 14396 14964 14427
rect 16316 14396 16344 14427
rect 16942 14424 16948 14476
rect 17000 14424 17006 14476
rect 17052 14464 17080 14504
rect 18877 14501 18889 14535
rect 18923 14532 18935 14535
rect 18966 14532 18972 14544
rect 18923 14504 18972 14532
rect 18923 14501 18935 14504
rect 18877 14495 18935 14501
rect 18966 14492 18972 14504
rect 19024 14492 19030 14544
rect 19058 14464 19064 14476
rect 17052 14436 19064 14464
rect 19058 14424 19064 14436
rect 19116 14424 19122 14476
rect 21453 14467 21511 14473
rect 21453 14433 21465 14467
rect 21499 14464 21511 14467
rect 21634 14464 21640 14476
rect 21499 14436 21640 14464
rect 21499 14433 21511 14436
rect 21453 14427 21511 14433
rect 21634 14424 21640 14436
rect 21692 14424 21698 14476
rect 16853 14399 16911 14405
rect 16853 14396 16865 14399
rect 14936 14368 16865 14396
rect 11296 14232 12434 14260
rect 14016 14260 14044 14356
rect 14185 14331 14243 14337
rect 14185 14297 14197 14331
rect 14231 14328 14243 14331
rect 14918 14328 14924 14340
rect 14231 14300 14924 14328
rect 14231 14297 14243 14300
rect 14185 14291 14243 14297
rect 14918 14288 14924 14300
rect 14976 14288 14982 14340
rect 15856 14272 15884 14368
rect 16853 14365 16865 14368
rect 16899 14365 16911 14399
rect 16853 14359 16911 14365
rect 18782 14288 18788 14340
rect 18840 14328 18846 14340
rect 19153 14331 19211 14337
rect 19153 14328 19165 14331
rect 18840 14300 19165 14328
rect 18840 14288 18846 14300
rect 19153 14297 19165 14300
rect 19199 14297 19211 14331
rect 19153 14291 19211 14297
rect 15010 14260 15016 14272
rect 14016 14232 15016 14260
rect 11296 14220 11302 14232
rect 15010 14220 15016 14232
rect 15068 14220 15074 14272
rect 15749 14263 15807 14269
rect 15749 14229 15761 14263
rect 15795 14260 15807 14263
rect 15838 14260 15844 14272
rect 15795 14232 15844 14260
rect 15795 14229 15807 14232
rect 15749 14223 15807 14229
rect 15838 14220 15844 14232
rect 15896 14220 15902 14272
rect 19334 14220 19340 14272
rect 19392 14220 19398 14272
rect 21637 14263 21695 14269
rect 21637 14229 21649 14263
rect 21683 14260 21695 14263
rect 22278 14260 22284 14272
rect 21683 14232 22284 14260
rect 21683 14229 21695 14232
rect 21637 14223 21695 14229
rect 22278 14220 22284 14232
rect 22336 14220 22342 14272
rect 552 14170 28428 14192
rect 552 14118 3882 14170
rect 3934 14118 3946 14170
rect 3998 14118 4010 14170
rect 4062 14118 4074 14170
rect 4126 14118 4138 14170
rect 4190 14118 10851 14170
rect 10903 14118 10915 14170
rect 10967 14118 10979 14170
rect 11031 14118 11043 14170
rect 11095 14118 11107 14170
rect 11159 14118 17820 14170
rect 17872 14118 17884 14170
rect 17936 14118 17948 14170
rect 18000 14118 18012 14170
rect 18064 14118 18076 14170
rect 18128 14118 24789 14170
rect 24841 14118 24853 14170
rect 24905 14118 24917 14170
rect 24969 14118 24981 14170
rect 25033 14118 25045 14170
rect 25097 14118 28428 14170
rect 552 14096 28428 14118
rect 5994 14016 6000 14068
rect 6052 14016 6058 14068
rect 7742 14056 7748 14068
rect 6840 14028 7748 14056
rect 6840 13929 6868 14028
rect 7484 13997 7512 14028
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 8938 14016 8944 14068
rect 8996 14016 9002 14068
rect 11330 14016 11336 14068
rect 11388 14056 11394 14068
rect 11425 14059 11483 14065
rect 11425 14056 11437 14059
rect 11388 14028 11437 14056
rect 11388 14016 11394 14028
rect 11425 14025 11437 14028
rect 11471 14025 11483 14059
rect 11425 14019 11483 14025
rect 19334 14016 19340 14068
rect 19392 14016 19398 14068
rect 7101 13991 7159 13997
rect 7101 13957 7113 13991
rect 7147 13988 7159 13991
rect 7469 13991 7527 13997
rect 7147 13960 7420 13988
rect 7147 13957 7159 13960
rect 7101 13951 7159 13957
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 5736 13892 6837 13920
rect 5736 13864 5764 13892
rect 6825 13889 6837 13892
rect 6871 13889 6883 13923
rect 7392 13920 7420 13960
rect 7469 13957 7481 13991
rect 7515 13957 7527 13991
rect 8956 13988 8984 14016
rect 7469 13951 7527 13957
rect 7576 13960 8984 13988
rect 7576 13920 7604 13960
rect 7392 13892 7604 13920
rect 6825 13883 6883 13889
rect 2038 13812 2044 13864
rect 2096 13812 2102 13864
rect 3973 13855 4031 13861
rect 3973 13821 3985 13855
rect 4019 13821 4031 13855
rect 3973 13815 4031 13821
rect 3234 13744 3240 13796
rect 3292 13784 3298 13796
rect 3988 13784 4016 13815
rect 4062 13812 4068 13864
rect 4120 13852 4126 13864
rect 4157 13855 4215 13861
rect 4157 13852 4169 13855
rect 4120 13824 4169 13852
rect 4120 13812 4126 13824
rect 4157 13821 4169 13824
rect 4203 13852 4215 13855
rect 4522 13852 4528 13864
rect 4203 13824 4528 13852
rect 4203 13821 4215 13824
rect 4157 13815 4215 13821
rect 4522 13812 4528 13824
rect 4580 13812 4586 13864
rect 4798 13812 4804 13864
rect 4856 13852 4862 13864
rect 5445 13855 5503 13861
rect 5445 13852 5457 13855
rect 4856 13824 5457 13852
rect 4856 13812 4862 13824
rect 5445 13821 5457 13824
rect 5491 13821 5503 13855
rect 5445 13815 5503 13821
rect 5718 13812 5724 13864
rect 5776 13812 5782 13864
rect 7852 13861 7880 13960
rect 10502 13948 10508 14000
rect 10560 13988 10566 14000
rect 10560 13960 12434 13988
rect 10560 13948 10566 13960
rect 11422 13920 11428 13932
rect 7944 13892 11428 13920
rect 5813 13855 5871 13861
rect 5813 13821 5825 13855
rect 5859 13852 5871 13855
rect 7837 13855 7895 13861
rect 5859 13824 7788 13852
rect 5859 13821 5871 13824
rect 5813 13815 5871 13821
rect 5074 13784 5080 13796
rect 3292 13756 5080 13784
rect 3292 13744 3298 13756
rect 5074 13744 5080 13756
rect 5132 13744 5138 13796
rect 5626 13744 5632 13796
rect 5684 13744 5690 13796
rect 1762 13676 1768 13728
rect 1820 13716 1826 13728
rect 1857 13719 1915 13725
rect 1857 13716 1869 13719
rect 1820 13688 1869 13716
rect 1820 13676 1826 13688
rect 1857 13685 1869 13688
rect 1903 13685 1915 13719
rect 1857 13679 1915 13685
rect 4154 13676 4160 13728
rect 4212 13676 4218 13728
rect 4522 13676 4528 13728
rect 4580 13716 4586 13728
rect 4706 13716 4712 13728
rect 4580 13688 4712 13716
rect 4580 13676 4586 13688
rect 4706 13676 4712 13688
rect 4764 13716 4770 13728
rect 5828 13716 5856 13815
rect 7190 13744 7196 13796
rect 7248 13784 7254 13796
rect 7760 13784 7788 13824
rect 7837 13821 7849 13855
rect 7883 13821 7895 13855
rect 7837 13815 7895 13821
rect 7944 13784 7972 13892
rect 11422 13880 11428 13892
rect 11480 13880 11486 13932
rect 12406 13920 12434 13960
rect 17218 13920 17224 13932
rect 12406 13892 17224 13920
rect 17218 13880 17224 13892
rect 17276 13880 17282 13932
rect 18966 13880 18972 13932
rect 19024 13920 19030 13932
rect 19153 13923 19211 13929
rect 19153 13920 19165 13923
rect 19024 13892 19165 13920
rect 19024 13880 19030 13892
rect 19153 13889 19165 13892
rect 19199 13889 19211 13923
rect 19153 13883 19211 13889
rect 8849 13855 8907 13861
rect 8849 13821 8861 13855
rect 8895 13852 8907 13855
rect 9858 13852 9864 13864
rect 8895 13824 9864 13852
rect 8895 13821 8907 13824
rect 8849 13815 8907 13821
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 10686 13812 10692 13864
rect 10744 13852 10750 13864
rect 11609 13855 11667 13861
rect 11609 13852 11621 13855
rect 10744 13824 11621 13852
rect 10744 13812 10750 13824
rect 11609 13821 11621 13824
rect 11655 13821 11667 13855
rect 11609 13815 11667 13821
rect 13630 13812 13636 13864
rect 13688 13812 13694 13864
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 18322 13812 18328 13864
rect 18380 13852 18386 13864
rect 18877 13855 18935 13861
rect 18877 13852 18889 13855
rect 18380 13824 18889 13852
rect 18380 13812 18386 13824
rect 18877 13821 18889 13824
rect 18923 13821 18935 13855
rect 18877 13815 18935 13821
rect 19058 13812 19064 13864
rect 19116 13812 19122 13864
rect 7248 13756 7420 13784
rect 7760 13756 7972 13784
rect 19168 13784 19196 13883
rect 19352 13861 19380 14016
rect 21177 13991 21235 13997
rect 21177 13988 21189 13991
rect 20824 13960 21189 13988
rect 19797 13923 19855 13929
rect 19797 13920 19809 13923
rect 19444 13892 19809 13920
rect 19444 13864 19472 13892
rect 19797 13889 19809 13892
rect 19843 13889 19855 13923
rect 19797 13883 19855 13889
rect 20257 13923 20315 13929
rect 20257 13889 20269 13923
rect 20303 13920 20315 13923
rect 20303 13892 20760 13920
rect 20303 13889 20315 13892
rect 20257 13883 20315 13889
rect 19337 13855 19395 13861
rect 19337 13821 19349 13855
rect 19383 13821 19395 13855
rect 19337 13815 19395 13821
rect 19426 13812 19432 13864
rect 19484 13812 19490 13864
rect 19518 13812 19524 13864
rect 19576 13812 19582 13864
rect 19886 13812 19892 13864
rect 19944 13852 19950 13864
rect 20346 13852 20352 13864
rect 19944 13824 20352 13852
rect 19944 13812 19950 13824
rect 20346 13812 20352 13824
rect 20404 13812 20410 13864
rect 20533 13855 20591 13861
rect 20533 13821 20545 13855
rect 20579 13852 20591 13855
rect 20622 13852 20628 13864
rect 20579 13824 20628 13852
rect 20579 13821 20591 13824
rect 20533 13815 20591 13821
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 20732 13861 20760 13892
rect 20824 13861 20852 13960
rect 21177 13957 21189 13960
rect 21223 13957 21235 13991
rect 21177 13951 21235 13957
rect 20717 13855 20775 13861
rect 20717 13821 20729 13855
rect 20763 13821 20775 13855
rect 20717 13815 20775 13821
rect 20809 13855 20867 13861
rect 20809 13821 20821 13855
rect 20855 13821 20867 13855
rect 20809 13815 20867 13821
rect 20901 13855 20959 13861
rect 20901 13821 20913 13855
rect 20947 13821 20959 13855
rect 22557 13855 22615 13861
rect 22557 13852 22569 13855
rect 20901 13815 20959 13821
rect 22112 13824 22569 13852
rect 20824 13784 20852 13815
rect 19168 13756 20852 13784
rect 7248 13744 7254 13756
rect 4764 13688 5856 13716
rect 4764 13676 4770 13688
rect 7282 13676 7288 13728
rect 7340 13676 7346 13728
rect 7392 13725 7420 13756
rect 7377 13719 7435 13725
rect 7377 13685 7389 13719
rect 7423 13685 7435 13719
rect 7377 13679 7435 13685
rect 7742 13676 7748 13728
rect 7800 13716 7806 13728
rect 13446 13716 13452 13728
rect 7800 13688 13452 13716
rect 7800 13676 7806 13688
rect 13446 13676 13452 13688
rect 13504 13676 13510 13728
rect 13722 13676 13728 13728
rect 13780 13676 13786 13728
rect 18693 13719 18751 13725
rect 18693 13685 18705 13719
rect 18739 13716 18751 13719
rect 18874 13716 18880 13728
rect 18739 13688 18880 13716
rect 18739 13685 18751 13688
rect 18693 13679 18751 13685
rect 18874 13676 18880 13688
rect 18932 13676 18938 13728
rect 19426 13676 19432 13728
rect 19484 13676 19490 13728
rect 19978 13676 19984 13728
rect 20036 13716 20042 13728
rect 20254 13716 20260 13728
rect 20036 13688 20260 13716
rect 20036 13676 20042 13688
rect 20254 13676 20260 13688
rect 20312 13716 20318 13728
rect 20916 13716 20944 13815
rect 22002 13744 22008 13796
rect 22060 13784 22066 13796
rect 22112 13784 22140 13824
rect 22557 13821 22569 13824
rect 22603 13821 22615 13855
rect 22557 13815 22615 13821
rect 22060 13756 22140 13784
rect 22060 13744 22066 13756
rect 22278 13744 22284 13796
rect 22336 13793 22342 13796
rect 22336 13747 22348 13793
rect 22336 13744 22342 13747
rect 20312 13688 20944 13716
rect 20312 13676 20318 13688
rect 21082 13676 21088 13728
rect 21140 13676 21146 13728
rect 552 13626 28587 13648
rect 552 13574 7366 13626
rect 7418 13574 7430 13626
rect 7482 13574 7494 13626
rect 7546 13574 7558 13626
rect 7610 13574 7622 13626
rect 7674 13574 14335 13626
rect 14387 13574 14399 13626
rect 14451 13574 14463 13626
rect 14515 13574 14527 13626
rect 14579 13574 14591 13626
rect 14643 13574 21304 13626
rect 21356 13574 21368 13626
rect 21420 13574 21432 13626
rect 21484 13574 21496 13626
rect 21548 13574 21560 13626
rect 21612 13574 28273 13626
rect 28325 13574 28337 13626
rect 28389 13574 28401 13626
rect 28453 13574 28465 13626
rect 28517 13574 28529 13626
rect 28581 13574 28587 13626
rect 552 13552 28587 13574
rect 5902 13512 5908 13524
rect 2746 13484 5908 13512
rect 1578 13404 1584 13456
rect 1636 13444 1642 13456
rect 2746 13444 2774 13484
rect 5902 13472 5908 13484
rect 5960 13512 5966 13524
rect 6089 13515 6147 13521
rect 6089 13512 6101 13515
rect 5960 13484 6101 13512
rect 5960 13472 5966 13484
rect 6089 13481 6101 13484
rect 6135 13481 6147 13515
rect 7742 13512 7748 13524
rect 6089 13475 6147 13481
rect 7484 13484 7748 13512
rect 1636 13416 2774 13444
rect 1636 13404 1642 13416
rect 3050 13404 3056 13456
rect 3108 13444 3114 13456
rect 4062 13444 4068 13456
rect 3108 13416 4068 13444
rect 3108 13404 3114 13416
rect 1489 13379 1547 13385
rect 1489 13345 1501 13379
rect 1535 13376 1547 13379
rect 1596 13376 1624 13404
rect 1762 13385 1768 13388
rect 1756 13376 1768 13385
rect 1535 13348 1624 13376
rect 1723 13348 1768 13376
rect 1535 13345 1547 13348
rect 1489 13339 1547 13345
rect 1756 13339 1768 13348
rect 1762 13336 1768 13339
rect 1820 13336 1826 13388
rect 3160 13385 3188 13416
rect 4062 13404 4068 13416
rect 4120 13404 4126 13456
rect 4154 13404 4160 13456
rect 4212 13444 4218 13456
rect 4249 13447 4307 13453
rect 4249 13444 4261 13447
rect 4212 13416 4261 13444
rect 4212 13404 4218 13416
rect 4249 13413 4261 13416
rect 4295 13413 4307 13447
rect 4249 13407 4307 13413
rect 4617 13447 4675 13453
rect 4617 13413 4629 13447
rect 4663 13444 4675 13447
rect 5074 13444 5080 13456
rect 4663 13416 5080 13444
rect 4663 13413 4675 13416
rect 4617 13407 4675 13413
rect 5074 13404 5080 13416
rect 5132 13404 5138 13456
rect 3145 13379 3203 13385
rect 3145 13345 3157 13379
rect 3191 13345 3203 13379
rect 3881 13379 3939 13385
rect 3881 13376 3893 13379
rect 3145 13339 3203 13345
rect 3528 13348 3893 13376
rect 3234 13268 3240 13320
rect 3292 13268 3298 13320
rect 2869 13243 2927 13249
rect 2869 13209 2881 13243
rect 2915 13240 2927 13243
rect 3252 13240 3280 13268
rect 3528 13252 3556 13348
rect 3881 13345 3893 13348
rect 3927 13345 3939 13379
rect 3881 13339 3939 13345
rect 4522 13336 4528 13388
rect 4580 13336 4586 13388
rect 4706 13336 4712 13388
rect 4764 13336 4770 13388
rect 4890 13336 4896 13388
rect 4948 13376 4954 13388
rect 7484 13376 7512 13484
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 10045 13515 10103 13521
rect 10045 13481 10057 13515
rect 10091 13512 10103 13515
rect 10318 13512 10324 13524
rect 10091 13484 10324 13512
rect 10091 13481 10103 13484
rect 10045 13475 10103 13481
rect 10318 13472 10324 13484
rect 10376 13472 10382 13524
rect 10410 13472 10416 13524
rect 10468 13512 10474 13524
rect 10597 13515 10655 13521
rect 10597 13512 10609 13515
rect 10468 13484 10609 13512
rect 10468 13472 10474 13484
rect 10597 13481 10609 13484
rect 10643 13481 10655 13515
rect 10597 13475 10655 13481
rect 13449 13515 13507 13521
rect 13449 13481 13461 13515
rect 13495 13481 13507 13515
rect 13449 13475 13507 13481
rect 7561 13447 7619 13453
rect 7561 13413 7573 13447
rect 7607 13444 7619 13447
rect 7837 13447 7895 13453
rect 7837 13444 7849 13447
rect 7607 13416 7849 13444
rect 7607 13413 7619 13416
rect 7561 13407 7619 13413
rect 7837 13413 7849 13416
rect 7883 13444 7895 13447
rect 8202 13444 8208 13456
rect 7883 13416 8208 13444
rect 7883 13413 7895 13416
rect 7837 13407 7895 13413
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 9585 13447 9643 13453
rect 9585 13413 9597 13447
rect 9631 13444 9643 13447
rect 11238 13444 11244 13456
rect 9631 13416 11244 13444
rect 9631 13413 9643 13416
rect 9585 13407 9643 13413
rect 11238 13404 11244 13416
rect 11296 13404 11302 13456
rect 11422 13404 11428 13456
rect 11480 13404 11486 13456
rect 13464 13444 13492 13475
rect 14182 13472 14188 13524
rect 14240 13512 14246 13524
rect 15749 13515 15807 13521
rect 14240 13484 14872 13512
rect 14240 13472 14246 13484
rect 13630 13444 13636 13456
rect 13464 13416 13636 13444
rect 13630 13404 13636 13416
rect 13688 13444 13694 13456
rect 13725 13447 13783 13453
rect 13725 13444 13737 13447
rect 13688 13416 13737 13444
rect 13688 13404 13694 13416
rect 13725 13413 13737 13416
rect 13771 13413 13783 13447
rect 13725 13407 13783 13413
rect 13814 13404 13820 13456
rect 13872 13444 13878 13456
rect 13909 13447 13967 13453
rect 13909 13444 13921 13447
rect 13872 13416 13921 13444
rect 13872 13404 13878 13416
rect 13909 13413 13921 13416
rect 13955 13444 13967 13447
rect 14093 13447 14151 13453
rect 14093 13444 14105 13447
rect 13955 13416 14105 13444
rect 13955 13413 13967 13416
rect 13909 13407 13967 13413
rect 14093 13413 14105 13416
rect 14139 13413 14151 13447
rect 14093 13407 14151 13413
rect 14599 13447 14657 13453
rect 14599 13413 14611 13447
rect 14645 13444 14657 13447
rect 14734 13444 14740 13456
rect 14645 13416 14740 13444
rect 14645 13413 14657 13416
rect 14599 13407 14657 13413
rect 14734 13404 14740 13416
rect 14792 13404 14798 13456
rect 4948 13348 7512 13376
rect 4948 13336 4954 13348
rect 9858 13336 9864 13388
rect 9916 13336 9922 13388
rect 10134 13336 10140 13388
rect 10192 13336 10198 13388
rect 10229 13379 10287 13385
rect 10229 13345 10241 13379
rect 10275 13345 10287 13379
rect 10229 13339 10287 13345
rect 13081 13379 13139 13385
rect 13081 13345 13093 13379
rect 13127 13376 13139 13379
rect 13127 13348 14136 13376
rect 13127 13345 13139 13348
rect 13081 13339 13139 13345
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13308 4123 13311
rect 4614 13308 4620 13320
rect 4111 13280 4620 13308
rect 4111 13277 4123 13280
rect 4065 13271 4123 13277
rect 4614 13268 4620 13280
rect 4672 13268 4678 13320
rect 9030 13268 9036 13320
rect 9088 13308 9094 13320
rect 9398 13308 9404 13320
rect 9088 13280 9404 13308
rect 9088 13268 9094 13280
rect 9398 13268 9404 13280
rect 9456 13308 9462 13320
rect 10244 13308 10272 13339
rect 9456 13280 10272 13308
rect 9456 13268 9462 13280
rect 10318 13268 10324 13320
rect 10376 13268 10382 13320
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13308 13047 13311
rect 13998 13308 14004 13320
rect 13035 13280 14004 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 2915 13212 3280 13240
rect 2915 13209 2927 13212
rect 2869 13203 2927 13209
rect 3510 13200 3516 13252
rect 3568 13200 3574 13252
rect 3786 13200 3792 13252
rect 3844 13240 3850 13252
rect 3881 13243 3939 13249
rect 3881 13240 3893 13243
rect 3844 13212 3893 13240
rect 3844 13200 3850 13212
rect 3881 13209 3893 13212
rect 3927 13209 3939 13243
rect 3881 13203 3939 13209
rect 13004 13184 13032 13271
rect 13998 13268 14004 13280
rect 14056 13268 14062 13320
rect 13906 13200 13912 13252
rect 13964 13240 13970 13252
rect 14108 13240 14136 13348
rect 14182 13336 14188 13388
rect 14240 13376 14246 13388
rect 14277 13379 14335 13385
rect 14277 13376 14289 13379
rect 14240 13348 14289 13376
rect 14240 13336 14246 13348
rect 14277 13345 14289 13348
rect 14323 13345 14335 13379
rect 14277 13339 14335 13345
rect 14366 13336 14372 13388
rect 14424 13336 14430 13388
rect 14461 13379 14519 13385
rect 14461 13345 14473 13379
rect 14507 13345 14519 13379
rect 14461 13339 14519 13345
rect 14844 13376 14872 13484
rect 15749 13481 15761 13515
rect 15795 13512 15807 13515
rect 16298 13512 16304 13524
rect 15795 13484 16304 13512
rect 15795 13481 15807 13484
rect 15749 13475 15807 13481
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 19334 13512 19340 13524
rect 18616 13484 19340 13512
rect 15212 13416 15516 13444
rect 15212 13388 15240 13416
rect 15194 13376 15200 13388
rect 14844 13348 15200 13376
rect 13964 13212 14136 13240
rect 13964 13200 13970 13212
rect 3418 13132 3424 13184
rect 3476 13172 3482 13184
rect 4341 13175 4399 13181
rect 4341 13172 4353 13175
rect 3476 13144 4353 13172
rect 3476 13132 3482 13144
rect 4341 13141 4353 13144
rect 4387 13141 4399 13175
rect 4341 13135 4399 13141
rect 9674 13132 9680 13184
rect 9732 13132 9738 13184
rect 10410 13132 10416 13184
rect 10468 13132 10474 13184
rect 11698 13132 11704 13184
rect 11756 13172 11762 13184
rect 12894 13172 12900 13184
rect 11756 13144 12900 13172
rect 11756 13132 11762 13144
rect 12894 13132 12900 13144
rect 12952 13132 12958 13184
rect 12986 13132 12992 13184
rect 13044 13132 13050 13184
rect 13538 13132 13544 13184
rect 13596 13132 13602 13184
rect 14476 13172 14504 13339
rect 14737 13311 14795 13317
rect 14737 13277 14749 13311
rect 14783 13308 14795 13311
rect 14844 13308 14872 13348
rect 15194 13336 15200 13348
rect 15252 13336 15258 13388
rect 15381 13379 15439 13385
rect 15381 13345 15393 13379
rect 15427 13345 15439 13379
rect 15488 13376 15516 13416
rect 15562 13404 15568 13456
rect 15620 13444 15626 13456
rect 15620 13416 16160 13444
rect 15620 13404 15626 13416
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15488 13348 15669 13376
rect 15381 13339 15439 13345
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 14783 13280 14872 13308
rect 15396 13308 15424 13339
rect 15838 13336 15844 13388
rect 15896 13336 15902 13388
rect 16132 13385 16160 13416
rect 16224 13416 17632 13444
rect 16224 13388 16252 13416
rect 16117 13379 16175 13385
rect 16117 13345 16129 13379
rect 16163 13345 16175 13379
rect 16117 13339 16175 13345
rect 16206 13336 16212 13388
rect 16264 13336 16270 13388
rect 16298 13336 16304 13388
rect 16356 13336 16362 13388
rect 17604 13376 17632 13416
rect 17678 13404 17684 13456
rect 17736 13444 17742 13456
rect 17782 13447 17840 13453
rect 17782 13444 17794 13447
rect 17736 13416 17794 13444
rect 17736 13404 17742 13416
rect 17782 13413 17794 13416
rect 17828 13413 17840 13447
rect 17782 13407 17840 13413
rect 18616 13376 18644 13484
rect 19334 13472 19340 13484
rect 19392 13472 19398 13524
rect 19518 13472 19524 13524
rect 19576 13472 19582 13524
rect 19797 13515 19855 13521
rect 19797 13481 19809 13515
rect 19843 13512 19855 13515
rect 19886 13512 19892 13524
rect 19843 13484 19892 13512
rect 19843 13481 19855 13484
rect 19797 13475 19855 13481
rect 19886 13472 19892 13484
rect 19944 13472 19950 13524
rect 21082 13472 21088 13524
rect 21140 13472 21146 13524
rect 21634 13472 21640 13524
rect 21692 13472 21698 13524
rect 18782 13404 18788 13456
rect 18840 13444 18846 13456
rect 19061 13447 19119 13453
rect 19061 13444 19073 13447
rect 18840 13416 19073 13444
rect 18840 13404 18846 13416
rect 19061 13413 19073 13416
rect 19107 13413 19119 13447
rect 19536 13444 19564 13472
rect 19613 13447 19671 13453
rect 19613 13444 19625 13447
rect 19536 13416 19625 13444
rect 19061 13407 19119 13413
rect 19613 13413 19625 13416
rect 19659 13413 19671 13447
rect 19904 13444 19932 13472
rect 19904 13416 20024 13444
rect 19613 13407 19671 13413
rect 17604 13348 18644 13376
rect 18693 13379 18751 13385
rect 18693 13345 18705 13379
rect 18739 13376 18751 13379
rect 19426 13376 19432 13388
rect 18739 13348 19432 13376
rect 18739 13345 18751 13348
rect 18693 13339 18751 13345
rect 19426 13336 19432 13348
rect 19484 13376 19490 13388
rect 19889 13379 19947 13385
rect 19889 13376 19901 13379
rect 19484 13348 19901 13376
rect 19484 13336 19490 13348
rect 19889 13345 19901 13348
rect 19935 13345 19947 13379
rect 19889 13339 19947 13345
rect 15856 13308 15884 13336
rect 15396 13280 16712 13308
rect 14783 13277 14795 13280
rect 14737 13271 14795 13277
rect 14550 13200 14556 13252
rect 14608 13240 14614 13252
rect 14608 13212 16160 13240
rect 14608 13200 14614 13212
rect 16132 13184 16160 13212
rect 14826 13172 14832 13184
rect 14476 13144 14832 13172
rect 14826 13132 14832 13144
rect 14884 13132 14890 13184
rect 15010 13132 15016 13184
rect 15068 13172 15074 13184
rect 15562 13172 15568 13184
rect 15068 13144 15568 13172
rect 15068 13132 15074 13144
rect 15562 13132 15568 13144
rect 15620 13132 15626 13184
rect 16114 13132 16120 13184
rect 16172 13132 16178 13184
rect 16684 13181 16712 13280
rect 18046 13268 18052 13320
rect 18104 13268 18110 13320
rect 18598 13268 18604 13320
rect 18656 13268 18662 13320
rect 18785 13311 18843 13317
rect 18785 13277 18797 13311
rect 18831 13277 18843 13311
rect 18785 13271 18843 13277
rect 16758 13200 16764 13252
rect 16816 13240 16822 13252
rect 16816 13212 17172 13240
rect 16816 13200 16822 13212
rect 16669 13175 16727 13181
rect 16669 13141 16681 13175
rect 16715 13172 16727 13175
rect 17034 13172 17040 13184
rect 16715 13144 17040 13172
rect 16715 13141 16727 13144
rect 16669 13135 16727 13141
rect 17034 13132 17040 13144
rect 17092 13132 17098 13184
rect 17144 13172 17172 13212
rect 18417 13175 18475 13181
rect 18417 13172 18429 13175
rect 17144 13144 18429 13172
rect 18417 13141 18429 13144
rect 18463 13141 18475 13175
rect 18800 13172 18828 13271
rect 18874 13268 18880 13320
rect 18932 13268 18938 13320
rect 18966 13200 18972 13252
rect 19024 13240 19030 13252
rect 19337 13243 19395 13249
rect 19337 13240 19349 13243
rect 19024 13212 19349 13240
rect 19024 13200 19030 13212
rect 19337 13209 19349 13212
rect 19383 13209 19395 13243
rect 19996 13240 20024 13416
rect 21100 13376 21128 13472
rect 21453 13379 21511 13385
rect 21453 13376 21465 13379
rect 21100 13348 21465 13376
rect 21453 13345 21465 13348
rect 21499 13345 21511 13379
rect 21453 13339 21511 13345
rect 20346 13268 20352 13320
rect 20404 13308 20410 13320
rect 21269 13311 21327 13317
rect 21269 13308 21281 13311
rect 20404 13280 21281 13308
rect 20404 13268 20410 13280
rect 21269 13277 21281 13280
rect 21315 13308 21327 13311
rect 21910 13308 21916 13320
rect 21315 13280 21916 13308
rect 21315 13277 21327 13280
rect 21269 13271 21327 13277
rect 21910 13268 21916 13280
rect 21968 13268 21974 13320
rect 19337 13203 19395 13209
rect 19444 13212 20024 13240
rect 19444 13172 19472 13212
rect 18800 13144 19472 13172
rect 18417 13135 18475 13141
rect 19610 13132 19616 13184
rect 19668 13132 19674 13184
rect 552 13082 28428 13104
rect 552 13030 3882 13082
rect 3934 13030 3946 13082
rect 3998 13030 4010 13082
rect 4062 13030 4074 13082
rect 4126 13030 4138 13082
rect 4190 13030 10851 13082
rect 10903 13030 10915 13082
rect 10967 13030 10979 13082
rect 11031 13030 11043 13082
rect 11095 13030 11107 13082
rect 11159 13030 17820 13082
rect 17872 13030 17884 13082
rect 17936 13030 17948 13082
rect 18000 13030 18012 13082
rect 18064 13030 18076 13082
rect 18128 13030 24789 13082
rect 24841 13030 24853 13082
rect 24905 13030 24917 13082
rect 24969 13030 24981 13082
rect 25033 13030 25045 13082
rect 25097 13030 28428 13082
rect 552 13008 28428 13030
rect 2038 12928 2044 12980
rect 2096 12928 2102 12980
rect 3418 12968 3424 12980
rect 2746 12940 3424 12968
rect 2746 12832 2774 12940
rect 3418 12928 3424 12940
rect 3476 12928 3482 12980
rect 3510 12928 3516 12980
rect 3568 12928 3574 12980
rect 4706 12968 4712 12980
rect 4172 12940 4712 12968
rect 2240 12804 2774 12832
rect 3528 12832 3556 12928
rect 4172 12909 4200 12940
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 5626 12928 5632 12980
rect 5684 12968 5690 12980
rect 5813 12971 5871 12977
rect 5813 12968 5825 12971
rect 5684 12940 5825 12968
rect 5684 12928 5690 12940
rect 5813 12937 5825 12940
rect 5859 12937 5871 12971
rect 5813 12931 5871 12937
rect 7653 12971 7711 12977
rect 7653 12937 7665 12971
rect 7699 12968 7711 12971
rect 7742 12968 7748 12980
rect 7699 12940 7748 12968
rect 7699 12937 7711 12940
rect 7653 12931 7711 12937
rect 7742 12928 7748 12940
rect 7800 12928 7806 12980
rect 7837 12971 7895 12977
rect 7837 12937 7849 12971
rect 7883 12968 7895 12971
rect 7883 12940 8984 12968
rect 7883 12937 7895 12940
rect 7837 12931 7895 12937
rect 4157 12903 4215 12909
rect 4157 12869 4169 12903
rect 4203 12869 4215 12903
rect 7929 12903 7987 12909
rect 7929 12900 7941 12903
rect 4157 12863 4215 12869
rect 6656 12872 7941 12900
rect 3697 12835 3755 12841
rect 3697 12832 3709 12835
rect 3528 12804 3709 12832
rect 2240 12773 2268 12804
rect 3697 12801 3709 12804
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 6273 12835 6331 12841
rect 6273 12801 6285 12835
rect 6319 12832 6331 12835
rect 6656 12832 6684 12872
rect 7929 12869 7941 12872
rect 7975 12869 7987 12903
rect 8956 12900 8984 12940
rect 9030 12928 9036 12980
rect 9088 12928 9094 12980
rect 9766 12928 9772 12980
rect 9824 12968 9830 12980
rect 10321 12971 10379 12977
rect 10321 12968 10333 12971
rect 9824 12940 10333 12968
rect 9824 12928 9830 12940
rect 10321 12937 10333 12940
rect 10367 12968 10379 12971
rect 10502 12968 10508 12980
rect 10367 12940 10508 12968
rect 10367 12937 10379 12940
rect 10321 12931 10379 12937
rect 10502 12928 10508 12940
rect 10560 12928 10566 12980
rect 10781 12971 10839 12977
rect 10781 12937 10793 12971
rect 10827 12937 10839 12971
rect 10781 12931 10839 12937
rect 10410 12900 10416 12912
rect 8956 12872 10416 12900
rect 7929 12863 7987 12869
rect 10410 12860 10416 12872
rect 10468 12900 10474 12912
rect 10796 12900 10824 12931
rect 11882 12928 11888 12980
rect 11940 12968 11946 12980
rect 12621 12971 12679 12977
rect 11940 12940 12296 12968
rect 11940 12928 11946 12940
rect 10468 12872 10824 12900
rect 10468 12860 10474 12872
rect 6319 12804 6684 12832
rect 6319 12801 6331 12804
rect 6273 12795 6331 12801
rect 2225 12767 2283 12773
rect 2225 12733 2237 12767
rect 2271 12733 2283 12767
rect 2225 12727 2283 12733
rect 2406 12724 2412 12776
rect 2464 12724 2470 12776
rect 3786 12724 3792 12776
rect 3844 12724 3850 12776
rect 6086 12724 6092 12776
rect 6144 12764 6150 12776
rect 6656 12773 6684 12804
rect 7190 12792 7196 12844
rect 7248 12832 7254 12844
rect 7469 12835 7527 12841
rect 7469 12832 7481 12835
rect 7248 12804 7481 12832
rect 7248 12792 7254 12804
rect 7469 12801 7481 12804
rect 7515 12832 7527 12835
rect 7515 12804 7972 12832
rect 7515 12801 7527 12804
rect 7469 12795 7527 12801
rect 6181 12767 6239 12773
rect 6181 12764 6193 12767
rect 6144 12736 6193 12764
rect 6144 12724 6150 12736
rect 6181 12733 6193 12736
rect 6227 12733 6239 12767
rect 6181 12727 6239 12733
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12733 6699 12767
rect 6641 12727 6699 12733
rect 6917 12767 6975 12773
rect 6917 12733 6929 12767
rect 6963 12764 6975 12767
rect 7208 12764 7236 12792
rect 6963 12736 7236 12764
rect 6963 12733 6975 12736
rect 6917 12727 6975 12733
rect 6196 12696 6224 12727
rect 7282 12724 7288 12776
rect 7340 12724 7346 12776
rect 7944 12773 7972 12804
rect 8754 12792 8760 12844
rect 8812 12792 8818 12844
rect 10045 12835 10103 12841
rect 10045 12801 10057 12835
rect 10091 12801 10103 12835
rect 10045 12795 10103 12801
rect 7653 12767 7711 12773
rect 7653 12733 7665 12767
rect 7699 12733 7711 12767
rect 7653 12727 7711 12733
rect 7929 12767 7987 12773
rect 7929 12733 7941 12767
rect 7975 12733 7987 12767
rect 7929 12727 7987 12733
rect 8113 12767 8171 12773
rect 8113 12733 8125 12767
rect 8159 12733 8171 12767
rect 8113 12727 8171 12733
rect 6733 12699 6791 12705
rect 6733 12696 6745 12699
rect 6196 12668 6745 12696
rect 6733 12665 6745 12668
rect 6779 12696 6791 12699
rect 7193 12699 7251 12705
rect 7193 12696 7205 12699
rect 6779 12668 7205 12696
rect 6779 12665 6791 12668
rect 6733 12659 6791 12665
rect 7193 12665 7205 12668
rect 7239 12665 7251 12699
rect 7300 12696 7328 12724
rect 7668 12696 7696 12727
rect 8128 12696 8156 12727
rect 8662 12724 8668 12776
rect 8720 12764 8726 12776
rect 8938 12764 8944 12776
rect 8720 12736 8944 12764
rect 8720 12724 8726 12736
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 9766 12724 9772 12776
rect 9824 12724 9830 12776
rect 9953 12767 10011 12773
rect 9953 12733 9965 12767
rect 9999 12764 10011 12767
rect 10060 12764 10088 12795
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 10778 12832 10784 12844
rect 10192 12804 10784 12832
rect 10192 12792 10198 12804
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 11238 12792 11244 12844
rect 11296 12792 11302 12844
rect 9999 12736 10088 12764
rect 9999 12733 10011 12736
rect 9953 12727 10011 12733
rect 10226 12724 10232 12776
rect 10284 12764 10290 12776
rect 10505 12767 10563 12773
rect 10505 12764 10517 12767
rect 10284 12736 10517 12764
rect 10284 12724 10290 12736
rect 10505 12733 10517 12736
rect 10551 12733 10563 12767
rect 10505 12727 10563 12733
rect 7300 12668 8156 12696
rect 7193 12659 7251 12665
rect 7098 12588 7104 12640
rect 7156 12588 7162 12640
rect 8956 12628 8984 12724
rect 9858 12656 9864 12708
rect 9916 12696 9922 12708
rect 10318 12696 10324 12708
rect 9916 12668 10324 12696
rect 9916 12656 9922 12668
rect 10318 12656 10324 12668
rect 10376 12696 10382 12708
rect 10965 12699 11023 12705
rect 10965 12696 10977 12699
rect 10376 12668 10977 12696
rect 10376 12656 10382 12668
rect 10965 12665 10977 12668
rect 11011 12665 11023 12699
rect 10965 12659 11023 12665
rect 11508 12699 11566 12705
rect 11508 12665 11520 12699
rect 11554 12696 11566 12699
rect 11882 12696 11888 12708
rect 11554 12668 11888 12696
rect 11554 12665 11566 12668
rect 11508 12659 11566 12665
rect 11882 12656 11888 12668
rect 11940 12656 11946 12708
rect 12268 12696 12296 12940
rect 12621 12937 12633 12971
rect 12667 12968 12679 12971
rect 12986 12968 12992 12980
rect 12667 12940 12992 12968
rect 12667 12937 12679 12940
rect 12621 12931 12679 12937
rect 12986 12928 12992 12940
rect 13044 12928 13050 12980
rect 13538 12928 13544 12980
rect 13596 12968 13602 12980
rect 13725 12971 13783 12977
rect 13725 12968 13737 12971
rect 13596 12940 13737 12968
rect 13596 12928 13602 12940
rect 13725 12937 13737 12940
rect 13771 12937 13783 12971
rect 15013 12971 15071 12977
rect 15013 12968 15025 12971
rect 13725 12931 13783 12937
rect 14936 12940 15025 12968
rect 14734 12860 14740 12912
rect 14792 12900 14798 12912
rect 14936 12900 14964 12940
rect 15013 12937 15025 12940
rect 15059 12937 15071 12971
rect 15013 12931 15071 12937
rect 17144 12940 17448 12968
rect 17144 12900 17172 12940
rect 14792 12872 14964 12900
rect 15028 12872 17172 12900
rect 14792 12860 14798 12872
rect 12894 12792 12900 12844
rect 12952 12832 12958 12844
rect 15028 12832 15056 12872
rect 12952 12804 15056 12832
rect 12952 12792 12958 12804
rect 15194 12792 15200 12844
rect 15252 12792 15258 12844
rect 16114 12792 16120 12844
rect 16172 12792 16178 12844
rect 16393 12835 16451 12841
rect 16393 12801 16405 12835
rect 16439 12832 16451 12835
rect 16439 12804 16988 12832
rect 16439 12801 16451 12804
rect 16393 12795 16451 12801
rect 13464 12736 13952 12764
rect 13464 12708 13492 12736
rect 13173 12699 13231 12705
rect 13173 12696 13185 12699
rect 12268 12668 13185 12696
rect 13173 12665 13185 12668
rect 13219 12665 13231 12699
rect 13173 12659 13231 12665
rect 13446 12656 13452 12708
rect 13504 12656 13510 12708
rect 13722 12705 13728 12708
rect 13709 12699 13728 12705
rect 13709 12665 13721 12699
rect 13709 12659 13728 12665
rect 13722 12656 13728 12659
rect 13780 12656 13786 12708
rect 13924 12705 13952 12736
rect 14366 12724 14372 12776
rect 14424 12764 14430 12776
rect 14737 12767 14795 12773
rect 14737 12764 14749 12767
rect 14424 12736 14749 12764
rect 14424 12724 14430 12736
rect 14737 12733 14749 12736
rect 14783 12733 14795 12767
rect 14737 12727 14795 12733
rect 15010 12724 15016 12776
rect 15068 12724 15074 12776
rect 15105 12767 15163 12773
rect 15105 12733 15117 12767
rect 15151 12764 15163 12767
rect 15212 12764 15240 12792
rect 15151 12736 15240 12764
rect 15151 12733 15163 12736
rect 15105 12727 15163 12733
rect 15286 12724 15292 12776
rect 15344 12724 15350 12776
rect 16025 12767 16083 12773
rect 16025 12733 16037 12767
rect 16071 12733 16083 12767
rect 16025 12727 16083 12733
rect 13909 12699 13967 12705
rect 13909 12665 13921 12699
rect 13955 12665 13967 12699
rect 13909 12659 13967 12665
rect 13998 12656 14004 12708
rect 14056 12656 14062 12708
rect 14826 12656 14832 12708
rect 14884 12696 14890 12708
rect 16040 12696 16068 12727
rect 16298 12724 16304 12776
rect 16356 12764 16362 12776
rect 16960 12773 16988 12804
rect 16761 12767 16819 12773
rect 16761 12764 16773 12767
rect 16356 12736 16773 12764
rect 16356 12724 16362 12736
rect 16761 12733 16773 12736
rect 16807 12733 16819 12767
rect 16761 12727 16819 12733
rect 16945 12767 17003 12773
rect 16945 12733 16957 12767
rect 16991 12733 17003 12767
rect 16945 12727 17003 12733
rect 14884 12668 16068 12696
rect 16776 12696 16804 12727
rect 17034 12724 17040 12776
rect 17092 12724 17098 12776
rect 17144 12773 17172 12872
rect 17313 12903 17371 12909
rect 17313 12869 17325 12903
rect 17359 12869 17371 12903
rect 17420 12900 17448 12940
rect 17678 12928 17684 12980
rect 17736 12968 17742 12980
rect 17865 12971 17923 12977
rect 17865 12968 17877 12971
rect 17736 12940 17877 12968
rect 17736 12928 17742 12940
rect 17865 12937 17877 12940
rect 17911 12937 17923 12971
rect 17865 12931 17923 12937
rect 17586 12900 17592 12912
rect 17420 12872 17592 12900
rect 17313 12863 17371 12869
rect 17218 12792 17224 12844
rect 17276 12792 17282 12844
rect 17328 12832 17356 12863
rect 17586 12860 17592 12872
rect 17644 12900 17650 12912
rect 19978 12900 19984 12912
rect 17644 12872 19984 12900
rect 17644 12860 17650 12872
rect 19978 12860 19984 12872
rect 20036 12860 20042 12912
rect 17328 12804 17632 12832
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12733 17187 12767
rect 17236 12764 17264 12792
rect 17604 12773 17632 12804
rect 17405 12767 17463 12773
rect 17405 12764 17417 12767
rect 17236 12736 17417 12764
rect 17129 12727 17187 12733
rect 17405 12733 17417 12736
rect 17451 12733 17463 12767
rect 17405 12727 17463 12733
rect 17589 12767 17647 12773
rect 17589 12733 17601 12767
rect 17635 12733 17647 12767
rect 17589 12727 17647 12733
rect 17773 12767 17831 12773
rect 17773 12733 17785 12767
rect 17819 12764 17831 12767
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 17819 12736 18061 12764
rect 17819 12733 17831 12736
rect 17773 12727 17831 12733
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 18049 12727 18107 12733
rect 19702 12696 19708 12708
rect 16776 12668 19708 12696
rect 14884 12656 14890 12668
rect 10226 12628 10232 12640
rect 8956 12600 10232 12628
rect 10226 12588 10232 12600
rect 10284 12588 10290 12640
rect 10594 12588 10600 12640
rect 10652 12588 10658 12640
rect 10778 12637 10784 12640
rect 10765 12631 10784 12637
rect 10765 12597 10777 12631
rect 10765 12591 10784 12597
rect 10778 12588 10784 12591
rect 10836 12588 10842 12640
rect 12802 12588 12808 12640
rect 12860 12588 12866 12640
rect 12973 12631 13031 12637
rect 12973 12597 12985 12631
rect 13019 12628 13031 12631
rect 13078 12628 13084 12640
rect 13019 12600 13084 12628
rect 13019 12597 13031 12600
rect 12973 12591 13031 12597
rect 13078 12588 13084 12600
rect 13136 12588 13142 12640
rect 13538 12588 13544 12640
rect 13596 12588 13602 12640
rect 14016 12628 14044 12656
rect 15102 12628 15108 12640
rect 14016 12600 15108 12628
rect 15102 12588 15108 12600
rect 15160 12588 15166 12640
rect 15194 12588 15200 12640
rect 15252 12588 15258 12640
rect 16040 12628 16068 12668
rect 19702 12656 19708 12668
rect 19760 12696 19766 12708
rect 20622 12696 20628 12708
rect 19760 12668 20628 12696
rect 19760 12656 19766 12668
rect 20622 12656 20628 12668
rect 20680 12656 20686 12708
rect 16758 12628 16764 12640
rect 16040 12600 16764 12628
rect 16758 12588 16764 12600
rect 16816 12588 16822 12640
rect 17218 12588 17224 12640
rect 17276 12628 17282 12640
rect 20346 12628 20352 12640
rect 17276 12600 20352 12628
rect 17276 12588 17282 12600
rect 20346 12588 20352 12600
rect 20404 12588 20410 12640
rect 552 12538 28587 12560
rect 552 12486 7366 12538
rect 7418 12486 7430 12538
rect 7482 12486 7494 12538
rect 7546 12486 7558 12538
rect 7610 12486 7622 12538
rect 7674 12486 14335 12538
rect 14387 12486 14399 12538
rect 14451 12486 14463 12538
rect 14515 12486 14527 12538
rect 14579 12486 14591 12538
rect 14643 12486 21304 12538
rect 21356 12486 21368 12538
rect 21420 12486 21432 12538
rect 21484 12486 21496 12538
rect 21548 12486 21560 12538
rect 21612 12486 28273 12538
rect 28325 12486 28337 12538
rect 28389 12486 28401 12538
rect 28453 12486 28465 12538
rect 28517 12486 28529 12538
rect 28581 12486 28587 12538
rect 552 12464 28587 12486
rect 4614 12384 4620 12436
rect 4672 12424 4678 12436
rect 4709 12427 4767 12433
rect 4709 12424 4721 12427
rect 4672 12396 4721 12424
rect 4672 12384 4678 12396
rect 4709 12393 4721 12396
rect 4755 12393 4767 12427
rect 9217 12427 9275 12433
rect 4709 12387 4767 12393
rect 5644 12396 6408 12424
rect 4338 12316 4344 12368
rect 4396 12316 4402 12368
rect 4724 12356 4752 12387
rect 4724 12328 5488 12356
rect 4356 12288 4384 12316
rect 5460 12300 5488 12328
rect 5644 12307 5672 12396
rect 5629 12301 5687 12307
rect 4801 12291 4859 12297
rect 4801 12288 4813 12291
rect 4356 12260 4813 12288
rect 4801 12257 4813 12260
rect 4847 12257 4859 12291
rect 4801 12251 4859 12257
rect 5442 12248 5448 12300
rect 5500 12248 5506 12300
rect 5629 12267 5641 12301
rect 5675 12267 5687 12301
rect 5629 12261 5687 12267
rect 5718 12248 5724 12300
rect 5776 12286 5782 12300
rect 6089 12291 6147 12297
rect 6089 12288 6101 12291
rect 5828 12286 6101 12288
rect 5776 12260 6101 12286
rect 5776 12258 5856 12260
rect 5776 12248 5782 12258
rect 6089 12257 6101 12260
rect 6135 12257 6147 12291
rect 6089 12251 6147 12257
rect 6178 12248 6184 12300
rect 6236 12248 6242 12300
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12257 6331 12291
rect 6273 12251 6331 12257
rect 5537 12155 5595 12161
rect 5537 12121 5549 12155
rect 5583 12152 5595 12155
rect 6288 12152 6316 12251
rect 5583 12124 6316 12152
rect 6380 12152 6408 12396
rect 6472 12396 9168 12424
rect 6472 12297 6500 12396
rect 7098 12356 7104 12368
rect 6840 12328 7104 12356
rect 6840 12297 6868 12328
rect 7098 12316 7104 12328
rect 7156 12356 7162 12368
rect 7156 12328 7604 12356
rect 7156 12316 7162 12328
rect 7576 12297 7604 12328
rect 7650 12316 7656 12368
rect 7708 12316 7714 12368
rect 8662 12356 8668 12368
rect 7760 12328 8668 12356
rect 6457 12291 6515 12297
rect 6457 12257 6469 12291
rect 6503 12257 6515 12291
rect 6457 12251 6515 12257
rect 6641 12291 6699 12297
rect 6641 12257 6653 12291
rect 6687 12257 6699 12291
rect 6641 12251 6699 12257
rect 6825 12291 6883 12297
rect 6825 12257 6837 12291
rect 6871 12257 6883 12291
rect 6825 12251 6883 12257
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12257 7343 12291
rect 7285 12251 7343 12257
rect 7561 12291 7619 12297
rect 7561 12257 7573 12291
rect 7607 12257 7619 12291
rect 7561 12251 7619 12257
rect 6656 12220 6684 12251
rect 6917 12223 6975 12229
rect 6917 12220 6929 12223
rect 6656 12192 6929 12220
rect 6917 12189 6929 12192
rect 6963 12220 6975 12223
rect 6963 12192 7144 12220
rect 6963 12189 6975 12192
rect 6917 12183 6975 12189
rect 7116 12152 7144 12192
rect 7190 12180 7196 12232
rect 7248 12180 7254 12232
rect 7300 12220 7328 12251
rect 7760 12220 7788 12328
rect 8662 12316 8668 12328
rect 8720 12316 8726 12368
rect 9140 12356 9168 12396
rect 9217 12393 9229 12427
rect 9263 12424 9275 12427
rect 9766 12424 9772 12436
rect 9263 12396 9772 12424
rect 9263 12393 9275 12396
rect 9217 12387 9275 12393
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 11348 12396 11928 12424
rect 11348 12356 11376 12396
rect 11900 12356 11928 12396
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 12158 12424 12164 12436
rect 12032 12396 12164 12424
rect 12032 12384 12038 12396
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 13078 12384 13084 12436
rect 13136 12424 13142 12436
rect 19153 12427 19211 12433
rect 13136 12396 16160 12424
rect 13136 12384 13142 12396
rect 16132 12368 16160 12396
rect 19153 12393 19165 12427
rect 19199 12424 19211 12427
rect 19199 12396 19840 12424
rect 19199 12393 19211 12396
rect 19153 12387 19211 12393
rect 13354 12356 13360 12368
rect 9140 12328 11376 12356
rect 11440 12328 11744 12356
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12257 7895 12291
rect 7837 12251 7895 12257
rect 8757 12291 8815 12297
rect 8757 12257 8769 12291
rect 8803 12288 8815 12291
rect 10502 12288 10508 12300
rect 8803 12260 10508 12288
rect 8803 12257 8815 12260
rect 8757 12251 8815 12257
rect 7300 12192 7788 12220
rect 7650 12152 7656 12164
rect 6380 12124 7052 12152
rect 7116 12124 7656 12152
rect 5583 12121 5595 12124
rect 5537 12115 5595 12121
rect 5810 12044 5816 12096
rect 5868 12044 5874 12096
rect 6822 12044 6828 12096
rect 6880 12044 6886 12096
rect 7024 12084 7052 12124
rect 7650 12112 7656 12124
rect 7708 12112 7714 12164
rect 7852 12152 7880 12251
rect 10502 12248 10508 12260
rect 10560 12248 10566 12300
rect 11440 12297 11468 12328
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12257 11483 12291
rect 11425 12251 11483 12257
rect 11609 12291 11667 12297
rect 11609 12257 11621 12291
rect 11655 12257 11667 12291
rect 11609 12251 11667 12257
rect 9858 12152 9864 12164
rect 7852 12124 9864 12152
rect 7852 12084 7880 12124
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 11624 12152 11652 12251
rect 11716 12220 11744 12328
rect 11900 12328 13360 12356
rect 11900 12288 11928 12328
rect 13354 12316 13360 12328
rect 13412 12316 13418 12368
rect 16114 12316 16120 12368
rect 16172 12316 16178 12368
rect 19812 12365 19840 12396
rect 19337 12359 19395 12365
rect 19337 12356 19349 12359
rect 18800 12328 19349 12356
rect 12069 12291 12127 12297
rect 12069 12288 12081 12291
rect 11900 12260 12081 12288
rect 12069 12257 12081 12260
rect 12115 12257 12127 12291
rect 12069 12251 12127 12257
rect 12345 12291 12403 12297
rect 12345 12257 12357 12291
rect 12391 12288 12403 12291
rect 12802 12288 12808 12300
rect 12391 12260 12808 12288
rect 12391 12257 12403 12260
rect 12345 12251 12403 12257
rect 12802 12248 12808 12260
rect 12860 12248 12866 12300
rect 18598 12248 18604 12300
rect 18656 12288 18662 12300
rect 18800 12297 18828 12328
rect 19337 12325 19349 12328
rect 19383 12325 19395 12359
rect 19337 12319 19395 12325
rect 19797 12359 19855 12365
rect 19797 12325 19809 12359
rect 19843 12325 19855 12359
rect 19797 12319 19855 12325
rect 18785 12291 18843 12297
rect 18785 12288 18797 12291
rect 18656 12260 18797 12288
rect 18656 12248 18662 12260
rect 18785 12257 18797 12260
rect 18831 12257 18843 12291
rect 18785 12251 18843 12257
rect 19150 12248 19156 12300
rect 19208 12248 19214 12300
rect 19242 12248 19248 12300
rect 19300 12248 19306 12300
rect 19613 12291 19671 12297
rect 19613 12257 19625 12291
rect 19659 12288 19671 12291
rect 19702 12288 19708 12300
rect 19659 12260 19708 12288
rect 19659 12257 19671 12260
rect 19613 12251 19671 12257
rect 19702 12248 19708 12260
rect 19760 12248 19766 12300
rect 19889 12291 19947 12297
rect 19889 12257 19901 12291
rect 19935 12257 19947 12291
rect 19889 12251 19947 12257
rect 11882 12220 11888 12232
rect 11716 12192 11888 12220
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 12253 12223 12311 12229
rect 12253 12189 12265 12223
rect 12299 12220 12311 12223
rect 13538 12220 13544 12232
rect 12299 12192 13544 12220
rect 12299 12189 12311 12192
rect 12253 12183 12311 12189
rect 13538 12180 13544 12192
rect 13596 12180 13602 12232
rect 18877 12223 18935 12229
rect 18877 12189 18889 12223
rect 18923 12189 18935 12223
rect 19168 12220 19196 12248
rect 19904 12220 19932 12251
rect 19978 12248 19984 12300
rect 20036 12248 20042 12300
rect 20346 12248 20352 12300
rect 20404 12248 20410 12300
rect 20441 12291 20499 12297
rect 20441 12257 20453 12291
rect 20487 12257 20499 12291
rect 20441 12251 20499 12257
rect 20625 12291 20683 12297
rect 20625 12257 20637 12291
rect 20671 12288 20683 12291
rect 20717 12291 20775 12297
rect 20717 12288 20729 12291
rect 20671 12260 20729 12288
rect 20671 12257 20683 12260
rect 20625 12251 20683 12257
rect 20717 12257 20729 12260
rect 20763 12257 20775 12291
rect 20717 12251 20775 12257
rect 20456 12220 20484 12251
rect 19168 12192 19932 12220
rect 20180 12192 20484 12220
rect 18877 12183 18935 12189
rect 13078 12152 13084 12164
rect 11624 12124 13084 12152
rect 13078 12112 13084 12124
rect 13136 12112 13142 12164
rect 13262 12112 13268 12164
rect 13320 12152 13326 12164
rect 18892 12152 18920 12183
rect 19610 12152 19616 12164
rect 13320 12124 16436 12152
rect 18892 12124 19616 12152
rect 13320 12112 13326 12124
rect 16408 12096 16436 12124
rect 19610 12112 19616 12124
rect 19668 12112 19674 12164
rect 20180 12161 20208 12192
rect 20165 12155 20223 12161
rect 20165 12121 20177 12155
rect 20211 12121 20223 12155
rect 20165 12115 20223 12121
rect 7024 12056 7880 12084
rect 8018 12044 8024 12096
rect 8076 12044 8082 12096
rect 8938 12044 8944 12096
rect 8996 12044 9002 12096
rect 9582 12044 9588 12096
rect 9640 12084 9646 12096
rect 11514 12084 11520 12096
rect 9640 12056 11520 12084
rect 9640 12044 9646 12056
rect 11514 12044 11520 12056
rect 11572 12044 11578 12096
rect 11885 12087 11943 12093
rect 11885 12053 11897 12087
rect 11931 12084 11943 12087
rect 12158 12084 12164 12096
rect 11931 12056 12164 12084
rect 11931 12053 11943 12056
rect 11885 12047 11943 12053
rect 12158 12044 12164 12056
rect 12216 12044 12222 12096
rect 13722 12044 13728 12096
rect 13780 12084 13786 12096
rect 14918 12084 14924 12096
rect 13780 12056 14924 12084
rect 13780 12044 13786 12056
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 16390 12044 16396 12096
rect 16448 12044 16454 12096
rect 20898 12044 20904 12096
rect 20956 12044 20962 12096
rect 552 11994 28428 12016
rect 552 11942 3882 11994
rect 3934 11942 3946 11994
rect 3998 11942 4010 11994
rect 4062 11942 4074 11994
rect 4126 11942 4138 11994
rect 4190 11942 10851 11994
rect 10903 11942 10915 11994
rect 10967 11942 10979 11994
rect 11031 11942 11043 11994
rect 11095 11942 11107 11994
rect 11159 11942 17820 11994
rect 17872 11942 17884 11994
rect 17936 11942 17948 11994
rect 18000 11942 18012 11994
rect 18064 11942 18076 11994
rect 18128 11942 24789 11994
rect 24841 11942 24853 11994
rect 24905 11942 24917 11994
rect 24969 11942 24981 11994
rect 25033 11942 25045 11994
rect 25097 11942 28428 11994
rect 552 11920 28428 11942
rect 3786 11840 3792 11892
rect 3844 11840 3850 11892
rect 5810 11840 5816 11892
rect 5868 11840 5874 11892
rect 6822 11840 6828 11892
rect 6880 11840 6886 11892
rect 8018 11880 8024 11892
rect 7024 11852 8024 11880
rect 5828 11744 5856 11840
rect 5092 11716 5856 11744
rect 4913 11679 4971 11685
rect 4913 11645 4925 11679
rect 4959 11676 4971 11679
rect 5092 11676 5120 11716
rect 4959 11648 5120 11676
rect 5169 11679 5227 11685
rect 4959 11645 4971 11648
rect 4913 11639 4971 11645
rect 5169 11645 5181 11679
rect 5215 11676 5227 11679
rect 5902 11676 5908 11688
rect 5215 11648 5908 11676
rect 5215 11645 5227 11648
rect 5169 11639 5227 11645
rect 5902 11636 5908 11648
rect 5960 11676 5966 11688
rect 6638 11676 6644 11688
rect 5960 11648 6644 11676
rect 5960 11636 5966 11648
rect 6638 11636 6644 11648
rect 6696 11636 6702 11688
rect 6840 11676 6868 11840
rect 7024 11685 7052 11852
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 8849 11883 8907 11889
rect 8849 11849 8861 11883
rect 8895 11880 8907 11883
rect 9306 11880 9312 11892
rect 8895 11852 9312 11880
rect 8895 11849 8907 11852
rect 8849 11843 8907 11849
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 9674 11840 9680 11892
rect 9732 11840 9738 11892
rect 10413 11883 10471 11889
rect 10413 11849 10425 11883
rect 10459 11880 10471 11883
rect 10594 11880 10600 11892
rect 10459 11852 10600 11880
rect 10459 11849 10471 11852
rect 10413 11843 10471 11849
rect 10594 11840 10600 11852
rect 10652 11840 10658 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11572 11852 13952 11880
rect 11572 11840 11578 11852
rect 7193 11815 7251 11821
rect 7193 11781 7205 11815
rect 7239 11812 7251 11815
rect 9582 11812 9588 11824
rect 7239 11784 9588 11812
rect 7239 11781 7251 11784
rect 7193 11775 7251 11781
rect 9582 11772 9588 11784
rect 9640 11772 9646 11824
rect 9398 11744 9404 11756
rect 8864 11716 9404 11744
rect 6917 11679 6975 11685
rect 6917 11676 6929 11679
rect 6840 11648 6929 11676
rect 6917 11645 6929 11648
rect 6963 11645 6975 11679
rect 6917 11639 6975 11645
rect 7009 11679 7067 11685
rect 7009 11645 7021 11679
rect 7055 11645 7067 11679
rect 7009 11639 7067 11645
rect 7285 11679 7343 11685
rect 7285 11645 7297 11679
rect 7331 11676 7343 11679
rect 8110 11676 8116 11688
rect 7331 11648 8116 11676
rect 7331 11645 7343 11648
rect 7285 11639 7343 11645
rect 7190 11608 7196 11620
rect 7024 11580 7196 11608
rect 7024 11552 7052 11580
rect 7190 11568 7196 11580
rect 7248 11608 7254 11620
rect 7300 11608 7328 11639
rect 8110 11636 8116 11648
rect 8168 11636 8174 11688
rect 8864 11685 8892 11716
rect 9398 11704 9404 11716
rect 9456 11704 9462 11756
rect 9493 11747 9551 11753
rect 9493 11713 9505 11747
rect 9539 11744 9551 11747
rect 9692 11744 9720 11840
rect 9858 11772 9864 11824
rect 9916 11812 9922 11824
rect 13081 11815 13139 11821
rect 9916 11784 10364 11812
rect 9916 11772 9922 11784
rect 10336 11753 10364 11784
rect 13081 11781 13093 11815
rect 13127 11812 13139 11815
rect 13127 11784 13709 11812
rect 13127 11781 13139 11784
rect 13081 11775 13139 11781
rect 10321 11747 10379 11753
rect 9539 11716 10088 11744
rect 9539 11713 9551 11716
rect 9493 11707 9551 11713
rect 8849 11679 8907 11685
rect 8849 11645 8861 11679
rect 8895 11645 8907 11679
rect 8849 11639 8907 11645
rect 9125 11679 9183 11685
rect 9125 11645 9137 11679
rect 9171 11676 9183 11679
rect 9508 11676 9536 11707
rect 9171 11648 9536 11676
rect 9585 11679 9643 11685
rect 9171 11645 9183 11648
rect 9125 11639 9183 11645
rect 9585 11645 9597 11679
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 9858 11676 9864 11688
rect 9723 11648 9864 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 7248 11580 7328 11608
rect 9033 11611 9091 11617
rect 7248 11568 7254 11580
rect 9033 11577 9045 11611
rect 9079 11608 9091 11611
rect 9600 11608 9628 11639
rect 9858 11636 9864 11648
rect 9916 11636 9922 11688
rect 10060 11685 10088 11716
rect 10321 11713 10333 11747
rect 10367 11744 10379 11747
rect 13446 11744 13452 11756
rect 10367 11716 12112 11744
rect 10367 11713 10379 11716
rect 10321 11707 10379 11713
rect 10045 11679 10103 11685
rect 10045 11645 10057 11679
rect 10091 11645 10103 11679
rect 10045 11639 10103 11645
rect 9766 11608 9772 11620
rect 9079 11580 9772 11608
rect 9079 11577 9091 11580
rect 9033 11571 9091 11577
rect 9766 11568 9772 11580
rect 9824 11568 9830 11620
rect 11977 11611 12035 11617
rect 11977 11608 11989 11611
rect 10152 11580 11989 11608
rect 10152 11552 10180 11580
rect 11977 11577 11989 11580
rect 12023 11577 12035 11611
rect 12084 11608 12112 11716
rect 12406 11716 13452 11744
rect 12161 11679 12219 11685
rect 12161 11645 12173 11679
rect 12207 11676 12219 11679
rect 12406 11676 12434 11716
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 12207 11648 12434 11676
rect 13265 11679 13323 11685
rect 12207 11645 12219 11648
rect 12161 11639 12219 11645
rect 13265 11645 13277 11679
rect 13311 11645 13323 11679
rect 13265 11639 13323 11645
rect 13078 11608 13084 11620
rect 12084 11580 13084 11608
rect 11977 11571 12035 11577
rect 6730 11500 6736 11552
rect 6788 11500 6794 11552
rect 7006 11500 7012 11552
rect 7064 11500 7070 11552
rect 9214 11500 9220 11552
rect 9272 11500 9278 11552
rect 10134 11500 10140 11552
rect 10192 11500 10198 11552
rect 10410 11500 10416 11552
rect 10468 11540 10474 11552
rect 10597 11543 10655 11549
rect 10597 11540 10609 11543
rect 10468 11512 10609 11540
rect 10468 11500 10474 11512
rect 10597 11509 10609 11512
rect 10643 11509 10655 11543
rect 10597 11503 10655 11509
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11664 11512 11805 11540
rect 11664 11500 11670 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11992 11540 12020 11571
rect 13078 11568 13084 11580
rect 13136 11568 13142 11620
rect 13280 11608 13308 11639
rect 13354 11636 13360 11688
rect 13412 11636 13418 11688
rect 13681 11685 13709 11784
rect 13924 11744 13952 11852
rect 14918 11840 14924 11892
rect 14976 11880 14982 11892
rect 14976 11852 15976 11880
rect 14976 11840 14982 11852
rect 14090 11772 14096 11824
rect 14148 11772 14154 11824
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 13924 11716 14197 11744
rect 14185 11713 14197 11716
rect 14231 11713 14243 11747
rect 14185 11707 14243 11713
rect 13666 11679 13724 11685
rect 13666 11645 13678 11679
rect 13712 11645 13724 11679
rect 14461 11679 14519 11685
rect 14461 11676 14473 11679
rect 13666 11639 13724 11645
rect 14108 11648 14473 11676
rect 14108 11608 14136 11648
rect 14461 11645 14473 11648
rect 14507 11676 14519 11679
rect 14734 11676 14740 11688
rect 14507 11648 14740 11676
rect 14507 11645 14519 11648
rect 14461 11639 14519 11645
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 14936 11676 14964 11840
rect 15013 11815 15071 11821
rect 15013 11781 15025 11815
rect 15059 11812 15071 11815
rect 15194 11812 15200 11824
rect 15059 11784 15200 11812
rect 15059 11781 15071 11784
rect 15013 11775 15071 11781
rect 15194 11772 15200 11784
rect 15252 11772 15258 11824
rect 15948 11812 15976 11852
rect 18138 11840 18144 11892
rect 18196 11880 18202 11892
rect 18196 11852 21220 11880
rect 18196 11840 18202 11852
rect 18417 11815 18475 11821
rect 15948 11784 16068 11812
rect 15212 11744 15240 11772
rect 15212 11716 15976 11744
rect 15197 11679 15255 11685
rect 15197 11676 15209 11679
rect 14936 11648 15209 11676
rect 15197 11645 15209 11648
rect 15243 11645 15255 11679
rect 15197 11639 15255 11645
rect 15378 11636 15384 11688
rect 15436 11676 15442 11688
rect 15948 11685 15976 11716
rect 16040 11685 16068 11784
rect 18417 11781 18429 11815
rect 18463 11812 18475 11815
rect 19242 11812 19248 11824
rect 18463 11784 19248 11812
rect 18463 11781 18475 11784
rect 18417 11775 18475 11781
rect 19242 11772 19248 11784
rect 19300 11772 19306 11824
rect 19797 11815 19855 11821
rect 19797 11781 19809 11815
rect 19843 11781 19855 11815
rect 19797 11775 19855 11781
rect 18141 11747 18199 11753
rect 18141 11713 18153 11747
rect 18187 11744 18199 11747
rect 19150 11744 19156 11756
rect 18187 11716 19156 11744
rect 18187 11713 18199 11716
rect 18141 11707 18199 11713
rect 19150 11704 19156 11716
rect 19208 11744 19214 11756
rect 19812 11744 19840 11775
rect 21192 11753 21220 11852
rect 22002 11840 22008 11892
rect 22060 11840 22066 11892
rect 19208 11716 19840 11744
rect 21177 11747 21235 11753
rect 19208 11704 19214 11716
rect 21177 11713 21189 11747
rect 21223 11744 21235 11747
rect 22020 11744 22048 11840
rect 21223 11716 22048 11744
rect 21223 11713 21235 11716
rect 21177 11707 21235 11713
rect 15657 11679 15715 11685
rect 15657 11676 15669 11679
rect 15436 11648 15669 11676
rect 15436 11636 15442 11648
rect 15657 11645 15669 11648
rect 15703 11645 15715 11679
rect 15657 11639 15715 11645
rect 15933 11679 15991 11685
rect 15933 11645 15945 11679
rect 15979 11645 15991 11679
rect 15933 11639 15991 11645
rect 16025 11679 16083 11685
rect 16025 11645 16037 11679
rect 16071 11645 16083 11679
rect 16025 11639 16083 11645
rect 18049 11679 18107 11685
rect 18049 11645 18061 11679
rect 18095 11676 18107 11679
rect 18782 11676 18788 11688
rect 18095 11648 18788 11676
rect 18095 11645 18107 11648
rect 18049 11639 18107 11645
rect 18782 11636 18788 11648
rect 18840 11636 18846 11688
rect 20898 11636 20904 11688
rect 20956 11685 20962 11688
rect 20956 11676 20968 11685
rect 20956 11648 21001 11676
rect 20956 11639 20968 11648
rect 20956 11636 20962 11639
rect 13280 11580 14136 11608
rect 14182 11568 14188 11620
rect 14240 11608 14246 11620
rect 14277 11611 14335 11617
rect 14277 11608 14289 11611
rect 14240 11580 14289 11608
rect 14240 11568 14246 11580
rect 14277 11577 14289 11580
rect 14323 11577 14335 11611
rect 14277 11571 14335 11577
rect 15286 11568 15292 11620
rect 15344 11608 15350 11620
rect 15841 11611 15899 11617
rect 15841 11608 15853 11611
rect 15344 11580 15853 11608
rect 15344 11568 15350 11580
rect 15841 11577 15853 11580
rect 15887 11577 15899 11611
rect 15841 11571 15899 11577
rect 13262 11540 13268 11552
rect 11992 11512 13268 11540
rect 11793 11503 11851 11509
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 13538 11500 13544 11552
rect 13596 11500 13602 11552
rect 13725 11543 13783 11549
rect 13725 11509 13737 11543
rect 13771 11540 13783 11543
rect 14645 11543 14703 11549
rect 14645 11540 14657 11543
rect 13771 11512 14657 11540
rect 13771 11509 13783 11512
rect 13725 11503 13783 11509
rect 14645 11509 14657 11512
rect 14691 11509 14703 11543
rect 14645 11503 14703 11509
rect 15378 11500 15384 11552
rect 15436 11500 15442 11552
rect 15562 11500 15568 11552
rect 15620 11500 15626 11552
rect 16206 11500 16212 11552
rect 16264 11500 16270 11552
rect 552 11450 28587 11472
rect 552 11398 7366 11450
rect 7418 11398 7430 11450
rect 7482 11398 7494 11450
rect 7546 11398 7558 11450
rect 7610 11398 7622 11450
rect 7674 11398 14335 11450
rect 14387 11398 14399 11450
rect 14451 11398 14463 11450
rect 14515 11398 14527 11450
rect 14579 11398 14591 11450
rect 14643 11398 21304 11450
rect 21356 11398 21368 11450
rect 21420 11398 21432 11450
rect 21484 11398 21496 11450
rect 21548 11398 21560 11450
rect 21612 11398 28273 11450
rect 28325 11398 28337 11450
rect 28389 11398 28401 11450
rect 28453 11398 28465 11450
rect 28517 11398 28529 11450
rect 28581 11398 28587 11450
rect 552 11376 28587 11398
rect 6178 11296 6184 11348
rect 6236 11336 6242 11348
rect 8665 11339 8723 11345
rect 8665 11336 8677 11339
rect 6236 11308 8677 11336
rect 6236 11296 6242 11308
rect 8665 11305 8677 11308
rect 8711 11336 8723 11339
rect 8938 11336 8944 11348
rect 8711 11308 8944 11336
rect 8711 11305 8723 11308
rect 8665 11299 8723 11305
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 9214 11336 9220 11348
rect 9048 11308 9220 11336
rect 9048 11268 9076 11308
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 10321 11339 10379 11345
rect 9646 11308 10272 11336
rect 8956 11240 9076 11268
rect 6730 11160 6736 11212
rect 6788 11160 6794 11212
rect 6917 11203 6975 11209
rect 6917 11169 6929 11203
rect 6963 11169 6975 11203
rect 6917 11163 6975 11169
rect 7101 11203 7159 11209
rect 7101 11169 7113 11203
rect 7147 11200 7159 11203
rect 7193 11203 7251 11209
rect 7193 11200 7205 11203
rect 7147 11172 7205 11200
rect 7147 11169 7159 11172
rect 7101 11163 7159 11169
rect 7193 11169 7205 11172
rect 7239 11169 7251 11203
rect 7193 11163 7251 11169
rect 8113 11203 8171 11209
rect 8113 11169 8125 11203
rect 8159 11169 8171 11203
rect 8113 11163 8171 11169
rect 8297 11203 8355 11209
rect 8297 11169 8309 11203
rect 8343 11200 8355 11203
rect 8662 11203 8720 11209
rect 8343 11172 8524 11200
rect 8343 11169 8355 11172
rect 8297 11163 8355 11169
rect 6932 11132 6960 11163
rect 8128 11132 8156 11163
rect 6932 11104 8156 11132
rect 7374 10956 7380 11008
rect 7432 10956 7438 11008
rect 8128 10996 8156 11104
rect 8202 11092 8208 11144
rect 8260 11092 8266 11144
rect 8496 11073 8524 11172
rect 8662 11169 8674 11203
rect 8708 11200 8720 11203
rect 8754 11200 8760 11212
rect 8708 11172 8760 11200
rect 8708 11169 8720 11172
rect 8662 11163 8720 11169
rect 8754 11160 8760 11172
rect 8812 11200 8818 11212
rect 8812 11172 8892 11200
rect 8812 11160 8818 11172
rect 8481 11067 8539 11073
rect 8481 11033 8493 11067
rect 8527 11033 8539 11067
rect 8864 11064 8892 11172
rect 8956 11132 8984 11240
rect 9122 11228 9128 11280
rect 9180 11268 9186 11280
rect 9646 11268 9674 11308
rect 9180 11240 9674 11268
rect 9180 11228 9186 11240
rect 10134 11228 10140 11280
rect 10192 11228 10198 11280
rect 10244 11268 10272 11308
rect 10321 11305 10333 11339
rect 10367 11336 10379 11339
rect 10597 11339 10655 11345
rect 10597 11336 10609 11339
rect 10367 11308 10609 11336
rect 10367 11305 10379 11308
rect 10321 11299 10379 11305
rect 10597 11305 10609 11308
rect 10643 11305 10655 11339
rect 10597 11299 10655 11305
rect 11698 11296 11704 11348
rect 11756 11296 11762 11348
rect 13081 11339 13139 11345
rect 13081 11305 13093 11339
rect 13127 11305 13139 11339
rect 13081 11299 13139 11305
rect 11716 11268 11744 11296
rect 10244 11240 11744 11268
rect 13096 11268 13124 11299
rect 13354 11296 13360 11348
rect 13412 11336 13418 11348
rect 13449 11339 13507 11345
rect 13449 11336 13461 11339
rect 13412 11308 13461 11336
rect 13412 11296 13418 11308
rect 13449 11305 13461 11308
rect 13495 11336 13507 11339
rect 14182 11336 14188 11348
rect 13495 11308 14188 11336
rect 13495 11305 13507 11308
rect 13449 11299 13507 11305
rect 14182 11296 14188 11308
rect 14240 11296 14246 11348
rect 14826 11336 14832 11348
rect 14568 11308 14832 11336
rect 14090 11268 14096 11280
rect 13096 11240 14096 11268
rect 10152 11200 10180 11228
rect 9646 11172 10180 11200
rect 9033 11135 9091 11141
rect 9033 11132 9045 11135
rect 8956 11104 9045 11132
rect 9033 11101 9045 11104
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 9306 11132 9312 11144
rect 9171 11104 9312 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 9306 11092 9312 11104
rect 9364 11092 9370 11144
rect 9214 11064 9220 11076
rect 8864 11036 9220 11064
rect 8481 11027 8539 11033
rect 9214 11024 9220 11036
rect 9272 11024 9278 11076
rect 9646 10996 9674 11172
rect 10410 11160 10416 11212
rect 10468 11160 10474 11212
rect 10520 11209 10548 11240
rect 10505 11203 10563 11209
rect 10505 11169 10517 11203
rect 10551 11169 10563 11203
rect 10505 11163 10563 11169
rect 10689 11203 10747 11209
rect 10689 11169 10701 11203
rect 10735 11200 10747 11203
rect 10965 11203 11023 11209
rect 10965 11200 10977 11203
rect 10735 11172 10977 11200
rect 10735 11169 10747 11172
rect 10689 11163 10747 11169
rect 10965 11169 10977 11172
rect 11011 11169 11023 11203
rect 11701 11203 11759 11209
rect 11701 11200 11713 11203
rect 10965 11163 11023 11169
rect 11256 11172 11713 11200
rect 11256 11144 11284 11172
rect 11701 11169 11713 11172
rect 11747 11169 11759 11203
rect 11701 11163 11759 11169
rect 11790 11160 11796 11212
rect 11848 11200 11854 11212
rect 11957 11203 12015 11209
rect 11957 11200 11969 11203
rect 11848 11172 11969 11200
rect 11848 11160 11854 11172
rect 11957 11169 11969 11172
rect 12003 11169 12015 11203
rect 11957 11163 12015 11169
rect 11238 11092 11244 11144
rect 11296 11092 11302 11144
rect 13740 11141 13768 11240
rect 14090 11228 14096 11240
rect 14148 11228 14154 11280
rect 14568 11209 14596 11308
rect 14826 11296 14832 11308
rect 14884 11296 14890 11348
rect 15197 11339 15255 11345
rect 15197 11305 15209 11339
rect 15243 11336 15255 11339
rect 15286 11336 15292 11348
rect 15243 11308 15292 11336
rect 15243 11305 15255 11308
rect 15197 11299 15255 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 15562 11296 15568 11348
rect 15620 11296 15626 11348
rect 16206 11296 16212 11348
rect 16264 11296 16270 11348
rect 14645 11271 14703 11277
rect 14645 11237 14657 11271
rect 14691 11268 14703 11271
rect 15378 11268 15384 11280
rect 14691 11240 15384 11268
rect 14691 11237 14703 11240
rect 14645 11231 14703 11237
rect 15378 11228 15384 11240
rect 15436 11228 15442 11280
rect 13817 11203 13875 11209
rect 13817 11169 13829 11203
rect 13863 11169 13875 11203
rect 13817 11163 13875 11169
rect 14553 11203 14611 11209
rect 14553 11169 14565 11203
rect 14599 11169 14611 11203
rect 14553 11163 14611 11169
rect 14737 11203 14795 11209
rect 14737 11169 14749 11203
rect 14783 11169 14795 11203
rect 14737 11163 14795 11169
rect 11517 11135 11575 11141
rect 11517 11101 11529 11135
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11101 13783 11135
rect 13832 11132 13860 11163
rect 14752 11132 14780 11163
rect 14826 11160 14832 11212
rect 14884 11160 14890 11212
rect 15010 11160 15016 11212
rect 15068 11160 15074 11212
rect 15580 11209 15608 11296
rect 16224 11268 16252 11296
rect 15948 11240 16252 11268
rect 15948 11209 15976 11240
rect 16390 11228 16396 11280
rect 16448 11228 16454 11280
rect 15565 11203 15623 11209
rect 15565 11169 15577 11203
rect 15611 11169 15623 11203
rect 15565 11163 15623 11169
rect 15933 11203 15991 11209
rect 15933 11169 15945 11203
rect 15979 11169 15991 11203
rect 15933 11163 15991 11169
rect 16117 11203 16175 11209
rect 16117 11169 16129 11203
rect 16163 11169 16175 11203
rect 16117 11163 16175 11169
rect 16209 11203 16267 11209
rect 16209 11169 16221 11203
rect 16255 11169 16267 11203
rect 17690 11203 17748 11209
rect 17690 11200 17702 11203
rect 16209 11163 16267 11169
rect 16960 11172 17702 11200
rect 15028 11132 15056 11160
rect 16132 11132 16160 11163
rect 13832 11104 15056 11132
rect 15396 11104 16160 11132
rect 16224 11132 16252 11163
rect 16850 11132 16856 11144
rect 16224 11104 16856 11132
rect 13725 11095 13783 11101
rect 10502 11024 10508 11076
rect 10560 11064 10566 11076
rect 11330 11064 11336 11076
rect 10560 11036 11336 11064
rect 10560 11024 10566 11036
rect 11330 11024 11336 11036
rect 11388 11064 11394 11076
rect 11532 11064 11560 11095
rect 11388 11036 11560 11064
rect 11388 11024 11394 11036
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 15396 11073 15424 11104
rect 16850 11092 16856 11104
rect 16908 11092 16914 11144
rect 15381 11067 15439 11073
rect 14884 11036 15332 11064
rect 14884 11024 14890 11036
rect 8128 10968 9674 10996
rect 10134 10956 10140 11008
rect 10192 10956 10198 11008
rect 15304 10996 15332 11036
rect 15381 11033 15393 11067
rect 15427 11033 15439 11067
rect 16393 11067 16451 11073
rect 15381 11027 15439 11033
rect 15488 11036 16344 11064
rect 15488 10996 15516 11036
rect 15304 10968 15516 10996
rect 15841 10999 15899 11005
rect 15841 10965 15853 10999
rect 15887 10996 15899 10999
rect 16114 10996 16120 11008
rect 15887 10968 16120 10996
rect 15887 10965 15899 10968
rect 15841 10959 15899 10965
rect 16114 10956 16120 10968
rect 16172 10956 16178 11008
rect 16316 10996 16344 11036
rect 16393 11033 16405 11067
rect 16439 11064 16451 11067
rect 16960 11064 16988 11172
rect 17690 11169 17702 11172
rect 17736 11169 17748 11203
rect 17690 11163 17748 11169
rect 17957 11203 18015 11209
rect 17957 11169 17969 11203
rect 18003 11200 18015 11203
rect 18138 11200 18144 11212
rect 18003 11172 18144 11200
rect 18003 11169 18015 11172
rect 17957 11163 18015 11169
rect 18138 11160 18144 11172
rect 18196 11160 18202 11212
rect 16439 11036 16988 11064
rect 16439 11033 16451 11036
rect 16393 11027 16451 11033
rect 16574 10996 16580 11008
rect 16316 10968 16580 10996
rect 16574 10956 16580 10968
rect 16632 10956 16638 11008
rect 552 10906 28428 10928
rect 552 10854 3882 10906
rect 3934 10854 3946 10906
rect 3998 10854 4010 10906
rect 4062 10854 4074 10906
rect 4126 10854 4138 10906
rect 4190 10854 10851 10906
rect 10903 10854 10915 10906
rect 10967 10854 10979 10906
rect 11031 10854 11043 10906
rect 11095 10854 11107 10906
rect 11159 10854 17820 10906
rect 17872 10854 17884 10906
rect 17936 10854 17948 10906
rect 18000 10854 18012 10906
rect 18064 10854 18076 10906
rect 18128 10854 24789 10906
rect 24841 10854 24853 10906
rect 24905 10854 24917 10906
rect 24969 10854 24981 10906
rect 25033 10854 25045 10906
rect 25097 10854 28428 10906
rect 552 10832 28428 10854
rect 6273 10795 6331 10801
rect 6273 10761 6285 10795
rect 6319 10792 6331 10795
rect 7006 10792 7012 10804
rect 6319 10764 7012 10792
rect 6319 10761 6331 10764
rect 6273 10755 6331 10761
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 11241 10795 11299 10801
rect 11241 10761 11253 10795
rect 11287 10792 11299 10795
rect 11330 10792 11336 10804
rect 11287 10764 11336 10792
rect 11287 10761 11299 10764
rect 11241 10755 11299 10761
rect 11330 10752 11336 10764
rect 11388 10752 11394 10804
rect 11609 10795 11667 10801
rect 11609 10761 11621 10795
rect 11655 10792 11667 10795
rect 11790 10792 11796 10804
rect 11655 10764 11796 10792
rect 11655 10761 11667 10764
rect 11609 10755 11667 10761
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 16850 10752 16856 10804
rect 16908 10792 16914 10804
rect 17497 10795 17555 10801
rect 17497 10792 17509 10795
rect 16908 10764 17509 10792
rect 16908 10752 16914 10764
rect 17497 10761 17509 10764
rect 17543 10761 17555 10795
rect 17497 10755 17555 10761
rect 11606 10616 11612 10668
rect 11664 10616 11670 10668
rect 16574 10616 16580 10668
rect 16632 10656 16638 10668
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 16632 10628 16681 10656
rect 16632 10616 16638 10628
rect 16669 10625 16681 10628
rect 16715 10625 16727 10659
rect 16669 10619 16727 10625
rect 6638 10548 6644 10600
rect 6696 10588 6702 10600
rect 7653 10591 7711 10597
rect 7653 10588 7665 10591
rect 6696 10560 7665 10588
rect 6696 10548 6702 10560
rect 7653 10557 7665 10560
rect 7699 10588 7711 10591
rect 9861 10591 9919 10597
rect 7699 10560 7880 10588
rect 7699 10557 7711 10560
rect 7653 10551 7711 10557
rect 7374 10480 7380 10532
rect 7432 10529 7438 10532
rect 7432 10520 7444 10529
rect 7432 10492 7477 10520
rect 7432 10483 7444 10492
rect 7432 10480 7438 10483
rect 7852 10464 7880 10560
rect 9861 10557 9873 10591
rect 9907 10588 9919 10591
rect 11238 10588 11244 10600
rect 9907 10560 11244 10588
rect 9907 10557 9919 10560
rect 9861 10551 9919 10557
rect 11238 10548 11244 10560
rect 11296 10548 11302 10600
rect 11425 10591 11483 10597
rect 11425 10557 11437 10591
rect 11471 10588 11483 10591
rect 11624 10588 11652 10616
rect 11471 10560 11652 10588
rect 17313 10591 17371 10597
rect 11471 10557 11483 10560
rect 11425 10551 11483 10557
rect 17313 10557 17325 10591
rect 17359 10588 17371 10591
rect 17405 10591 17463 10597
rect 17405 10588 17417 10591
rect 17359 10560 17417 10588
rect 17359 10557 17371 10560
rect 17313 10551 17371 10557
rect 17405 10557 17417 10560
rect 17451 10557 17463 10591
rect 17405 10551 17463 10557
rect 17586 10548 17592 10600
rect 17644 10548 17650 10600
rect 10134 10529 10140 10532
rect 10128 10520 10140 10529
rect 10095 10492 10140 10520
rect 10128 10483 10140 10492
rect 10134 10480 10140 10483
rect 10192 10480 10198 10532
rect 7834 10412 7840 10464
rect 7892 10412 7898 10464
rect 552 10362 28587 10384
rect 552 10310 7366 10362
rect 7418 10310 7430 10362
rect 7482 10310 7494 10362
rect 7546 10310 7558 10362
rect 7610 10310 7622 10362
rect 7674 10310 14335 10362
rect 14387 10310 14399 10362
rect 14451 10310 14463 10362
rect 14515 10310 14527 10362
rect 14579 10310 14591 10362
rect 14643 10310 21304 10362
rect 21356 10310 21368 10362
rect 21420 10310 21432 10362
rect 21484 10310 21496 10362
rect 21548 10310 21560 10362
rect 21612 10310 28273 10362
rect 28325 10310 28337 10362
rect 28389 10310 28401 10362
rect 28453 10310 28465 10362
rect 28517 10310 28529 10362
rect 28581 10310 28587 10362
rect 552 10288 28587 10310
rect 9214 10208 9220 10260
rect 9272 10208 9278 10260
rect 8104 10183 8162 10189
rect 8104 10149 8116 10183
rect 8150 10180 8162 10183
rect 8202 10180 8208 10192
rect 8150 10152 8208 10180
rect 8150 10149 8162 10152
rect 8104 10143 8162 10149
rect 8202 10140 8208 10152
rect 8260 10140 8266 10192
rect 7834 10072 7840 10124
rect 7892 10072 7898 10124
rect 552 9818 28428 9840
rect 552 9766 3882 9818
rect 3934 9766 3946 9818
rect 3998 9766 4010 9818
rect 4062 9766 4074 9818
rect 4126 9766 4138 9818
rect 4190 9766 10851 9818
rect 10903 9766 10915 9818
rect 10967 9766 10979 9818
rect 11031 9766 11043 9818
rect 11095 9766 11107 9818
rect 11159 9766 17820 9818
rect 17872 9766 17884 9818
rect 17936 9766 17948 9818
rect 18000 9766 18012 9818
rect 18064 9766 18076 9818
rect 18128 9766 24789 9818
rect 24841 9766 24853 9818
rect 24905 9766 24917 9818
rect 24969 9766 24981 9818
rect 25033 9766 25045 9818
rect 25097 9766 28428 9818
rect 552 9744 28428 9766
rect 552 9274 28587 9296
rect 552 9222 7366 9274
rect 7418 9222 7430 9274
rect 7482 9222 7494 9274
rect 7546 9222 7558 9274
rect 7610 9222 7622 9274
rect 7674 9222 14335 9274
rect 14387 9222 14399 9274
rect 14451 9222 14463 9274
rect 14515 9222 14527 9274
rect 14579 9222 14591 9274
rect 14643 9222 21304 9274
rect 21356 9222 21368 9274
rect 21420 9222 21432 9274
rect 21484 9222 21496 9274
rect 21548 9222 21560 9274
rect 21612 9222 28273 9274
rect 28325 9222 28337 9274
rect 28389 9222 28401 9274
rect 28453 9222 28465 9274
rect 28517 9222 28529 9274
rect 28581 9222 28587 9274
rect 552 9200 28587 9222
rect 552 8730 28428 8752
rect 552 8678 3882 8730
rect 3934 8678 3946 8730
rect 3998 8678 4010 8730
rect 4062 8678 4074 8730
rect 4126 8678 4138 8730
rect 4190 8678 10851 8730
rect 10903 8678 10915 8730
rect 10967 8678 10979 8730
rect 11031 8678 11043 8730
rect 11095 8678 11107 8730
rect 11159 8678 17820 8730
rect 17872 8678 17884 8730
rect 17936 8678 17948 8730
rect 18000 8678 18012 8730
rect 18064 8678 18076 8730
rect 18128 8678 24789 8730
rect 24841 8678 24853 8730
rect 24905 8678 24917 8730
rect 24969 8678 24981 8730
rect 25033 8678 25045 8730
rect 25097 8678 28428 8730
rect 552 8656 28428 8678
rect 552 8186 28587 8208
rect 552 8134 7366 8186
rect 7418 8134 7430 8186
rect 7482 8134 7494 8186
rect 7546 8134 7558 8186
rect 7610 8134 7622 8186
rect 7674 8134 14335 8186
rect 14387 8134 14399 8186
rect 14451 8134 14463 8186
rect 14515 8134 14527 8186
rect 14579 8134 14591 8186
rect 14643 8134 21304 8186
rect 21356 8134 21368 8186
rect 21420 8134 21432 8186
rect 21484 8134 21496 8186
rect 21548 8134 21560 8186
rect 21612 8134 28273 8186
rect 28325 8134 28337 8186
rect 28389 8134 28401 8186
rect 28453 8134 28465 8186
rect 28517 8134 28529 8186
rect 28581 8134 28587 8186
rect 552 8112 28587 8134
rect 552 7642 28428 7664
rect 552 7590 3882 7642
rect 3934 7590 3946 7642
rect 3998 7590 4010 7642
rect 4062 7590 4074 7642
rect 4126 7590 4138 7642
rect 4190 7590 10851 7642
rect 10903 7590 10915 7642
rect 10967 7590 10979 7642
rect 11031 7590 11043 7642
rect 11095 7590 11107 7642
rect 11159 7590 17820 7642
rect 17872 7590 17884 7642
rect 17936 7590 17948 7642
rect 18000 7590 18012 7642
rect 18064 7590 18076 7642
rect 18128 7590 24789 7642
rect 24841 7590 24853 7642
rect 24905 7590 24917 7642
rect 24969 7590 24981 7642
rect 25033 7590 25045 7642
rect 25097 7590 28428 7642
rect 552 7568 28428 7590
rect 552 7098 28587 7120
rect 552 7046 7366 7098
rect 7418 7046 7430 7098
rect 7482 7046 7494 7098
rect 7546 7046 7558 7098
rect 7610 7046 7622 7098
rect 7674 7046 14335 7098
rect 14387 7046 14399 7098
rect 14451 7046 14463 7098
rect 14515 7046 14527 7098
rect 14579 7046 14591 7098
rect 14643 7046 21304 7098
rect 21356 7046 21368 7098
rect 21420 7046 21432 7098
rect 21484 7046 21496 7098
rect 21548 7046 21560 7098
rect 21612 7046 28273 7098
rect 28325 7046 28337 7098
rect 28389 7046 28401 7098
rect 28453 7046 28465 7098
rect 28517 7046 28529 7098
rect 28581 7046 28587 7098
rect 552 7024 28587 7046
rect 552 6554 28428 6576
rect 552 6502 3882 6554
rect 3934 6502 3946 6554
rect 3998 6502 4010 6554
rect 4062 6502 4074 6554
rect 4126 6502 4138 6554
rect 4190 6502 10851 6554
rect 10903 6502 10915 6554
rect 10967 6502 10979 6554
rect 11031 6502 11043 6554
rect 11095 6502 11107 6554
rect 11159 6502 17820 6554
rect 17872 6502 17884 6554
rect 17936 6502 17948 6554
rect 18000 6502 18012 6554
rect 18064 6502 18076 6554
rect 18128 6502 24789 6554
rect 24841 6502 24853 6554
rect 24905 6502 24917 6554
rect 24969 6502 24981 6554
rect 25033 6502 25045 6554
rect 25097 6502 28428 6554
rect 552 6480 28428 6502
rect 552 6010 28587 6032
rect 552 5958 7366 6010
rect 7418 5958 7430 6010
rect 7482 5958 7494 6010
rect 7546 5958 7558 6010
rect 7610 5958 7622 6010
rect 7674 5958 14335 6010
rect 14387 5958 14399 6010
rect 14451 5958 14463 6010
rect 14515 5958 14527 6010
rect 14579 5958 14591 6010
rect 14643 5958 21304 6010
rect 21356 5958 21368 6010
rect 21420 5958 21432 6010
rect 21484 5958 21496 6010
rect 21548 5958 21560 6010
rect 21612 5958 28273 6010
rect 28325 5958 28337 6010
rect 28389 5958 28401 6010
rect 28453 5958 28465 6010
rect 28517 5958 28529 6010
rect 28581 5958 28587 6010
rect 552 5936 28587 5958
rect 552 5466 28428 5488
rect 552 5414 3882 5466
rect 3934 5414 3946 5466
rect 3998 5414 4010 5466
rect 4062 5414 4074 5466
rect 4126 5414 4138 5466
rect 4190 5414 10851 5466
rect 10903 5414 10915 5466
rect 10967 5414 10979 5466
rect 11031 5414 11043 5466
rect 11095 5414 11107 5466
rect 11159 5414 17820 5466
rect 17872 5414 17884 5466
rect 17936 5414 17948 5466
rect 18000 5414 18012 5466
rect 18064 5414 18076 5466
rect 18128 5414 24789 5466
rect 24841 5414 24853 5466
rect 24905 5414 24917 5466
rect 24969 5414 24981 5466
rect 25033 5414 25045 5466
rect 25097 5414 28428 5466
rect 552 5392 28428 5414
rect 552 4922 28587 4944
rect 552 4870 7366 4922
rect 7418 4870 7430 4922
rect 7482 4870 7494 4922
rect 7546 4870 7558 4922
rect 7610 4870 7622 4922
rect 7674 4870 14335 4922
rect 14387 4870 14399 4922
rect 14451 4870 14463 4922
rect 14515 4870 14527 4922
rect 14579 4870 14591 4922
rect 14643 4870 21304 4922
rect 21356 4870 21368 4922
rect 21420 4870 21432 4922
rect 21484 4870 21496 4922
rect 21548 4870 21560 4922
rect 21612 4870 28273 4922
rect 28325 4870 28337 4922
rect 28389 4870 28401 4922
rect 28453 4870 28465 4922
rect 28517 4870 28529 4922
rect 28581 4870 28587 4922
rect 552 4848 28587 4870
rect 552 4378 28428 4400
rect 552 4326 3882 4378
rect 3934 4326 3946 4378
rect 3998 4326 4010 4378
rect 4062 4326 4074 4378
rect 4126 4326 4138 4378
rect 4190 4326 10851 4378
rect 10903 4326 10915 4378
rect 10967 4326 10979 4378
rect 11031 4326 11043 4378
rect 11095 4326 11107 4378
rect 11159 4326 17820 4378
rect 17872 4326 17884 4378
rect 17936 4326 17948 4378
rect 18000 4326 18012 4378
rect 18064 4326 18076 4378
rect 18128 4326 24789 4378
rect 24841 4326 24853 4378
rect 24905 4326 24917 4378
rect 24969 4326 24981 4378
rect 25033 4326 25045 4378
rect 25097 4326 28428 4378
rect 552 4304 28428 4326
rect 552 3834 28587 3856
rect 552 3782 7366 3834
rect 7418 3782 7430 3834
rect 7482 3782 7494 3834
rect 7546 3782 7558 3834
rect 7610 3782 7622 3834
rect 7674 3782 14335 3834
rect 14387 3782 14399 3834
rect 14451 3782 14463 3834
rect 14515 3782 14527 3834
rect 14579 3782 14591 3834
rect 14643 3782 21304 3834
rect 21356 3782 21368 3834
rect 21420 3782 21432 3834
rect 21484 3782 21496 3834
rect 21548 3782 21560 3834
rect 21612 3782 28273 3834
rect 28325 3782 28337 3834
rect 28389 3782 28401 3834
rect 28453 3782 28465 3834
rect 28517 3782 28529 3834
rect 28581 3782 28587 3834
rect 552 3760 28587 3782
rect 552 3290 28428 3312
rect 552 3238 3882 3290
rect 3934 3238 3946 3290
rect 3998 3238 4010 3290
rect 4062 3238 4074 3290
rect 4126 3238 4138 3290
rect 4190 3238 10851 3290
rect 10903 3238 10915 3290
rect 10967 3238 10979 3290
rect 11031 3238 11043 3290
rect 11095 3238 11107 3290
rect 11159 3238 17820 3290
rect 17872 3238 17884 3290
rect 17936 3238 17948 3290
rect 18000 3238 18012 3290
rect 18064 3238 18076 3290
rect 18128 3238 24789 3290
rect 24841 3238 24853 3290
rect 24905 3238 24917 3290
rect 24969 3238 24981 3290
rect 25033 3238 25045 3290
rect 25097 3238 28428 3290
rect 552 3216 28428 3238
rect 552 2746 28587 2768
rect 552 2694 7366 2746
rect 7418 2694 7430 2746
rect 7482 2694 7494 2746
rect 7546 2694 7558 2746
rect 7610 2694 7622 2746
rect 7674 2694 14335 2746
rect 14387 2694 14399 2746
rect 14451 2694 14463 2746
rect 14515 2694 14527 2746
rect 14579 2694 14591 2746
rect 14643 2694 21304 2746
rect 21356 2694 21368 2746
rect 21420 2694 21432 2746
rect 21484 2694 21496 2746
rect 21548 2694 21560 2746
rect 21612 2694 28273 2746
rect 28325 2694 28337 2746
rect 28389 2694 28401 2746
rect 28453 2694 28465 2746
rect 28517 2694 28529 2746
rect 28581 2694 28587 2746
rect 552 2672 28587 2694
rect 552 2202 28428 2224
rect 552 2150 3882 2202
rect 3934 2150 3946 2202
rect 3998 2150 4010 2202
rect 4062 2150 4074 2202
rect 4126 2150 4138 2202
rect 4190 2150 10851 2202
rect 10903 2150 10915 2202
rect 10967 2150 10979 2202
rect 11031 2150 11043 2202
rect 11095 2150 11107 2202
rect 11159 2150 17820 2202
rect 17872 2150 17884 2202
rect 17936 2150 17948 2202
rect 18000 2150 18012 2202
rect 18064 2150 18076 2202
rect 18128 2150 24789 2202
rect 24841 2150 24853 2202
rect 24905 2150 24917 2202
rect 24969 2150 24981 2202
rect 25033 2150 25045 2202
rect 25097 2150 28428 2202
rect 552 2128 28428 2150
rect 552 1658 28587 1680
rect 552 1606 7366 1658
rect 7418 1606 7430 1658
rect 7482 1606 7494 1658
rect 7546 1606 7558 1658
rect 7610 1606 7622 1658
rect 7674 1606 14335 1658
rect 14387 1606 14399 1658
rect 14451 1606 14463 1658
rect 14515 1606 14527 1658
rect 14579 1606 14591 1658
rect 14643 1606 21304 1658
rect 21356 1606 21368 1658
rect 21420 1606 21432 1658
rect 21484 1606 21496 1658
rect 21548 1606 21560 1658
rect 21612 1606 28273 1658
rect 28325 1606 28337 1658
rect 28389 1606 28401 1658
rect 28453 1606 28465 1658
rect 28517 1606 28529 1658
rect 28581 1606 28587 1658
rect 552 1584 28587 1606
rect 552 1114 28428 1136
rect 552 1062 3882 1114
rect 3934 1062 3946 1114
rect 3998 1062 4010 1114
rect 4062 1062 4074 1114
rect 4126 1062 4138 1114
rect 4190 1062 10851 1114
rect 10903 1062 10915 1114
rect 10967 1062 10979 1114
rect 11031 1062 11043 1114
rect 11095 1062 11107 1114
rect 11159 1062 17820 1114
rect 17872 1062 17884 1114
rect 17936 1062 17948 1114
rect 18000 1062 18012 1114
rect 18064 1062 18076 1114
rect 18128 1062 24789 1114
rect 24841 1062 24853 1114
rect 24905 1062 24917 1114
rect 24969 1062 24981 1114
rect 25033 1062 25045 1114
rect 25097 1062 28428 1114
rect 552 1040 28428 1062
rect 552 570 28587 592
rect 552 518 7366 570
rect 7418 518 7430 570
rect 7482 518 7494 570
rect 7546 518 7558 570
rect 7610 518 7622 570
rect 7674 518 14335 570
rect 14387 518 14399 570
rect 14451 518 14463 570
rect 14515 518 14527 570
rect 14579 518 14591 570
rect 14643 518 21304 570
rect 21356 518 21368 570
rect 21420 518 21432 570
rect 21484 518 21496 570
rect 21548 518 21560 570
rect 21612 518 28273 570
rect 28325 518 28337 570
rect 28389 518 28401 570
rect 28453 518 28465 570
rect 28517 518 28529 570
rect 28581 518 28587 570
rect 552 496 28587 518
<< via1 >>
rect 3882 28262 3934 28314
rect 3946 28262 3998 28314
rect 4010 28262 4062 28314
rect 4074 28262 4126 28314
rect 4138 28262 4190 28314
rect 10851 28262 10903 28314
rect 10915 28262 10967 28314
rect 10979 28262 11031 28314
rect 11043 28262 11095 28314
rect 11107 28262 11159 28314
rect 17820 28262 17872 28314
rect 17884 28262 17936 28314
rect 17948 28262 18000 28314
rect 18012 28262 18064 28314
rect 18076 28262 18128 28314
rect 24789 28262 24841 28314
rect 24853 28262 24905 28314
rect 24917 28262 24969 28314
rect 24981 28262 25033 28314
rect 25045 28262 25097 28314
rect 11428 28160 11480 28212
rect 19524 28160 19576 28212
rect 11152 27999 11204 28008
rect 11152 27965 11161 27999
rect 11161 27965 11195 27999
rect 11195 27965 11204 27999
rect 11152 27956 11204 27965
rect 15660 27999 15712 28008
rect 15660 27965 15669 27999
rect 15669 27965 15703 27999
rect 15703 27965 15712 27999
rect 15660 27956 15712 27965
rect 17500 27956 17552 28008
rect 19248 27999 19300 28008
rect 19248 27965 19257 27999
rect 19257 27965 19291 27999
rect 19291 27965 19300 27999
rect 19248 27956 19300 27965
rect 16212 27820 16264 27872
rect 18144 27820 18196 27872
rect 19892 27863 19944 27872
rect 19892 27829 19901 27863
rect 19901 27829 19935 27863
rect 19935 27829 19944 27863
rect 19892 27820 19944 27829
rect 20076 27863 20128 27872
rect 20076 27829 20085 27863
rect 20085 27829 20119 27863
rect 20119 27829 20128 27863
rect 20076 27820 20128 27829
rect 21548 27956 21600 28008
rect 23572 27956 23624 28008
rect 25596 27956 25648 28008
rect 21640 27863 21692 27872
rect 21640 27829 21649 27863
rect 21649 27829 21683 27863
rect 21683 27829 21692 27863
rect 21640 27820 21692 27829
rect 23848 27863 23900 27872
rect 23848 27829 23857 27863
rect 23857 27829 23891 27863
rect 23891 27829 23900 27863
rect 23848 27820 23900 27829
rect 25872 27863 25924 27872
rect 25872 27829 25881 27863
rect 25881 27829 25915 27863
rect 25915 27829 25924 27863
rect 25872 27820 25924 27829
rect 7366 27718 7418 27770
rect 7430 27718 7482 27770
rect 7494 27718 7546 27770
rect 7558 27718 7610 27770
rect 7622 27718 7674 27770
rect 14335 27718 14387 27770
rect 14399 27718 14451 27770
rect 14463 27718 14515 27770
rect 14527 27718 14579 27770
rect 14591 27718 14643 27770
rect 21304 27718 21356 27770
rect 21368 27718 21420 27770
rect 21432 27718 21484 27770
rect 21496 27718 21548 27770
rect 21560 27718 21612 27770
rect 28273 27718 28325 27770
rect 28337 27718 28389 27770
rect 28401 27718 28453 27770
rect 28465 27718 28517 27770
rect 28529 27718 28581 27770
rect 1308 27548 1360 27600
rect 3332 27548 3384 27600
rect 5356 27548 5408 27600
rect 2228 27480 2280 27532
rect 2596 27523 2648 27532
rect 2596 27489 2630 27523
rect 2630 27489 2648 27523
rect 2596 27480 2648 27489
rect 2320 27455 2372 27464
rect 2320 27421 2329 27455
rect 2329 27421 2363 27455
rect 2363 27421 2372 27455
rect 2320 27412 2372 27421
rect 4344 27412 4396 27464
rect 4896 27523 4948 27532
rect 4896 27489 4905 27523
rect 4905 27489 4939 27523
rect 4939 27489 4948 27523
rect 4896 27480 4948 27489
rect 5540 27523 5592 27532
rect 5540 27489 5549 27523
rect 5549 27489 5583 27523
rect 5583 27489 5592 27523
rect 5540 27480 5592 27489
rect 5908 27480 5960 27532
rect 7012 27480 7064 27532
rect 6092 27412 6144 27464
rect 6920 27344 6972 27396
rect 7288 27344 7340 27396
rect 7932 27480 7984 27532
rect 8944 27523 8996 27532
rect 8944 27489 8953 27523
rect 8953 27489 8987 27523
rect 8987 27489 8996 27523
rect 8944 27480 8996 27489
rect 9496 27480 9548 27532
rect 9956 27480 10008 27532
rect 11244 27480 11296 27532
rect 7840 27412 7892 27464
rect 11152 27344 11204 27396
rect 13268 27480 13320 27532
rect 15016 27591 15068 27600
rect 15016 27557 15025 27591
rect 15025 27557 15059 27591
rect 15059 27557 15068 27591
rect 15016 27548 15068 27557
rect 15660 27616 15712 27668
rect 19248 27616 19300 27668
rect 21640 27616 21692 27668
rect 15476 27548 15528 27600
rect 15200 27480 15252 27532
rect 16212 27480 16264 27532
rect 19892 27548 19944 27600
rect 18328 27480 18380 27532
rect 16120 27455 16172 27464
rect 16120 27421 16129 27455
rect 16129 27421 16163 27455
rect 16163 27421 16172 27455
rect 16120 27412 16172 27421
rect 14188 27344 14240 27396
rect 3700 27319 3752 27328
rect 3700 27285 3709 27319
rect 3709 27285 3743 27319
rect 3743 27285 3752 27319
rect 3700 27276 3752 27285
rect 4436 27319 4488 27328
rect 4436 27285 4445 27319
rect 4445 27285 4479 27319
rect 4479 27285 4488 27319
rect 4436 27276 4488 27285
rect 4988 27319 5040 27328
rect 4988 27285 4997 27319
rect 4997 27285 5031 27319
rect 5031 27285 5040 27319
rect 4988 27276 5040 27285
rect 6000 27276 6052 27328
rect 7472 27276 7524 27328
rect 10692 27276 10744 27328
rect 13452 27276 13504 27328
rect 14832 27276 14884 27328
rect 15108 27276 15160 27328
rect 22836 27480 22888 27532
rect 23296 27523 23348 27532
rect 23296 27489 23330 27523
rect 23330 27489 23348 27523
rect 23296 27480 23348 27489
rect 20628 27344 20680 27396
rect 19432 27276 19484 27328
rect 20720 27319 20772 27328
rect 20720 27285 20729 27319
rect 20729 27285 20763 27319
rect 20763 27285 20772 27319
rect 20720 27276 20772 27285
rect 20904 27276 20956 27328
rect 22928 27276 22980 27328
rect 24400 27319 24452 27328
rect 24400 27285 24409 27319
rect 24409 27285 24443 27319
rect 24443 27285 24452 27319
rect 24400 27276 24452 27285
rect 3882 27174 3934 27226
rect 3946 27174 3998 27226
rect 4010 27174 4062 27226
rect 4074 27174 4126 27226
rect 4138 27174 4190 27226
rect 10851 27174 10903 27226
rect 10915 27174 10967 27226
rect 10979 27174 11031 27226
rect 11043 27174 11095 27226
rect 11107 27174 11159 27226
rect 17820 27174 17872 27226
rect 17884 27174 17936 27226
rect 17948 27174 18000 27226
rect 18012 27174 18064 27226
rect 18076 27174 18128 27226
rect 24789 27174 24841 27226
rect 24853 27174 24905 27226
rect 24917 27174 24969 27226
rect 24981 27174 25033 27226
rect 25045 27174 25097 27226
rect 2596 27072 2648 27124
rect 4528 27072 4580 27124
rect 7840 27115 7892 27124
rect 7840 27081 7849 27115
rect 7849 27081 7883 27115
rect 7883 27081 7892 27115
rect 7840 27072 7892 27081
rect 9404 27072 9456 27124
rect 10692 27072 10744 27124
rect 3700 27004 3752 27056
rect 4896 27047 4948 27056
rect 3700 26868 3752 26920
rect 4896 27013 4905 27047
rect 4905 27013 4939 27047
rect 4939 27013 4948 27047
rect 4896 27004 4948 27013
rect 7748 27047 7800 27056
rect 7748 27013 7757 27047
rect 7757 27013 7791 27047
rect 7791 27013 7800 27047
rect 7748 27004 7800 27013
rect 6000 26911 6052 26920
rect 6000 26877 6018 26911
rect 6018 26877 6052 26911
rect 6000 26868 6052 26877
rect 6276 26911 6328 26920
rect 6276 26877 6285 26911
rect 6285 26877 6319 26911
rect 6319 26877 6328 26911
rect 6276 26868 6328 26877
rect 8760 26911 8812 26920
rect 8760 26877 8769 26911
rect 8769 26877 8803 26911
rect 8803 26877 8812 26911
rect 8760 26868 8812 26877
rect 13268 27072 13320 27124
rect 15016 27115 15068 27124
rect 15016 27081 15025 27115
rect 15025 27081 15059 27115
rect 15059 27081 15068 27115
rect 15016 27072 15068 27081
rect 18328 27115 18380 27124
rect 18328 27081 18337 27115
rect 18337 27081 18371 27115
rect 18371 27081 18380 27115
rect 18328 27072 18380 27081
rect 16764 27047 16816 27056
rect 16764 27013 16773 27047
rect 16773 27013 16807 27047
rect 16807 27013 16816 27047
rect 16764 27004 16816 27013
rect 11152 26936 11204 26988
rect 7288 26800 7340 26852
rect 12440 26911 12492 26920
rect 12440 26877 12449 26911
rect 12449 26877 12483 26911
rect 12483 26877 12492 26911
rect 12440 26868 12492 26877
rect 15200 26936 15252 26988
rect 12808 26911 12860 26920
rect 12808 26877 12817 26911
rect 12817 26877 12851 26911
rect 12851 26877 12860 26911
rect 12808 26868 12860 26877
rect 14740 26868 14792 26920
rect 15292 26911 15344 26920
rect 15292 26877 15301 26911
rect 15301 26877 15335 26911
rect 15335 26877 15344 26911
rect 15292 26868 15344 26877
rect 16672 26868 16724 26920
rect 18144 26868 18196 26920
rect 20444 26868 20496 26920
rect 20904 26911 20956 26920
rect 20904 26877 20938 26911
rect 20938 26877 20956 26911
rect 20904 26868 20956 26877
rect 4252 26775 4304 26784
rect 4252 26741 4261 26775
rect 4261 26741 4295 26775
rect 4295 26741 4304 26775
rect 4252 26732 4304 26741
rect 4344 26732 4396 26784
rect 7472 26732 7524 26784
rect 11428 26732 11480 26784
rect 11980 26775 12032 26784
rect 11980 26741 11989 26775
rect 11989 26741 12023 26775
rect 12023 26741 12032 26775
rect 11980 26732 12032 26741
rect 12624 26732 12676 26784
rect 13912 26732 13964 26784
rect 15108 26732 15160 26784
rect 16948 26775 17000 26784
rect 16948 26741 16957 26775
rect 16957 26741 16991 26775
rect 16991 26741 17000 26775
rect 16948 26732 17000 26741
rect 18144 26732 18196 26784
rect 19432 26800 19484 26852
rect 20076 26800 20128 26852
rect 22836 27072 22888 27124
rect 23296 27072 23348 27124
rect 24400 27072 24452 27124
rect 23848 26868 23900 26920
rect 23756 26800 23808 26852
rect 25872 26800 25924 26852
rect 20352 26732 20404 26784
rect 24216 26732 24268 26784
rect 7366 26630 7418 26682
rect 7430 26630 7482 26682
rect 7494 26630 7546 26682
rect 7558 26630 7610 26682
rect 7622 26630 7674 26682
rect 14335 26630 14387 26682
rect 14399 26630 14451 26682
rect 14463 26630 14515 26682
rect 14527 26630 14579 26682
rect 14591 26630 14643 26682
rect 21304 26630 21356 26682
rect 21368 26630 21420 26682
rect 21432 26630 21484 26682
rect 21496 26630 21548 26682
rect 21560 26630 21612 26682
rect 28273 26630 28325 26682
rect 28337 26630 28389 26682
rect 28401 26630 28453 26682
rect 28465 26630 28517 26682
rect 28529 26630 28581 26682
rect 4988 26528 5040 26580
rect 6092 26571 6144 26580
rect 6092 26537 6101 26571
rect 6101 26537 6135 26571
rect 6135 26537 6144 26571
rect 6092 26528 6144 26537
rect 7288 26528 7340 26580
rect 7564 26528 7616 26580
rect 7748 26571 7800 26580
rect 7748 26537 7757 26571
rect 7757 26537 7791 26571
rect 7791 26537 7800 26571
rect 7748 26528 7800 26537
rect 6828 26392 6880 26444
rect 4528 26324 4580 26376
rect 5908 26324 5960 26376
rect 6552 26367 6604 26376
rect 6552 26333 6561 26367
rect 6561 26333 6595 26367
rect 6595 26333 6604 26367
rect 6552 26324 6604 26333
rect 7564 26435 7616 26444
rect 7564 26401 7573 26435
rect 7573 26401 7607 26435
rect 7607 26401 7616 26435
rect 7564 26392 7616 26401
rect 7840 26435 7892 26444
rect 7840 26401 7849 26435
rect 7849 26401 7883 26435
rect 7883 26401 7892 26435
rect 7840 26392 7892 26401
rect 10048 26435 10100 26444
rect 10048 26401 10057 26435
rect 10057 26401 10091 26435
rect 10091 26401 10100 26435
rect 10048 26392 10100 26401
rect 6368 26256 6420 26308
rect 4436 26188 4488 26240
rect 11152 26528 11204 26580
rect 11980 26528 12032 26580
rect 12808 26528 12860 26580
rect 14188 26571 14240 26580
rect 14188 26537 14197 26571
rect 14197 26537 14231 26571
rect 14231 26537 14240 26571
rect 14188 26528 14240 26537
rect 14740 26571 14792 26580
rect 14740 26537 14749 26571
rect 14749 26537 14783 26571
rect 14783 26537 14792 26571
rect 14740 26528 14792 26537
rect 15292 26528 15344 26580
rect 16948 26528 17000 26580
rect 12256 26435 12308 26444
rect 12256 26401 12265 26435
rect 12265 26401 12299 26435
rect 12299 26401 12308 26435
rect 12256 26392 12308 26401
rect 12348 26392 12400 26444
rect 12532 26435 12584 26444
rect 12532 26401 12541 26435
rect 12541 26401 12575 26435
rect 12575 26401 12584 26435
rect 12532 26392 12584 26401
rect 12624 26435 12676 26444
rect 12624 26401 12633 26435
rect 12633 26401 12667 26435
rect 12667 26401 12676 26435
rect 12624 26392 12676 26401
rect 11612 26256 11664 26308
rect 11796 26256 11848 26308
rect 13912 26460 13964 26512
rect 13084 26256 13136 26308
rect 14004 26231 14056 26240
rect 14004 26197 14013 26231
rect 14013 26197 14047 26231
rect 14047 26197 14056 26231
rect 14740 26324 14792 26376
rect 16120 26392 16172 26444
rect 16580 26392 16632 26444
rect 20812 26435 20864 26444
rect 20812 26401 20830 26435
rect 20830 26401 20864 26435
rect 20812 26392 20864 26401
rect 15200 26324 15252 26376
rect 14004 26188 14056 26197
rect 16764 26188 16816 26240
rect 16856 26188 16908 26240
rect 19708 26299 19760 26308
rect 19708 26265 19717 26299
rect 19717 26265 19751 26299
rect 19751 26265 19760 26299
rect 19708 26256 19760 26265
rect 18236 26188 18288 26240
rect 20444 26188 20496 26240
rect 3882 26086 3934 26138
rect 3946 26086 3998 26138
rect 4010 26086 4062 26138
rect 4074 26086 4126 26138
rect 4138 26086 4190 26138
rect 10851 26086 10903 26138
rect 10915 26086 10967 26138
rect 10979 26086 11031 26138
rect 11043 26086 11095 26138
rect 11107 26086 11159 26138
rect 17820 26086 17872 26138
rect 17884 26086 17936 26138
rect 17948 26086 18000 26138
rect 18012 26086 18064 26138
rect 18076 26086 18128 26138
rect 24789 26086 24841 26138
rect 24853 26086 24905 26138
rect 24917 26086 24969 26138
rect 24981 26086 25033 26138
rect 25045 26086 25097 26138
rect 1400 25780 1452 25832
rect 2320 25780 2372 25832
rect 2412 25712 2464 25764
rect 6000 26027 6052 26036
rect 6000 25993 6009 26027
rect 6009 25993 6043 26027
rect 6043 25993 6052 26027
rect 6000 25984 6052 25993
rect 6552 25984 6604 26036
rect 7932 25984 7984 26036
rect 4712 25712 4764 25764
rect 6276 25780 6328 25832
rect 6736 25916 6788 25968
rect 7012 25916 7064 25968
rect 11336 25916 11388 25968
rect 12532 26027 12584 26036
rect 12532 25993 12541 26027
rect 12541 25993 12575 26027
rect 12575 25993 12584 26027
rect 12532 25984 12584 25993
rect 13084 26027 13136 26036
rect 13084 25993 13093 26027
rect 13093 25993 13127 26027
rect 13127 25993 13136 26027
rect 13084 25984 13136 25993
rect 13912 25916 13964 25968
rect 7932 25780 7984 25832
rect 8668 25780 8720 25832
rect 6828 25755 6880 25764
rect 6828 25721 6837 25755
rect 6837 25721 6871 25755
rect 6871 25721 6880 25755
rect 6828 25712 6880 25721
rect 7748 25712 7800 25764
rect 12256 25780 12308 25832
rect 3148 25644 3200 25696
rect 6000 25644 6052 25696
rect 6368 25644 6420 25696
rect 8760 25687 8812 25696
rect 8760 25653 8769 25687
rect 8769 25653 8803 25687
rect 8803 25653 8812 25687
rect 8760 25644 8812 25653
rect 11888 25644 11940 25696
rect 14832 25848 14884 25900
rect 16580 25984 16632 26036
rect 20812 25984 20864 26036
rect 12624 25712 12676 25764
rect 12716 25755 12768 25764
rect 12716 25721 12725 25755
rect 12725 25721 12759 25755
rect 12759 25721 12768 25755
rect 14004 25780 14056 25832
rect 14924 25823 14976 25832
rect 14924 25789 14933 25823
rect 14933 25789 14967 25823
rect 14967 25789 14976 25823
rect 14924 25780 14976 25789
rect 18144 25916 18196 25968
rect 18420 25780 18472 25832
rect 19984 25780 20036 25832
rect 20444 25848 20496 25900
rect 20352 25823 20404 25832
rect 20352 25789 20361 25823
rect 20361 25789 20395 25823
rect 20395 25789 20404 25823
rect 20352 25780 20404 25789
rect 22928 25780 22980 25832
rect 23848 25780 23900 25832
rect 12716 25712 12768 25721
rect 15292 25687 15344 25696
rect 15292 25653 15301 25687
rect 15301 25653 15335 25687
rect 15335 25653 15344 25687
rect 15292 25644 15344 25653
rect 21732 25712 21784 25764
rect 18696 25687 18748 25696
rect 18696 25653 18705 25687
rect 18705 25653 18739 25687
rect 18739 25653 18748 25687
rect 18696 25644 18748 25653
rect 22652 25687 22704 25696
rect 22652 25653 22661 25687
rect 22661 25653 22695 25687
rect 22695 25653 22704 25687
rect 22652 25644 22704 25653
rect 7366 25542 7418 25594
rect 7430 25542 7482 25594
rect 7494 25542 7546 25594
rect 7558 25542 7610 25594
rect 7622 25542 7674 25594
rect 14335 25542 14387 25594
rect 14399 25542 14451 25594
rect 14463 25542 14515 25594
rect 14527 25542 14579 25594
rect 14591 25542 14643 25594
rect 21304 25542 21356 25594
rect 21368 25542 21420 25594
rect 21432 25542 21484 25594
rect 21496 25542 21548 25594
rect 21560 25542 21612 25594
rect 28273 25542 28325 25594
rect 28337 25542 28389 25594
rect 28401 25542 28453 25594
rect 28465 25542 28517 25594
rect 28529 25542 28581 25594
rect 2412 25440 2464 25492
rect 3148 25483 3200 25492
rect 3148 25449 3157 25483
rect 3157 25449 3191 25483
rect 3191 25449 3200 25483
rect 3148 25440 3200 25449
rect 3700 25483 3752 25492
rect 3700 25449 3709 25483
rect 3709 25449 3743 25483
rect 3743 25449 3752 25483
rect 3700 25440 3752 25449
rect 4344 25440 4396 25492
rect 3332 25347 3384 25356
rect 3332 25313 3341 25347
rect 3341 25313 3375 25347
rect 3375 25313 3384 25347
rect 3332 25304 3384 25313
rect 4712 25483 4764 25492
rect 4712 25449 4721 25483
rect 4721 25449 4755 25483
rect 4755 25449 4764 25483
rect 4712 25440 4764 25449
rect 7932 25483 7984 25492
rect 7932 25449 7941 25483
rect 7941 25449 7975 25483
rect 7975 25449 7984 25483
rect 7932 25440 7984 25449
rect 8668 25440 8720 25492
rect 8760 25440 8812 25492
rect 8944 25440 8996 25492
rect 12256 25483 12308 25492
rect 12256 25449 12265 25483
rect 12265 25449 12299 25483
rect 12299 25449 12308 25483
rect 12256 25440 12308 25449
rect 4896 25347 4948 25356
rect 4896 25313 4905 25347
rect 4905 25313 4939 25347
rect 4939 25313 4948 25347
rect 4896 25304 4948 25313
rect 5448 25304 5500 25356
rect 3792 25236 3844 25288
rect 6644 25236 6696 25288
rect 8300 25347 8352 25356
rect 8300 25313 8309 25347
rect 8309 25313 8343 25347
rect 8343 25313 8352 25347
rect 8300 25304 8352 25313
rect 11612 25372 11664 25424
rect 14004 25372 14056 25424
rect 14372 25483 14424 25492
rect 14372 25449 14397 25483
rect 14397 25449 14424 25483
rect 14372 25440 14424 25449
rect 14832 25440 14884 25492
rect 15292 25483 15344 25492
rect 15292 25449 15301 25483
rect 15301 25449 15335 25483
rect 15335 25449 15344 25483
rect 15292 25440 15344 25449
rect 18420 25483 18472 25492
rect 18420 25449 18429 25483
rect 18429 25449 18463 25483
rect 18463 25449 18472 25483
rect 18420 25440 18472 25449
rect 21732 25483 21784 25492
rect 21732 25449 21741 25483
rect 21741 25449 21775 25483
rect 21775 25449 21784 25483
rect 21732 25440 21784 25449
rect 13728 25304 13780 25356
rect 8668 25279 8720 25288
rect 8668 25245 8677 25279
rect 8677 25245 8711 25279
rect 8711 25245 8720 25279
rect 8668 25236 8720 25245
rect 12532 25236 12584 25288
rect 16856 25372 16908 25424
rect 16764 25347 16816 25356
rect 16764 25313 16773 25347
rect 16773 25313 16807 25347
rect 16807 25313 16816 25347
rect 16764 25304 16816 25313
rect 18328 25372 18380 25424
rect 18604 25372 18656 25424
rect 19616 25347 19668 25356
rect 19616 25313 19650 25347
rect 19650 25313 19668 25347
rect 19616 25304 19668 25313
rect 23848 25372 23900 25424
rect 4344 25100 4396 25152
rect 5356 25100 5408 25152
rect 5448 25100 5500 25152
rect 9588 25100 9640 25152
rect 12716 25100 12768 25152
rect 13084 25100 13136 25152
rect 14556 25236 14608 25288
rect 14924 25236 14976 25288
rect 18696 25236 18748 25288
rect 21456 25347 21508 25356
rect 21456 25313 21465 25347
rect 21465 25313 21499 25347
rect 21499 25313 21508 25347
rect 21456 25304 21508 25313
rect 24216 25304 24268 25356
rect 14096 25100 14148 25152
rect 17132 25143 17184 25152
rect 17132 25109 17141 25143
rect 17141 25109 17175 25143
rect 17175 25109 17184 25143
rect 17132 25100 17184 25109
rect 18144 25100 18196 25152
rect 23204 25236 23256 25288
rect 19984 25100 20036 25152
rect 20996 25100 21048 25152
rect 22928 25143 22980 25152
rect 22928 25109 22937 25143
rect 22937 25109 22971 25143
rect 22971 25109 22980 25143
rect 22928 25100 22980 25109
rect 3882 24998 3934 25050
rect 3946 24998 3998 25050
rect 4010 24998 4062 25050
rect 4074 24998 4126 25050
rect 4138 24998 4190 25050
rect 10851 24998 10903 25050
rect 10915 24998 10967 25050
rect 10979 24998 11031 25050
rect 11043 24998 11095 25050
rect 11107 24998 11159 25050
rect 17820 24998 17872 25050
rect 17884 24998 17936 25050
rect 17948 24998 18000 25050
rect 18012 24998 18064 25050
rect 18076 24998 18128 25050
rect 24789 24998 24841 25050
rect 24853 24998 24905 25050
rect 24917 24998 24969 25050
rect 24981 24998 25033 25050
rect 25045 24998 25097 25050
rect 6644 24939 6696 24948
rect 3792 24828 3844 24880
rect 6644 24905 6653 24939
rect 6653 24905 6687 24939
rect 6687 24905 6696 24939
rect 6644 24896 6696 24905
rect 7012 24896 7064 24948
rect 9864 24896 9916 24948
rect 11888 24896 11940 24948
rect 12532 24939 12584 24948
rect 12532 24905 12541 24939
rect 12541 24905 12575 24939
rect 12575 24905 12584 24939
rect 12532 24896 12584 24905
rect 14188 24896 14240 24948
rect 14740 24896 14792 24948
rect 18328 24896 18380 24948
rect 19248 24896 19300 24948
rect 19616 24939 19668 24948
rect 19616 24905 19625 24939
rect 19625 24905 19659 24939
rect 19659 24905 19668 24939
rect 19616 24896 19668 24905
rect 21456 24896 21508 24948
rect 22652 24896 22704 24948
rect 11704 24828 11756 24880
rect 12348 24803 12400 24812
rect 12348 24769 12357 24803
rect 12357 24769 12391 24803
rect 12391 24769 12400 24803
rect 12348 24760 12400 24769
rect 14832 24871 14884 24880
rect 14832 24837 14841 24871
rect 14841 24837 14875 24871
rect 14875 24837 14884 24871
rect 14832 24828 14884 24837
rect 5908 24624 5960 24676
rect 7288 24556 7340 24608
rect 9496 24692 9548 24744
rect 9588 24692 9640 24744
rect 11060 24692 11112 24744
rect 12624 24692 12676 24744
rect 12716 24692 12768 24744
rect 13912 24735 13964 24744
rect 13912 24701 13921 24735
rect 13921 24701 13955 24735
rect 13955 24701 13964 24735
rect 13912 24692 13964 24701
rect 14004 24692 14056 24744
rect 10600 24624 10652 24676
rect 10784 24667 10836 24676
rect 10784 24633 10818 24667
rect 10818 24633 10836 24667
rect 10784 24624 10836 24633
rect 14096 24667 14148 24676
rect 14096 24633 14105 24667
rect 14105 24633 14139 24667
rect 14139 24633 14148 24667
rect 14096 24624 14148 24633
rect 14556 24667 14608 24676
rect 14556 24633 14565 24667
rect 14565 24633 14599 24667
rect 14599 24633 14608 24667
rect 14556 24624 14608 24633
rect 10416 24599 10468 24608
rect 10416 24565 10425 24599
rect 10425 24565 10459 24599
rect 10459 24565 10468 24599
rect 10416 24556 10468 24565
rect 10968 24556 11020 24608
rect 11704 24556 11756 24608
rect 14188 24556 14240 24608
rect 16120 24760 16172 24812
rect 20812 24760 20864 24812
rect 22008 24760 22060 24812
rect 18144 24624 18196 24676
rect 18512 24556 18564 24608
rect 18788 24556 18840 24608
rect 21824 24692 21876 24744
rect 19248 24556 19300 24608
rect 19616 24624 19668 24676
rect 19432 24556 19484 24608
rect 20628 24556 20680 24608
rect 21088 24599 21140 24608
rect 21088 24565 21097 24599
rect 21097 24565 21131 24599
rect 21131 24565 21140 24599
rect 21088 24556 21140 24565
rect 22652 24599 22704 24608
rect 22652 24565 22661 24599
rect 22661 24565 22695 24599
rect 22695 24565 22704 24599
rect 22652 24556 22704 24565
rect 7366 24454 7418 24506
rect 7430 24454 7482 24506
rect 7494 24454 7546 24506
rect 7558 24454 7610 24506
rect 7622 24454 7674 24506
rect 14335 24454 14387 24506
rect 14399 24454 14451 24506
rect 14463 24454 14515 24506
rect 14527 24454 14579 24506
rect 14591 24454 14643 24506
rect 21304 24454 21356 24506
rect 21368 24454 21420 24506
rect 21432 24454 21484 24506
rect 21496 24454 21548 24506
rect 21560 24454 21612 24506
rect 28273 24454 28325 24506
rect 28337 24454 28389 24506
rect 28401 24454 28453 24506
rect 28465 24454 28517 24506
rect 28529 24454 28581 24506
rect 1308 24259 1360 24268
rect 1308 24225 1317 24259
rect 1317 24225 1351 24259
rect 1351 24225 1360 24259
rect 1308 24216 1360 24225
rect 1400 24148 1452 24200
rect 2136 24216 2188 24268
rect 3516 24216 3568 24268
rect 3700 24216 3752 24268
rect 5356 24352 5408 24404
rect 7748 24352 7800 24404
rect 8668 24352 8720 24404
rect 9220 24352 9272 24404
rect 10416 24352 10468 24404
rect 10600 24352 10652 24404
rect 10784 24352 10836 24404
rect 5356 24148 5408 24200
rect 5908 24148 5960 24200
rect 6368 24216 6420 24268
rect 1124 24055 1176 24064
rect 1124 24021 1133 24055
rect 1133 24021 1167 24055
rect 1167 24021 1176 24055
rect 1124 24012 1176 24021
rect 4252 24012 4304 24064
rect 6184 24080 6236 24132
rect 7748 24216 7800 24268
rect 11152 24352 11204 24404
rect 12992 24352 13044 24404
rect 13912 24352 13964 24404
rect 14004 24352 14056 24404
rect 5264 24012 5316 24064
rect 5356 24055 5408 24064
rect 5356 24021 5365 24055
rect 5365 24021 5399 24055
rect 5399 24021 5408 24055
rect 5356 24012 5408 24021
rect 5816 24055 5868 24064
rect 5816 24021 5825 24055
rect 5825 24021 5859 24055
rect 5859 24021 5868 24055
rect 5816 24012 5868 24021
rect 6000 24012 6052 24064
rect 6092 24012 6144 24064
rect 6460 24055 6512 24064
rect 6460 24021 6469 24055
rect 6469 24021 6503 24055
rect 6503 24021 6512 24055
rect 6460 24012 6512 24021
rect 7288 24080 7340 24132
rect 11612 24259 11664 24268
rect 11612 24225 11621 24259
rect 11621 24225 11655 24259
rect 11655 24225 11664 24259
rect 11612 24216 11664 24225
rect 10968 24148 11020 24200
rect 11060 24148 11112 24200
rect 11152 24191 11204 24200
rect 11152 24157 11161 24191
rect 11161 24157 11195 24191
rect 11195 24157 11204 24191
rect 11152 24148 11204 24157
rect 11796 24259 11848 24268
rect 11796 24225 11805 24259
rect 11805 24225 11839 24259
rect 11839 24225 11848 24259
rect 11796 24216 11848 24225
rect 13084 24216 13136 24268
rect 14188 24352 14240 24404
rect 15568 24352 15620 24404
rect 7748 24012 7800 24064
rect 9036 24055 9088 24064
rect 9036 24021 9045 24055
rect 9045 24021 9079 24055
rect 9079 24021 9088 24055
rect 9036 24012 9088 24021
rect 9588 24123 9640 24132
rect 9588 24089 9597 24123
rect 9597 24089 9631 24123
rect 9631 24089 9640 24123
rect 9588 24080 9640 24089
rect 9772 24055 9824 24064
rect 9772 24021 9781 24055
rect 9781 24021 9815 24055
rect 9815 24021 9824 24055
rect 9772 24012 9824 24021
rect 10692 24012 10744 24064
rect 12072 24148 12124 24200
rect 12808 24148 12860 24200
rect 14096 24148 14148 24200
rect 11704 24080 11756 24132
rect 11796 24055 11848 24064
rect 11796 24021 11805 24055
rect 11805 24021 11839 24055
rect 11839 24021 11848 24055
rect 11796 24012 11848 24021
rect 13912 24012 13964 24064
rect 14648 24055 14700 24064
rect 14648 24021 14657 24055
rect 14657 24021 14691 24055
rect 14691 24021 14700 24055
rect 14648 24012 14700 24021
rect 16120 24259 16172 24268
rect 16120 24225 16129 24259
rect 16129 24225 16163 24259
rect 16163 24225 16172 24259
rect 16120 24216 16172 24225
rect 18052 24216 18104 24268
rect 18512 24259 18564 24268
rect 18512 24225 18521 24259
rect 18521 24225 18555 24259
rect 18555 24225 18564 24259
rect 18512 24216 18564 24225
rect 18604 24216 18656 24268
rect 18788 24395 18840 24404
rect 18788 24361 18797 24395
rect 18797 24361 18831 24395
rect 18831 24361 18840 24395
rect 18788 24352 18840 24361
rect 22468 24352 22520 24404
rect 22652 24352 22704 24404
rect 20352 24259 20404 24268
rect 20352 24225 20361 24259
rect 20361 24225 20395 24259
rect 20395 24225 20404 24259
rect 20352 24216 20404 24225
rect 21640 24216 21692 24268
rect 18788 24148 18840 24200
rect 19616 24148 19668 24200
rect 20536 24191 20588 24200
rect 20536 24157 20545 24191
rect 20545 24157 20579 24191
rect 20579 24157 20588 24191
rect 20536 24148 20588 24157
rect 20996 24080 21048 24132
rect 21824 24080 21876 24132
rect 22560 24259 22612 24268
rect 22560 24225 22569 24259
rect 22569 24225 22603 24259
rect 22603 24225 22612 24259
rect 22560 24216 22612 24225
rect 23204 24216 23256 24268
rect 22192 24148 22244 24200
rect 17040 24012 17092 24064
rect 17684 24012 17736 24064
rect 18328 24055 18380 24064
rect 18328 24021 18337 24055
rect 18337 24021 18371 24055
rect 18371 24021 18380 24055
rect 18328 24012 18380 24021
rect 18420 24055 18472 24064
rect 18420 24021 18429 24055
rect 18429 24021 18463 24055
rect 18463 24021 18472 24055
rect 18420 24012 18472 24021
rect 22468 24055 22520 24064
rect 22468 24021 22477 24055
rect 22477 24021 22511 24055
rect 22511 24021 22520 24055
rect 22468 24012 22520 24021
rect 23112 24080 23164 24132
rect 23572 24259 23624 24268
rect 23572 24225 23581 24259
rect 23581 24225 23615 24259
rect 23615 24225 23624 24259
rect 23572 24216 23624 24225
rect 24492 24216 24544 24268
rect 23848 24191 23900 24200
rect 23848 24157 23857 24191
rect 23857 24157 23891 24191
rect 23891 24157 23900 24191
rect 23848 24148 23900 24157
rect 23204 24055 23256 24064
rect 23204 24021 23213 24055
rect 23213 24021 23247 24055
rect 23247 24021 23256 24055
rect 23204 24012 23256 24021
rect 24216 24012 24268 24064
rect 24584 24012 24636 24064
rect 3882 23910 3934 23962
rect 3946 23910 3998 23962
rect 4010 23910 4062 23962
rect 4074 23910 4126 23962
rect 4138 23910 4190 23962
rect 10851 23910 10903 23962
rect 10915 23910 10967 23962
rect 10979 23910 11031 23962
rect 11043 23910 11095 23962
rect 11107 23910 11159 23962
rect 17820 23910 17872 23962
rect 17884 23910 17936 23962
rect 17948 23910 18000 23962
rect 18012 23910 18064 23962
rect 18076 23910 18128 23962
rect 24789 23910 24841 23962
rect 24853 23910 24905 23962
rect 24917 23910 24969 23962
rect 24981 23910 25033 23962
rect 25045 23910 25097 23962
rect 2136 23808 2188 23860
rect 3700 23808 3752 23860
rect 4252 23851 4304 23860
rect 4252 23817 4261 23851
rect 4261 23817 4295 23851
rect 4295 23817 4304 23851
rect 4252 23808 4304 23817
rect 4896 23808 4948 23860
rect 5816 23808 5868 23860
rect 6092 23808 6144 23860
rect 7288 23808 7340 23860
rect 9036 23808 9088 23860
rect 9128 23808 9180 23860
rect 11520 23808 11572 23860
rect 12716 23808 12768 23860
rect 14096 23808 14148 23860
rect 15660 23808 15712 23860
rect 16120 23851 16172 23860
rect 16120 23817 16129 23851
rect 16129 23817 16163 23851
rect 16163 23817 16172 23851
rect 16120 23808 16172 23817
rect 19984 23851 20036 23860
rect 19984 23817 19993 23851
rect 19993 23817 20027 23851
rect 20027 23817 20036 23851
rect 19984 23808 20036 23817
rect 20536 23851 20588 23860
rect 20536 23817 20545 23851
rect 20545 23817 20579 23851
rect 20579 23817 20588 23851
rect 20536 23808 20588 23817
rect 23572 23808 23624 23860
rect 24216 23808 24268 23860
rect 24492 23851 24544 23860
rect 24492 23817 24501 23851
rect 24501 23817 24535 23851
rect 24535 23817 24544 23851
rect 24492 23808 24544 23817
rect 9220 23740 9272 23792
rect 15568 23740 15620 23792
rect 16764 23740 16816 23792
rect 17684 23740 17736 23792
rect 1124 23579 1176 23588
rect 1124 23545 1158 23579
rect 1158 23545 1176 23579
rect 1124 23536 1176 23545
rect 1400 23604 1452 23656
rect 2872 23647 2924 23656
rect 2872 23613 2881 23647
rect 2881 23613 2915 23647
rect 2915 23613 2924 23647
rect 2872 23604 2924 23613
rect 4252 23604 4304 23656
rect 3700 23536 3752 23588
rect 5264 23604 5316 23656
rect 6460 23647 6512 23656
rect 6460 23613 6469 23647
rect 6469 23613 6503 23647
rect 6503 23613 6512 23647
rect 6460 23604 6512 23613
rect 9036 23604 9088 23656
rect 9772 23672 9824 23724
rect 12992 23672 13044 23724
rect 13820 23672 13872 23724
rect 9220 23604 9272 23656
rect 9404 23647 9456 23656
rect 9404 23613 9413 23647
rect 9413 23613 9447 23647
rect 9447 23613 9456 23647
rect 9404 23604 9456 23613
rect 1216 23468 1268 23520
rect 2412 23511 2464 23520
rect 2412 23477 2421 23511
rect 2421 23477 2455 23511
rect 2455 23477 2464 23511
rect 2412 23468 2464 23477
rect 3608 23468 3660 23520
rect 7840 23536 7892 23588
rect 13084 23604 13136 23656
rect 12808 23536 12860 23588
rect 12992 23536 13044 23588
rect 16856 23536 16908 23588
rect 17132 23604 17184 23656
rect 18788 23672 18840 23724
rect 20812 23715 20864 23724
rect 20812 23681 20821 23715
rect 20821 23681 20855 23715
rect 20855 23681 20864 23715
rect 21640 23715 21692 23724
rect 20812 23672 20864 23681
rect 21640 23681 21649 23715
rect 21649 23681 21683 23715
rect 21683 23681 21692 23715
rect 21640 23672 21692 23681
rect 18972 23604 19024 23656
rect 20996 23604 21048 23656
rect 21916 23604 21968 23656
rect 22468 23672 22520 23724
rect 17408 23579 17460 23588
rect 17408 23545 17417 23579
rect 17417 23545 17451 23579
rect 17451 23545 17460 23579
rect 17408 23536 17460 23545
rect 17868 23579 17920 23588
rect 17868 23545 17877 23579
rect 17877 23545 17911 23579
rect 17911 23545 17920 23579
rect 17868 23536 17920 23545
rect 8852 23468 8904 23520
rect 8944 23511 8996 23520
rect 8944 23477 8953 23511
rect 8953 23477 8987 23511
rect 8987 23477 8996 23511
rect 8944 23468 8996 23477
rect 9680 23468 9732 23520
rect 11612 23468 11664 23520
rect 12256 23468 12308 23520
rect 12532 23511 12584 23520
rect 12532 23477 12541 23511
rect 12541 23477 12575 23511
rect 12575 23477 12584 23511
rect 12532 23468 12584 23477
rect 13636 23468 13688 23520
rect 14188 23511 14240 23520
rect 14188 23477 14197 23511
rect 14197 23477 14231 23511
rect 14231 23477 14240 23511
rect 14188 23468 14240 23477
rect 22376 23647 22428 23656
rect 22376 23613 22385 23647
rect 22385 23613 22419 23647
rect 22419 23613 22428 23647
rect 22376 23604 22428 23613
rect 23204 23604 23256 23656
rect 23388 23604 23440 23656
rect 18144 23511 18196 23520
rect 18144 23477 18153 23511
rect 18153 23477 18187 23511
rect 18187 23477 18196 23511
rect 18144 23468 18196 23477
rect 22560 23468 22612 23520
rect 22652 23468 22704 23520
rect 24400 23647 24452 23656
rect 24400 23613 24409 23647
rect 24409 23613 24443 23647
rect 24443 23613 24452 23647
rect 24400 23604 24452 23613
rect 24584 23604 24636 23656
rect 7366 23366 7418 23418
rect 7430 23366 7482 23418
rect 7494 23366 7546 23418
rect 7558 23366 7610 23418
rect 7622 23366 7674 23418
rect 14335 23366 14387 23418
rect 14399 23366 14451 23418
rect 14463 23366 14515 23418
rect 14527 23366 14579 23418
rect 14591 23366 14643 23418
rect 21304 23366 21356 23418
rect 21368 23366 21420 23418
rect 21432 23366 21484 23418
rect 21496 23366 21548 23418
rect 21560 23366 21612 23418
rect 28273 23366 28325 23418
rect 28337 23366 28389 23418
rect 28401 23366 28453 23418
rect 28465 23366 28517 23418
rect 28529 23366 28581 23418
rect 1308 23264 1360 23316
rect 1768 23239 1820 23248
rect 1768 23205 1777 23239
rect 1777 23205 1811 23239
rect 1811 23205 1820 23239
rect 1768 23196 1820 23205
rect 2136 23196 2188 23248
rect 2412 23060 2464 23112
rect 3240 23239 3292 23248
rect 3240 23205 3265 23239
rect 3265 23205 3292 23239
rect 3240 23196 3292 23205
rect 3516 23307 3568 23316
rect 3516 23273 3525 23307
rect 3525 23273 3559 23307
rect 3559 23273 3568 23307
rect 3516 23264 3568 23273
rect 9404 23264 9456 23316
rect 4528 23196 4580 23248
rect 8760 23196 8812 23248
rect 9036 23196 9088 23248
rect 9680 23239 9732 23248
rect 4436 23171 4488 23180
rect 4436 23137 4445 23171
rect 4445 23137 4479 23171
rect 4479 23137 4488 23171
rect 4436 23128 4488 23137
rect 4620 23171 4672 23180
rect 4620 23137 4629 23171
rect 4629 23137 4663 23171
rect 4663 23137 4672 23171
rect 4620 23128 4672 23137
rect 5356 23128 5408 23180
rect 6644 23171 6696 23180
rect 6644 23137 6653 23171
rect 6653 23137 6687 23171
rect 6687 23137 6696 23171
rect 6644 23128 6696 23137
rect 7840 23128 7892 23180
rect 8668 23171 8720 23180
rect 8668 23137 8677 23171
rect 8677 23137 8711 23171
rect 8711 23137 8720 23171
rect 8668 23128 8720 23137
rect 6736 23103 6788 23112
rect 6736 23069 6745 23103
rect 6745 23069 6779 23103
rect 6779 23069 6788 23103
rect 6736 23060 6788 23069
rect 8300 23103 8352 23112
rect 8300 23069 8309 23103
rect 8309 23069 8343 23103
rect 8343 23069 8352 23103
rect 9680 23205 9714 23239
rect 9714 23205 9732 23239
rect 9680 23196 9732 23205
rect 9496 23128 9548 23180
rect 10692 23264 10744 23316
rect 11336 23264 11388 23316
rect 11888 23264 11940 23316
rect 12992 23264 13044 23316
rect 13820 23307 13872 23316
rect 13820 23273 13829 23307
rect 13829 23273 13863 23307
rect 13863 23273 13872 23307
rect 13820 23264 13872 23273
rect 14004 23264 14056 23316
rect 14096 23264 14148 23316
rect 11796 23128 11848 23180
rect 12164 23171 12216 23180
rect 12164 23137 12173 23171
rect 12173 23137 12207 23171
rect 12207 23137 12216 23171
rect 12164 23128 12216 23137
rect 12256 23171 12308 23180
rect 12256 23137 12265 23171
rect 12265 23137 12299 23171
rect 12299 23137 12308 23171
rect 12256 23128 12308 23137
rect 12348 23128 12400 23180
rect 12532 23128 12584 23180
rect 12900 23171 12952 23180
rect 12900 23137 12902 23171
rect 12902 23137 12936 23171
rect 12936 23137 12952 23171
rect 8300 23060 8352 23069
rect 11336 23103 11388 23112
rect 11336 23069 11345 23103
rect 11345 23069 11379 23103
rect 11379 23069 11388 23103
rect 11336 23060 11388 23069
rect 11704 23060 11756 23112
rect 12900 23128 12952 23137
rect 13084 23128 13136 23180
rect 13360 23171 13412 23180
rect 13360 23137 13369 23171
rect 13369 23137 13403 23171
rect 13403 23137 13412 23171
rect 15016 23196 15068 23248
rect 15292 23196 15344 23248
rect 15568 23196 15620 23248
rect 17868 23264 17920 23316
rect 13360 23128 13412 23137
rect 14832 23171 14884 23180
rect 14832 23137 14841 23171
rect 14841 23137 14875 23171
rect 14875 23137 14884 23171
rect 14832 23128 14884 23137
rect 2872 22992 2924 23044
rect 1676 22924 1728 22976
rect 3792 22924 3844 22976
rect 4528 22967 4580 22976
rect 4528 22933 4537 22967
rect 4537 22933 4571 22967
rect 4571 22933 4580 22967
rect 4528 22924 4580 22933
rect 8944 22924 8996 22976
rect 10048 22924 10100 22976
rect 10692 22924 10744 22976
rect 11612 22924 11664 22976
rect 12624 22992 12676 23044
rect 13176 23035 13228 23044
rect 13176 23001 13185 23035
rect 13185 23001 13219 23035
rect 13219 23001 13228 23035
rect 13176 22992 13228 23001
rect 14740 23060 14792 23112
rect 14004 22992 14056 23044
rect 16764 23171 16816 23180
rect 16764 23137 16773 23171
rect 16773 23137 16807 23171
rect 16807 23137 16816 23171
rect 16764 23128 16816 23137
rect 16856 23171 16908 23180
rect 16856 23137 16866 23171
rect 16866 23137 16900 23171
rect 16900 23137 16908 23171
rect 20996 23264 21048 23316
rect 21640 23307 21692 23316
rect 21640 23273 21649 23307
rect 21649 23273 21683 23307
rect 21683 23273 21692 23307
rect 21640 23264 21692 23273
rect 16856 23128 16908 23137
rect 17224 23171 17276 23180
rect 17224 23137 17233 23171
rect 17233 23137 17267 23171
rect 17267 23137 17276 23171
rect 17224 23128 17276 23137
rect 17316 23128 17368 23180
rect 18328 23128 18380 23180
rect 18420 23128 18472 23180
rect 18696 23171 18748 23180
rect 18696 23137 18705 23171
rect 18705 23137 18739 23171
rect 18739 23137 18748 23171
rect 18696 23128 18748 23137
rect 18788 23171 18840 23180
rect 18788 23137 18797 23171
rect 18797 23137 18831 23171
rect 18831 23137 18840 23171
rect 18788 23128 18840 23137
rect 18880 23171 18932 23180
rect 18880 23137 18925 23171
rect 18925 23137 18932 23171
rect 18880 23128 18932 23137
rect 19064 23171 19116 23180
rect 19064 23137 19073 23171
rect 19073 23137 19107 23171
rect 19107 23137 19116 23171
rect 19064 23128 19116 23137
rect 21916 23196 21968 23248
rect 18052 23060 18104 23112
rect 13636 22967 13688 22976
rect 13636 22933 13645 22967
rect 13645 22933 13679 22967
rect 13679 22933 13688 22967
rect 13636 22924 13688 22933
rect 13728 22967 13780 22976
rect 13728 22933 13737 22967
rect 13737 22933 13771 22967
rect 13771 22933 13780 22967
rect 13728 22924 13780 22933
rect 14464 22924 14516 22976
rect 21732 22992 21784 23044
rect 15108 22967 15160 22976
rect 15108 22933 15117 22967
rect 15117 22933 15151 22967
rect 15151 22933 15160 22967
rect 15108 22924 15160 22933
rect 15844 22967 15896 22976
rect 15844 22933 15853 22967
rect 15853 22933 15887 22967
rect 15887 22933 15896 22967
rect 15844 22924 15896 22933
rect 16856 22924 16908 22976
rect 17592 22967 17644 22976
rect 17592 22933 17601 22967
rect 17601 22933 17635 22967
rect 17635 22933 17644 22967
rect 17592 22924 17644 22933
rect 18144 22924 18196 22976
rect 18972 22924 19024 22976
rect 19156 22924 19208 22976
rect 21824 22967 21876 22976
rect 21824 22933 21833 22967
rect 21833 22933 21867 22967
rect 21867 22933 21876 22967
rect 21824 22924 21876 22933
rect 3882 22822 3934 22874
rect 3946 22822 3998 22874
rect 4010 22822 4062 22874
rect 4074 22822 4126 22874
rect 4138 22822 4190 22874
rect 10851 22822 10903 22874
rect 10915 22822 10967 22874
rect 10979 22822 11031 22874
rect 11043 22822 11095 22874
rect 11107 22822 11159 22874
rect 17820 22822 17872 22874
rect 17884 22822 17936 22874
rect 17948 22822 18000 22874
rect 18012 22822 18064 22874
rect 18076 22822 18128 22874
rect 24789 22822 24841 22874
rect 24853 22822 24905 22874
rect 24917 22822 24969 22874
rect 24981 22822 25033 22874
rect 25045 22822 25097 22874
rect 1768 22720 1820 22772
rect 2136 22763 2188 22772
rect 2136 22729 2145 22763
rect 2145 22729 2179 22763
rect 2179 22729 2188 22763
rect 2136 22720 2188 22729
rect 3240 22763 3292 22772
rect 3240 22729 3249 22763
rect 3249 22729 3283 22763
rect 3283 22729 3292 22763
rect 3240 22720 3292 22729
rect 3700 22720 3752 22772
rect 3792 22763 3844 22772
rect 3792 22729 3801 22763
rect 3801 22729 3835 22763
rect 3835 22729 3844 22763
rect 3792 22720 3844 22729
rect 4528 22720 4580 22772
rect 2412 22559 2464 22568
rect 2412 22525 2421 22559
rect 2421 22525 2455 22559
rect 2455 22525 2464 22559
rect 2412 22516 2464 22525
rect 3424 22559 3476 22568
rect 3424 22525 3433 22559
rect 3433 22525 3467 22559
rect 3467 22525 3476 22559
rect 3424 22516 3476 22525
rect 6000 22720 6052 22772
rect 6184 22720 6236 22772
rect 6920 22720 6972 22772
rect 8944 22720 8996 22772
rect 9864 22720 9916 22772
rect 10416 22720 10468 22772
rect 11428 22720 11480 22772
rect 11796 22720 11848 22772
rect 11888 22720 11940 22772
rect 12164 22763 12216 22772
rect 12164 22729 12173 22763
rect 12173 22729 12207 22763
rect 12207 22729 12216 22763
rect 12164 22720 12216 22729
rect 12624 22720 12676 22772
rect 6552 22652 6604 22704
rect 3608 22491 3660 22500
rect 3608 22457 3617 22491
rect 3617 22457 3651 22491
rect 3651 22457 3660 22491
rect 3608 22448 3660 22457
rect 3424 22380 3476 22432
rect 4344 22491 4396 22500
rect 4344 22457 4353 22491
rect 4353 22457 4387 22491
rect 4387 22457 4396 22491
rect 4344 22448 4396 22457
rect 4896 22516 4948 22568
rect 5356 22516 5408 22568
rect 6368 22584 6420 22636
rect 6460 22627 6512 22636
rect 6460 22593 6469 22627
rect 6469 22593 6503 22627
rect 6503 22593 6512 22627
rect 6460 22584 6512 22593
rect 11612 22652 11664 22704
rect 8024 22516 8076 22568
rect 8760 22627 8812 22636
rect 8760 22593 8769 22627
rect 8769 22593 8803 22627
rect 8803 22593 8812 22627
rect 8760 22584 8812 22593
rect 6736 22448 6788 22500
rect 7748 22448 7800 22500
rect 8300 22448 8352 22500
rect 9680 22516 9732 22568
rect 10692 22516 10744 22568
rect 12716 22584 12768 22636
rect 13636 22652 13688 22704
rect 14004 22652 14056 22704
rect 16396 22763 16448 22772
rect 16396 22729 16405 22763
rect 16405 22729 16439 22763
rect 16439 22729 16448 22763
rect 16396 22720 16448 22729
rect 19064 22720 19116 22772
rect 15292 22652 15344 22704
rect 12808 22559 12860 22568
rect 4620 22380 4672 22432
rect 5816 22380 5868 22432
rect 6000 22423 6052 22432
rect 6000 22389 6009 22423
rect 6009 22389 6043 22423
rect 6043 22389 6052 22423
rect 6000 22380 6052 22389
rect 8760 22380 8812 22432
rect 8944 22423 8996 22432
rect 8944 22389 8953 22423
rect 8953 22389 8987 22423
rect 8987 22389 8996 22423
rect 8944 22380 8996 22389
rect 12808 22525 12817 22559
rect 12817 22525 12851 22559
rect 12851 22525 12860 22559
rect 12808 22516 12860 22525
rect 11704 22448 11756 22500
rect 12532 22380 12584 22432
rect 13360 22448 13412 22500
rect 18972 22652 19024 22704
rect 20812 22720 20864 22772
rect 22376 22720 22428 22772
rect 19340 22652 19392 22704
rect 20260 22695 20312 22704
rect 20260 22661 20269 22695
rect 20269 22661 20303 22695
rect 20303 22661 20312 22695
rect 20260 22652 20312 22661
rect 15844 22627 15896 22636
rect 15844 22593 15853 22627
rect 15853 22593 15887 22627
rect 15887 22593 15896 22627
rect 15844 22584 15896 22593
rect 18236 22584 18288 22636
rect 19156 22627 19208 22636
rect 19156 22593 19165 22627
rect 19165 22593 19199 22627
rect 19199 22593 19208 22627
rect 19156 22584 19208 22593
rect 20720 22652 20772 22704
rect 21180 22695 21232 22704
rect 21180 22661 21189 22695
rect 21189 22661 21223 22695
rect 21223 22661 21232 22695
rect 21180 22652 21232 22661
rect 14188 22516 14240 22568
rect 14832 22516 14884 22568
rect 14464 22448 14516 22500
rect 12900 22380 12952 22432
rect 19064 22559 19116 22568
rect 19064 22525 19073 22559
rect 19073 22525 19107 22559
rect 19107 22525 19116 22559
rect 19064 22516 19116 22525
rect 18144 22448 18196 22500
rect 16488 22380 16540 22432
rect 20536 22516 20588 22568
rect 20260 22448 20312 22500
rect 20996 22559 21048 22568
rect 20996 22525 21005 22559
rect 21005 22525 21039 22559
rect 21039 22525 21048 22559
rect 20996 22516 21048 22525
rect 22192 22584 22244 22636
rect 22652 22584 22704 22636
rect 23296 22627 23348 22636
rect 23296 22593 23305 22627
rect 23305 22593 23339 22627
rect 23339 22593 23348 22627
rect 23296 22584 23348 22593
rect 23848 22627 23900 22636
rect 23848 22593 23857 22627
rect 23857 22593 23891 22627
rect 23891 22593 23900 22627
rect 23848 22584 23900 22593
rect 22560 22559 22612 22568
rect 22560 22525 22569 22559
rect 22569 22525 22603 22559
rect 22603 22525 22612 22559
rect 22560 22516 22612 22525
rect 23480 22559 23532 22568
rect 23480 22525 23489 22559
rect 23489 22525 23523 22559
rect 23523 22525 23532 22559
rect 23480 22516 23532 22525
rect 23112 22448 23164 22500
rect 24308 22448 24360 22500
rect 20536 22380 20588 22432
rect 21640 22380 21692 22432
rect 22100 22423 22152 22432
rect 22100 22389 22109 22423
rect 22109 22389 22143 22423
rect 22143 22389 22152 22423
rect 22100 22380 22152 22389
rect 22284 22380 22336 22432
rect 23664 22423 23716 22432
rect 23664 22389 23673 22423
rect 23673 22389 23707 22423
rect 23707 22389 23716 22423
rect 23664 22380 23716 22389
rect 25228 22423 25280 22432
rect 25228 22389 25237 22423
rect 25237 22389 25271 22423
rect 25271 22389 25280 22423
rect 25228 22380 25280 22389
rect 7366 22278 7418 22330
rect 7430 22278 7482 22330
rect 7494 22278 7546 22330
rect 7558 22278 7610 22330
rect 7622 22278 7674 22330
rect 14335 22278 14387 22330
rect 14399 22278 14451 22330
rect 14463 22278 14515 22330
rect 14527 22278 14579 22330
rect 14591 22278 14643 22330
rect 21304 22278 21356 22330
rect 21368 22278 21420 22330
rect 21432 22278 21484 22330
rect 21496 22278 21548 22330
rect 21560 22278 21612 22330
rect 28273 22278 28325 22330
rect 28337 22278 28389 22330
rect 28401 22278 28453 22330
rect 28465 22278 28517 22330
rect 28529 22278 28581 22330
rect 4896 22176 4948 22228
rect 5816 22176 5868 22228
rect 6460 22176 6512 22228
rect 8944 22176 8996 22228
rect 4436 22151 4488 22160
rect 4436 22117 4445 22151
rect 4445 22117 4479 22151
rect 4479 22117 4488 22151
rect 4436 22108 4488 22117
rect 5356 22108 5408 22160
rect 1492 22083 1544 22092
rect 1492 22049 1501 22083
rect 1501 22049 1535 22083
rect 1535 22049 1544 22083
rect 1492 22040 1544 22049
rect 1860 22040 1912 22092
rect 3424 21972 3476 22024
rect 6736 22040 6788 22092
rect 8484 22083 8536 22092
rect 8484 22049 8493 22083
rect 8493 22049 8527 22083
rect 8527 22049 8536 22083
rect 8484 22040 8536 22049
rect 9680 22108 9732 22160
rect 10600 22151 10652 22160
rect 10600 22117 10609 22151
rect 10609 22117 10643 22151
rect 10643 22117 10652 22151
rect 10600 22108 10652 22117
rect 9588 22083 9640 22092
rect 9588 22049 9597 22083
rect 9597 22049 9631 22083
rect 9631 22049 9640 22083
rect 9588 22040 9640 22049
rect 10508 22083 10560 22092
rect 10508 22049 10517 22083
rect 10517 22049 10551 22083
rect 10551 22049 10560 22083
rect 10508 22040 10560 22049
rect 11060 22040 11112 22092
rect 12256 22108 12308 22160
rect 13360 22151 13412 22160
rect 13360 22117 13369 22151
rect 13369 22117 13403 22151
rect 13403 22117 13412 22151
rect 13360 22108 13412 22117
rect 13636 22108 13688 22160
rect 16120 22108 16172 22160
rect 17224 22108 17276 22160
rect 14740 22040 14792 22092
rect 6460 21904 6512 21956
rect 1768 21879 1820 21888
rect 1768 21845 1777 21879
rect 1777 21845 1811 21879
rect 1811 21845 1820 21879
rect 1768 21836 1820 21845
rect 2044 21879 2096 21888
rect 2044 21845 2053 21879
rect 2053 21845 2087 21879
rect 2087 21845 2096 21879
rect 2044 21836 2096 21845
rect 2412 21836 2464 21888
rect 6644 21836 6696 21888
rect 8300 21879 8352 21888
rect 8300 21845 8309 21879
rect 8309 21845 8343 21879
rect 8343 21845 8352 21879
rect 8300 21836 8352 21845
rect 12440 21972 12492 22024
rect 12624 21972 12676 22024
rect 15108 21972 15160 22024
rect 16488 22015 16540 22024
rect 16488 21981 16497 22015
rect 16497 21981 16531 22015
rect 16531 21981 16540 22015
rect 16488 21972 16540 21981
rect 9956 21904 10008 21956
rect 11152 21904 11204 21956
rect 11980 21904 12032 21956
rect 18880 22108 18932 22160
rect 19708 22176 19760 22228
rect 20996 22176 21048 22228
rect 22560 22176 22612 22228
rect 21732 22151 21784 22160
rect 21732 22117 21741 22151
rect 21741 22117 21775 22151
rect 21775 22117 21784 22151
rect 21732 22108 21784 22117
rect 19432 22040 19484 22092
rect 18788 22015 18840 22024
rect 18788 21981 18797 22015
rect 18797 21981 18831 22015
rect 18831 21981 18840 22015
rect 18788 21972 18840 21981
rect 20260 22040 20312 22092
rect 20536 22040 20588 22092
rect 22100 22108 22152 22160
rect 22284 22108 22336 22160
rect 23664 22176 23716 22228
rect 24308 22219 24360 22228
rect 24308 22185 24317 22219
rect 24317 22185 24351 22219
rect 24351 22185 24360 22219
rect 24308 22176 24360 22185
rect 22652 22083 22704 22092
rect 22652 22049 22661 22083
rect 22661 22049 22695 22083
rect 22695 22049 22704 22083
rect 22652 22040 22704 22049
rect 22928 22083 22980 22092
rect 22928 22049 22937 22083
rect 22937 22049 22971 22083
rect 22971 22049 22980 22083
rect 22928 22040 22980 22049
rect 20996 21972 21048 22024
rect 20352 21904 20404 21956
rect 21640 21904 21692 21956
rect 22468 21972 22520 22024
rect 23480 22083 23532 22092
rect 23480 22049 23489 22083
rect 23489 22049 23523 22083
rect 23523 22049 23532 22083
rect 23480 22040 23532 22049
rect 23572 21904 23624 21956
rect 8668 21836 8720 21888
rect 9036 21836 9088 21888
rect 9312 21836 9364 21888
rect 9864 21836 9916 21888
rect 11428 21836 11480 21888
rect 15108 21836 15160 21888
rect 16672 21836 16724 21888
rect 17684 21836 17736 21888
rect 20260 21836 20312 21888
rect 21732 21836 21784 21888
rect 22928 21836 22980 21888
rect 3882 21734 3934 21786
rect 3946 21734 3998 21786
rect 4010 21734 4062 21786
rect 4074 21734 4126 21786
rect 4138 21734 4190 21786
rect 10851 21734 10903 21786
rect 10915 21734 10967 21786
rect 10979 21734 11031 21786
rect 11043 21734 11095 21786
rect 11107 21734 11159 21786
rect 17820 21734 17872 21786
rect 17884 21734 17936 21786
rect 17948 21734 18000 21786
rect 18012 21734 18064 21786
rect 18076 21734 18128 21786
rect 24789 21734 24841 21786
rect 24853 21734 24905 21786
rect 24917 21734 24969 21786
rect 24981 21734 25033 21786
rect 25045 21734 25097 21786
rect 2412 21675 2464 21684
rect 2412 21641 2421 21675
rect 2421 21641 2455 21675
rect 2455 21641 2464 21675
rect 2412 21632 2464 21641
rect 6920 21632 6972 21684
rect 1124 21428 1176 21480
rect 1768 21428 1820 21480
rect 5172 21564 5224 21616
rect 5356 21564 5408 21616
rect 5540 21539 5592 21548
rect 2872 21335 2924 21344
rect 2872 21301 2881 21335
rect 2881 21301 2915 21335
rect 2915 21301 2924 21335
rect 2872 21292 2924 21301
rect 3056 21403 3108 21412
rect 3056 21369 3065 21403
rect 3065 21369 3099 21403
rect 3099 21369 3108 21403
rect 3056 21360 3108 21369
rect 5540 21505 5549 21539
rect 5549 21505 5583 21539
rect 5583 21505 5592 21539
rect 5540 21496 5592 21505
rect 5356 21428 5408 21480
rect 7012 21428 7064 21480
rect 7104 21471 7156 21480
rect 7104 21437 7113 21471
rect 7113 21437 7147 21471
rect 7147 21437 7156 21471
rect 7104 21428 7156 21437
rect 8300 21632 8352 21684
rect 9312 21632 9364 21684
rect 9588 21632 9640 21684
rect 14004 21632 14056 21684
rect 8024 21496 8076 21548
rect 7748 21471 7800 21480
rect 7748 21437 7757 21471
rect 7757 21437 7791 21471
rect 7791 21437 7800 21471
rect 7748 21428 7800 21437
rect 3332 21292 3384 21344
rect 5816 21403 5868 21412
rect 5816 21369 5850 21403
rect 5850 21369 5868 21403
rect 5816 21360 5868 21369
rect 4804 21335 4856 21344
rect 4804 21301 4813 21335
rect 4813 21301 4847 21335
rect 4847 21301 4856 21335
rect 4804 21292 4856 21301
rect 6736 21292 6788 21344
rect 8392 21428 8444 21480
rect 8668 21428 8720 21480
rect 9312 21496 9364 21548
rect 9036 21428 9088 21480
rect 9864 21496 9916 21548
rect 10048 21471 10100 21480
rect 10048 21437 10057 21471
rect 10057 21437 10091 21471
rect 10091 21437 10100 21471
rect 10048 21428 10100 21437
rect 10508 21471 10560 21480
rect 10508 21437 10517 21471
rect 10517 21437 10551 21471
rect 10551 21437 10560 21471
rect 10508 21428 10560 21437
rect 9588 21292 9640 21344
rect 10232 21360 10284 21412
rect 10324 21292 10376 21344
rect 11888 21607 11940 21616
rect 11888 21573 11897 21607
rect 11897 21573 11931 21607
rect 11931 21573 11940 21607
rect 11888 21564 11940 21573
rect 12072 21496 12124 21548
rect 15660 21632 15712 21684
rect 15844 21632 15896 21684
rect 17224 21632 17276 21684
rect 18880 21632 18932 21684
rect 21088 21632 21140 21684
rect 22744 21632 22796 21684
rect 22836 21632 22888 21684
rect 12716 21428 12768 21480
rect 11796 21292 11848 21344
rect 14096 21360 14148 21412
rect 15016 21428 15068 21480
rect 14832 21360 14884 21412
rect 22284 21564 22336 21616
rect 17684 21539 17736 21548
rect 17684 21505 17693 21539
rect 17693 21505 17727 21539
rect 17727 21505 17736 21539
rect 17684 21496 17736 21505
rect 16304 21471 16356 21480
rect 16304 21437 16313 21471
rect 16313 21437 16347 21471
rect 16347 21437 16356 21471
rect 16304 21428 16356 21437
rect 15844 21335 15896 21344
rect 15844 21301 15853 21335
rect 15853 21301 15887 21335
rect 15887 21301 15896 21335
rect 15844 21292 15896 21301
rect 17224 21471 17276 21480
rect 17224 21437 17233 21471
rect 17233 21437 17267 21471
rect 17267 21437 17276 21471
rect 17224 21428 17276 21437
rect 17592 21428 17644 21480
rect 18052 21471 18104 21480
rect 18052 21437 18061 21471
rect 18061 21437 18095 21471
rect 18095 21437 18104 21471
rect 18052 21428 18104 21437
rect 20720 21496 20772 21548
rect 18972 21471 19024 21480
rect 18972 21437 18981 21471
rect 18981 21437 19015 21471
rect 19015 21437 19024 21471
rect 18972 21428 19024 21437
rect 19340 21428 19392 21480
rect 16764 21292 16816 21344
rect 20352 21428 20404 21480
rect 19708 21360 19760 21412
rect 19984 21360 20036 21412
rect 20996 21428 21048 21480
rect 22652 21496 22704 21548
rect 22928 21496 22980 21548
rect 21640 21428 21692 21480
rect 22192 21471 22244 21480
rect 22192 21437 22201 21471
rect 22201 21437 22235 21471
rect 22235 21437 22244 21471
rect 22192 21428 22244 21437
rect 24308 21496 24360 21548
rect 25228 21428 25280 21480
rect 19524 21292 19576 21344
rect 20260 21292 20312 21344
rect 21916 21292 21968 21344
rect 23020 21335 23072 21344
rect 23020 21301 23029 21335
rect 23029 21301 23063 21335
rect 23063 21301 23072 21335
rect 23020 21292 23072 21301
rect 23848 21335 23900 21344
rect 23848 21301 23857 21335
rect 23857 21301 23891 21335
rect 23891 21301 23900 21335
rect 23848 21292 23900 21301
rect 7366 21190 7418 21242
rect 7430 21190 7482 21242
rect 7494 21190 7546 21242
rect 7558 21190 7610 21242
rect 7622 21190 7674 21242
rect 14335 21190 14387 21242
rect 14399 21190 14451 21242
rect 14463 21190 14515 21242
rect 14527 21190 14579 21242
rect 14591 21190 14643 21242
rect 21304 21190 21356 21242
rect 21368 21190 21420 21242
rect 21432 21190 21484 21242
rect 21496 21190 21548 21242
rect 21560 21190 21612 21242
rect 28273 21190 28325 21242
rect 28337 21190 28389 21242
rect 28401 21190 28453 21242
rect 28465 21190 28517 21242
rect 28529 21190 28581 21242
rect 1860 21088 1912 21140
rect 3056 21088 3108 21140
rect 5264 21088 5316 21140
rect 5540 21088 5592 21140
rect 9496 21088 9548 21140
rect 9772 21088 9824 21140
rect 10324 21088 10376 21140
rect 1676 20952 1728 21004
rect 2044 20995 2096 21004
rect 2044 20961 2053 20995
rect 2053 20961 2087 20995
rect 2087 20961 2096 20995
rect 2044 20952 2096 20961
rect 2872 20952 2924 21004
rect 4804 20952 4856 21004
rect 4988 20995 5040 21004
rect 4988 20961 4997 20995
rect 4997 20961 5031 20995
rect 5031 20961 5040 20995
rect 4988 20952 5040 20961
rect 9680 21063 9732 21072
rect 9680 21029 9689 21063
rect 9689 21029 9723 21063
rect 9723 21029 9732 21063
rect 9680 21020 9732 21029
rect 12532 21088 12584 21140
rect 13544 21088 13596 21140
rect 11520 21020 11572 21072
rect 11980 21063 12032 21072
rect 11980 21029 11989 21063
rect 11989 21029 12023 21063
rect 12023 21029 12032 21063
rect 11980 21020 12032 21029
rect 1492 20748 1544 20800
rect 5080 20884 5132 20936
rect 5448 20952 5500 21004
rect 6276 20952 6328 21004
rect 8208 20952 8260 21004
rect 10232 20952 10284 21004
rect 13912 21020 13964 21072
rect 12808 20995 12860 21004
rect 12808 20961 12842 20995
rect 12842 20961 12860 20995
rect 5540 20927 5592 20936
rect 5540 20893 5549 20927
rect 5549 20893 5583 20927
rect 5583 20893 5592 20927
rect 5540 20884 5592 20893
rect 9864 20927 9916 20936
rect 9864 20893 9873 20927
rect 9873 20893 9907 20927
rect 9907 20893 9916 20927
rect 9864 20884 9916 20893
rect 9956 20927 10008 20936
rect 9956 20893 9965 20927
rect 9965 20893 9999 20927
rect 9999 20893 10008 20927
rect 9956 20884 10008 20893
rect 10048 20884 10100 20936
rect 3332 20816 3384 20868
rect 6092 20816 6144 20868
rect 11704 20884 11756 20936
rect 11980 20884 12032 20936
rect 12808 20952 12860 20961
rect 11244 20816 11296 20868
rect 3700 20748 3752 20800
rect 5632 20748 5684 20800
rect 6000 20748 6052 20800
rect 14188 20995 14240 21004
rect 14188 20961 14197 20995
rect 14197 20961 14231 20995
rect 14231 20961 14240 20995
rect 14188 20952 14240 20961
rect 14832 21131 14884 21140
rect 14832 21097 14841 21131
rect 14841 21097 14875 21131
rect 14875 21097 14884 21131
rect 14832 21088 14884 21097
rect 15844 21088 15896 21140
rect 16488 21088 16540 21140
rect 15016 20995 15068 21004
rect 15016 20961 15025 20995
rect 15025 20961 15059 20995
rect 15059 20961 15068 20995
rect 15016 20952 15068 20961
rect 17132 20952 17184 21004
rect 17592 20952 17644 21004
rect 17684 20952 17736 21004
rect 18972 21088 19024 21140
rect 20812 21088 20864 21140
rect 22744 21131 22796 21140
rect 22744 21097 22753 21131
rect 22753 21097 22787 21131
rect 22787 21097 22796 21131
rect 22744 21088 22796 21097
rect 23848 21088 23900 21140
rect 19524 21020 19576 21072
rect 19984 21063 20036 21072
rect 19984 21029 19994 21063
rect 19994 21029 20028 21063
rect 20028 21029 20036 21063
rect 19984 21020 20036 21029
rect 21732 21020 21784 21072
rect 16764 20884 16816 20936
rect 18972 20884 19024 20936
rect 19708 20952 19760 21004
rect 19432 20884 19484 20936
rect 20076 20995 20128 21004
rect 20076 20961 20111 20995
rect 20111 20961 20128 20995
rect 20076 20952 20128 20961
rect 20260 20995 20312 21004
rect 20260 20961 20269 20995
rect 20269 20961 20303 20995
rect 20303 20961 20312 20995
rect 20260 20952 20312 20961
rect 21824 20995 21876 21004
rect 21824 20961 21833 20995
rect 21833 20961 21867 20995
rect 21867 20961 21876 20995
rect 21824 20952 21876 20961
rect 22836 21020 22888 21072
rect 23020 20952 23072 21004
rect 22468 20816 22520 20868
rect 24400 20816 24452 20868
rect 14096 20748 14148 20800
rect 14740 20748 14792 20800
rect 17224 20748 17276 20800
rect 19248 20748 19300 20800
rect 20076 20748 20128 20800
rect 20904 20748 20956 20800
rect 22192 20748 22244 20800
rect 23388 20791 23440 20800
rect 23388 20757 23397 20791
rect 23397 20757 23431 20791
rect 23431 20757 23440 20791
rect 23388 20748 23440 20757
rect 3882 20646 3934 20698
rect 3946 20646 3998 20698
rect 4010 20646 4062 20698
rect 4074 20646 4126 20698
rect 4138 20646 4190 20698
rect 10851 20646 10903 20698
rect 10915 20646 10967 20698
rect 10979 20646 11031 20698
rect 11043 20646 11095 20698
rect 11107 20646 11159 20698
rect 17820 20646 17872 20698
rect 17884 20646 17936 20698
rect 17948 20646 18000 20698
rect 18012 20646 18064 20698
rect 18076 20646 18128 20698
rect 24789 20646 24841 20698
rect 24853 20646 24905 20698
rect 24917 20646 24969 20698
rect 24981 20646 25033 20698
rect 25045 20646 25097 20698
rect 5816 20587 5868 20596
rect 5816 20553 5825 20587
rect 5825 20553 5859 20587
rect 5859 20553 5868 20587
rect 5816 20544 5868 20553
rect 6828 20544 6880 20596
rect 9956 20544 10008 20596
rect 11060 20544 11112 20596
rect 12808 20587 12860 20596
rect 12808 20553 12817 20587
rect 12817 20553 12851 20587
rect 12851 20553 12860 20587
rect 12808 20544 12860 20553
rect 16304 20587 16356 20596
rect 16304 20553 16313 20587
rect 16313 20553 16347 20587
rect 16347 20553 16356 20587
rect 16304 20544 16356 20553
rect 16396 20544 16448 20596
rect 19340 20544 19392 20596
rect 19524 20544 19576 20596
rect 20904 20587 20956 20596
rect 20904 20553 20913 20587
rect 20913 20553 20947 20587
rect 20947 20553 20956 20587
rect 20904 20544 20956 20553
rect 21180 20544 21232 20596
rect 21824 20544 21876 20596
rect 22192 20587 22244 20596
rect 22192 20553 22201 20587
rect 22201 20553 22235 20587
rect 22235 20553 22244 20587
rect 22192 20544 22244 20553
rect 23388 20544 23440 20596
rect 6736 20519 6788 20528
rect 6736 20485 6745 20519
rect 6745 20485 6779 20519
rect 6779 20485 6788 20519
rect 6736 20476 6788 20485
rect 6092 20408 6144 20460
rect 7196 20408 7248 20460
rect 7288 20408 7340 20460
rect 8392 20451 8444 20460
rect 8392 20417 8401 20451
rect 8401 20417 8435 20451
rect 8435 20417 8444 20451
rect 8392 20408 8444 20417
rect 8484 20408 8536 20460
rect 12716 20476 12768 20528
rect 1952 20340 2004 20392
rect 5632 20340 5684 20392
rect 6000 20383 6052 20392
rect 6000 20349 6009 20383
rect 6009 20349 6043 20383
rect 6043 20349 6052 20383
rect 6000 20340 6052 20349
rect 6920 20383 6972 20392
rect 6920 20349 6929 20383
rect 6929 20349 6963 20383
rect 6963 20349 6972 20383
rect 6920 20340 6972 20349
rect 7104 20383 7156 20392
rect 7104 20349 7113 20383
rect 7113 20349 7147 20383
rect 7147 20349 7156 20383
rect 7104 20340 7156 20349
rect 9588 20451 9640 20460
rect 9588 20417 9597 20451
rect 9597 20417 9631 20451
rect 9631 20417 9640 20451
rect 9588 20408 9640 20417
rect 5356 20272 5408 20324
rect 5724 20272 5776 20324
rect 6736 20272 6788 20324
rect 9312 20383 9364 20392
rect 9312 20349 9321 20383
rect 9321 20349 9355 20383
rect 9355 20349 9364 20383
rect 9312 20340 9364 20349
rect 11244 20340 11296 20392
rect 12624 20408 12676 20460
rect 11980 20383 12032 20392
rect 11980 20349 11989 20383
rect 11989 20349 12023 20383
rect 12023 20349 12032 20383
rect 11980 20340 12032 20349
rect 12992 20340 13044 20392
rect 14004 20408 14056 20460
rect 14740 20408 14792 20460
rect 15384 20451 15436 20460
rect 15384 20417 15393 20451
rect 15393 20417 15427 20451
rect 15427 20417 15436 20451
rect 15384 20408 15436 20417
rect 13176 20340 13228 20392
rect 13636 20383 13688 20392
rect 13636 20349 13645 20383
rect 13645 20349 13679 20383
rect 13679 20349 13688 20383
rect 13636 20340 13688 20349
rect 11428 20272 11480 20324
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 4988 20204 5040 20256
rect 6092 20204 6144 20256
rect 7012 20247 7064 20256
rect 7012 20213 7021 20247
rect 7021 20213 7055 20247
rect 7055 20213 7064 20247
rect 7012 20204 7064 20213
rect 7196 20204 7248 20256
rect 11336 20247 11388 20256
rect 11336 20213 11345 20247
rect 11345 20213 11379 20247
rect 11379 20213 11388 20247
rect 11336 20204 11388 20213
rect 12164 20315 12216 20324
rect 12164 20281 12173 20315
rect 12173 20281 12207 20315
rect 12207 20281 12216 20315
rect 12164 20272 12216 20281
rect 16764 20451 16816 20460
rect 16764 20417 16773 20451
rect 16773 20417 16807 20451
rect 16807 20417 16816 20451
rect 16764 20408 16816 20417
rect 16948 20451 17000 20460
rect 16948 20417 16957 20451
rect 16957 20417 16991 20451
rect 16991 20417 17000 20451
rect 16948 20408 17000 20417
rect 17132 20408 17184 20460
rect 16580 20340 16632 20392
rect 18972 20272 19024 20324
rect 20536 20383 20588 20392
rect 20536 20349 20545 20383
rect 20545 20349 20579 20383
rect 20579 20349 20588 20383
rect 20536 20340 20588 20349
rect 20996 20383 21048 20392
rect 20996 20349 21005 20383
rect 21005 20349 21039 20383
rect 21039 20349 21048 20383
rect 20996 20340 21048 20349
rect 21732 20383 21784 20392
rect 21732 20349 21741 20383
rect 21741 20349 21775 20383
rect 21775 20349 21784 20383
rect 21732 20340 21784 20349
rect 22100 20383 22152 20392
rect 22100 20349 22109 20383
rect 22109 20349 22143 20383
rect 22143 20349 22152 20383
rect 22100 20340 22152 20349
rect 22468 20383 22520 20392
rect 22468 20349 22477 20383
rect 22477 20349 22511 20383
rect 22511 20349 22520 20383
rect 22468 20340 22520 20349
rect 23480 20340 23532 20392
rect 12348 20204 12400 20256
rect 12900 20204 12952 20256
rect 13176 20204 13228 20256
rect 14832 20247 14884 20256
rect 14832 20213 14841 20247
rect 14841 20213 14875 20247
rect 14875 20213 14884 20247
rect 14832 20204 14884 20213
rect 17224 20204 17276 20256
rect 18144 20204 18196 20256
rect 21640 20204 21692 20256
rect 22836 20204 22888 20256
rect 7366 20102 7418 20154
rect 7430 20102 7482 20154
rect 7494 20102 7546 20154
rect 7558 20102 7610 20154
rect 7622 20102 7674 20154
rect 14335 20102 14387 20154
rect 14399 20102 14451 20154
rect 14463 20102 14515 20154
rect 14527 20102 14579 20154
rect 14591 20102 14643 20154
rect 21304 20102 21356 20154
rect 21368 20102 21420 20154
rect 21432 20102 21484 20154
rect 21496 20102 21548 20154
rect 21560 20102 21612 20154
rect 28273 20102 28325 20154
rect 28337 20102 28389 20154
rect 28401 20102 28453 20154
rect 28465 20102 28517 20154
rect 28529 20102 28581 20154
rect 1584 19975 1636 19984
rect 1584 19941 1618 19975
rect 1618 19941 1636 19975
rect 1584 19932 1636 19941
rect 1124 19864 1176 19916
rect 1492 19660 1544 19712
rect 2872 19660 2924 19712
rect 3608 19932 3660 19984
rect 7012 20000 7064 20052
rect 4804 19864 4856 19916
rect 4988 19839 5040 19848
rect 4988 19805 4997 19839
rect 4997 19805 5031 19839
rect 5031 19805 5040 19839
rect 4988 19796 5040 19805
rect 5080 19839 5132 19848
rect 5080 19805 5089 19839
rect 5089 19805 5123 19839
rect 5123 19805 5132 19839
rect 5080 19796 5132 19805
rect 5724 19796 5776 19848
rect 6184 19864 6236 19916
rect 6736 19907 6788 19916
rect 6736 19873 6745 19907
rect 6745 19873 6779 19907
rect 6779 19873 6788 19907
rect 6736 19864 6788 19873
rect 6920 19864 6972 19916
rect 7380 19975 7432 19984
rect 7380 19941 7408 19975
rect 7408 19941 7432 19975
rect 9036 20000 9088 20052
rect 9312 20000 9364 20052
rect 11336 20000 11388 20052
rect 11980 20000 12032 20052
rect 12992 20000 13044 20052
rect 13268 20000 13320 20052
rect 13544 20043 13596 20052
rect 13544 20009 13553 20043
rect 13553 20009 13587 20043
rect 13587 20009 13596 20043
rect 13544 20000 13596 20009
rect 13636 20043 13688 20052
rect 13636 20009 13645 20043
rect 13645 20009 13679 20043
rect 13679 20009 13688 20043
rect 13636 20000 13688 20009
rect 14740 20000 14792 20052
rect 14924 20000 14976 20052
rect 15384 20000 15436 20052
rect 16396 20000 16448 20052
rect 16764 20000 16816 20052
rect 17224 20043 17276 20052
rect 17224 20009 17233 20043
rect 17233 20009 17267 20043
rect 17267 20009 17276 20043
rect 17224 20000 17276 20009
rect 20996 20000 21048 20052
rect 7380 19932 7432 19941
rect 8576 19932 8628 19984
rect 8116 19864 8168 19916
rect 7288 19796 7340 19848
rect 9772 19864 9824 19916
rect 9956 19907 10008 19916
rect 9956 19873 9965 19907
rect 9965 19873 9999 19907
rect 9999 19873 10008 19907
rect 9956 19864 10008 19873
rect 12808 19864 12860 19916
rect 16120 19932 16172 19984
rect 22100 20043 22152 20052
rect 22100 20009 22109 20043
rect 22109 20009 22143 20043
rect 22143 20009 22152 20043
rect 22100 20000 22152 20009
rect 23020 20000 23072 20052
rect 24308 20043 24360 20052
rect 24308 20009 24317 20043
rect 24317 20009 24351 20043
rect 24351 20009 24360 20043
rect 24308 20000 24360 20009
rect 21916 19975 21968 19984
rect 13176 19907 13228 19916
rect 13176 19873 13185 19907
rect 13185 19873 13219 19907
rect 13219 19873 13228 19907
rect 13176 19864 13228 19873
rect 13820 19864 13872 19916
rect 13912 19864 13964 19916
rect 14188 19864 14240 19916
rect 3792 19728 3844 19780
rect 4436 19660 4488 19712
rect 4528 19703 4580 19712
rect 4528 19669 4537 19703
rect 4537 19669 4571 19703
rect 4571 19669 4580 19703
rect 4528 19660 4580 19669
rect 5540 19660 5592 19712
rect 6460 19703 6512 19712
rect 6460 19669 6469 19703
rect 6469 19669 6503 19703
rect 6503 19669 6512 19703
rect 6460 19660 6512 19669
rect 6644 19660 6696 19712
rect 8024 19660 8076 19712
rect 10232 19660 10284 19712
rect 10324 19703 10376 19712
rect 10324 19669 10333 19703
rect 10333 19669 10367 19703
rect 10367 19669 10376 19703
rect 10324 19660 10376 19669
rect 12900 19796 12952 19848
rect 13636 19796 13688 19848
rect 13452 19728 13504 19780
rect 11244 19660 11296 19712
rect 12532 19660 12584 19712
rect 12992 19703 13044 19712
rect 12992 19669 13001 19703
rect 13001 19669 13035 19703
rect 13035 19669 13044 19703
rect 12992 19660 13044 19669
rect 13268 19703 13320 19712
rect 13268 19669 13277 19703
rect 13277 19669 13311 19703
rect 13311 19669 13320 19703
rect 13268 19660 13320 19669
rect 13636 19660 13688 19712
rect 19340 19796 19392 19848
rect 20076 19839 20128 19848
rect 20076 19805 20085 19839
rect 20085 19805 20119 19839
rect 20119 19805 20128 19839
rect 20076 19796 20128 19805
rect 21180 19864 21232 19916
rect 21640 19864 21692 19916
rect 21916 19941 21925 19975
rect 21925 19941 21959 19975
rect 21959 19941 21968 19975
rect 21916 19932 21968 19941
rect 22284 19864 22336 19916
rect 23204 19907 23256 19916
rect 23204 19873 23238 19907
rect 23238 19873 23256 19907
rect 23204 19864 23256 19873
rect 22928 19839 22980 19848
rect 22928 19805 22937 19839
rect 22937 19805 22971 19839
rect 22971 19805 22980 19839
rect 22928 19796 22980 19805
rect 18236 19660 18288 19712
rect 18880 19660 18932 19712
rect 21272 19703 21324 19712
rect 21272 19669 21281 19703
rect 21281 19669 21315 19703
rect 21315 19669 21324 19703
rect 21272 19660 21324 19669
rect 3882 19558 3934 19610
rect 3946 19558 3998 19610
rect 4010 19558 4062 19610
rect 4074 19558 4126 19610
rect 4138 19558 4190 19610
rect 10851 19558 10903 19610
rect 10915 19558 10967 19610
rect 10979 19558 11031 19610
rect 11043 19558 11095 19610
rect 11107 19558 11159 19610
rect 17820 19558 17872 19610
rect 17884 19558 17936 19610
rect 17948 19558 18000 19610
rect 18012 19558 18064 19610
rect 18076 19558 18128 19610
rect 24789 19558 24841 19610
rect 24853 19558 24905 19610
rect 24917 19558 24969 19610
rect 24981 19558 25033 19610
rect 25045 19558 25097 19610
rect 1676 19456 1728 19508
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 3700 19456 3752 19508
rect 4436 19456 4488 19508
rect 5724 19456 5776 19508
rect 1492 19388 1544 19440
rect 3608 19363 3660 19372
rect 3608 19329 3617 19363
rect 3617 19329 3651 19363
rect 3651 19329 3660 19363
rect 3608 19320 3660 19329
rect 2872 19227 2924 19236
rect 2872 19193 2881 19227
rect 2881 19193 2915 19227
rect 2915 19193 2924 19227
rect 2872 19184 2924 19193
rect 3792 19252 3844 19304
rect 2136 19116 2188 19168
rect 3976 19295 4028 19304
rect 3976 19261 3985 19295
rect 3985 19261 4019 19295
rect 4019 19261 4028 19295
rect 3976 19252 4028 19261
rect 5448 19252 5500 19304
rect 6460 19456 6512 19508
rect 6920 19499 6972 19508
rect 6920 19465 6929 19499
rect 6929 19465 6963 19499
rect 6963 19465 6972 19499
rect 6920 19456 6972 19465
rect 8116 19456 8168 19508
rect 8208 19456 8260 19508
rect 7380 19388 7432 19440
rect 16948 19456 17000 19508
rect 20076 19499 20128 19508
rect 20076 19465 20085 19499
rect 20085 19465 20119 19499
rect 20119 19465 20128 19499
rect 20076 19456 20128 19465
rect 21272 19456 21324 19508
rect 22100 19456 22152 19508
rect 23204 19499 23256 19508
rect 23204 19465 23213 19499
rect 23213 19465 23247 19499
rect 23247 19465 23256 19499
rect 23204 19456 23256 19465
rect 6184 19320 6236 19372
rect 8024 19320 8076 19372
rect 6828 19252 6880 19304
rect 4896 19184 4948 19236
rect 5080 19184 5132 19236
rect 9588 19388 9640 19440
rect 9956 19388 10008 19440
rect 10048 19431 10100 19440
rect 10048 19397 10057 19431
rect 10057 19397 10091 19431
rect 10091 19397 10100 19431
rect 10048 19388 10100 19397
rect 13176 19388 13228 19440
rect 13728 19388 13780 19440
rect 17408 19388 17460 19440
rect 20720 19431 20772 19440
rect 20720 19397 20729 19431
rect 20729 19397 20763 19431
rect 20763 19397 20772 19431
rect 20720 19388 20772 19397
rect 11244 19320 11296 19372
rect 9772 19252 9824 19304
rect 9956 19252 10008 19304
rect 12808 19320 12860 19372
rect 13544 19320 13596 19372
rect 15384 19252 15436 19304
rect 17408 19252 17460 19304
rect 17684 19252 17736 19304
rect 17960 19295 18012 19304
rect 17960 19261 17969 19295
rect 17969 19261 18003 19295
rect 18003 19261 18012 19295
rect 17960 19252 18012 19261
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 18236 19295 18288 19304
rect 18236 19261 18245 19295
rect 18245 19261 18279 19295
rect 18279 19261 18288 19295
rect 18236 19252 18288 19261
rect 18328 19295 18380 19304
rect 18328 19261 18337 19295
rect 18337 19261 18371 19295
rect 18371 19261 18380 19295
rect 18328 19252 18380 19261
rect 18512 19320 18564 19372
rect 20168 19320 20220 19372
rect 11980 19227 12032 19236
rect 11980 19193 12014 19227
rect 12014 19193 12032 19227
rect 11980 19184 12032 19193
rect 15016 19184 15068 19236
rect 20996 19295 21048 19304
rect 20996 19261 21005 19295
rect 21005 19261 21039 19295
rect 21039 19261 21048 19295
rect 20996 19252 21048 19261
rect 21548 19252 21600 19304
rect 22100 19295 22152 19304
rect 22100 19261 22109 19295
rect 22109 19261 22143 19295
rect 22143 19261 22152 19295
rect 22100 19252 22152 19261
rect 22284 19295 22336 19304
rect 22284 19261 22293 19295
rect 22293 19261 22327 19295
rect 22327 19261 22336 19295
rect 22284 19252 22336 19261
rect 22560 19295 22612 19304
rect 22560 19261 22569 19295
rect 22569 19261 22603 19295
rect 22603 19261 22612 19295
rect 22560 19252 22612 19261
rect 22836 19252 22888 19304
rect 6092 19159 6144 19168
rect 6092 19125 6119 19159
rect 6119 19125 6144 19159
rect 6092 19116 6144 19125
rect 6644 19116 6696 19168
rect 8392 19159 8444 19168
rect 8392 19125 8401 19159
rect 8401 19125 8435 19159
rect 8435 19125 8444 19159
rect 8392 19116 8444 19125
rect 8668 19116 8720 19168
rect 9036 19159 9088 19168
rect 9036 19125 9045 19159
rect 9045 19125 9079 19159
rect 9079 19125 9088 19159
rect 9036 19116 9088 19125
rect 10968 19116 11020 19168
rect 13360 19116 13412 19168
rect 14004 19116 14056 19168
rect 16580 19116 16632 19168
rect 21916 19184 21968 19236
rect 20444 19116 20496 19168
rect 21180 19116 21232 19168
rect 21640 19159 21692 19168
rect 21640 19125 21649 19159
rect 21649 19125 21683 19159
rect 21683 19125 21692 19159
rect 21640 19116 21692 19125
rect 7366 19014 7418 19066
rect 7430 19014 7482 19066
rect 7494 19014 7546 19066
rect 7558 19014 7610 19066
rect 7622 19014 7674 19066
rect 14335 19014 14387 19066
rect 14399 19014 14451 19066
rect 14463 19014 14515 19066
rect 14527 19014 14579 19066
rect 14591 19014 14643 19066
rect 21304 19014 21356 19066
rect 21368 19014 21420 19066
rect 21432 19014 21484 19066
rect 21496 19014 21548 19066
rect 21560 19014 21612 19066
rect 28273 19014 28325 19066
rect 28337 19014 28389 19066
rect 28401 19014 28453 19066
rect 28465 19014 28517 19066
rect 28529 19014 28581 19066
rect 3976 18912 4028 18964
rect 4528 18912 4580 18964
rect 4896 18955 4948 18964
rect 4896 18921 4905 18955
rect 4905 18921 4939 18955
rect 4939 18921 4948 18955
rect 4896 18912 4948 18921
rect 5448 18912 5500 18964
rect 8760 18912 8812 18964
rect 11796 18955 11848 18964
rect 11796 18921 11805 18955
rect 11805 18921 11839 18955
rect 11839 18921 11848 18955
rect 11796 18912 11848 18921
rect 11980 18955 12032 18964
rect 11980 18921 11989 18955
rect 11989 18921 12023 18955
rect 12023 18921 12032 18955
rect 11980 18912 12032 18921
rect 12992 18912 13044 18964
rect 3608 18819 3660 18828
rect 3608 18785 3617 18819
rect 3617 18785 3651 18819
rect 3651 18785 3660 18819
rect 3608 18776 3660 18785
rect 9036 18887 9088 18896
rect 9036 18853 9045 18887
rect 9045 18853 9079 18887
rect 9079 18853 9088 18887
rect 9036 18844 9088 18853
rect 13176 18887 13228 18896
rect 13176 18853 13185 18887
rect 13185 18853 13219 18887
rect 13219 18853 13228 18887
rect 13176 18844 13228 18853
rect 13360 18844 13412 18896
rect 6736 18819 6788 18828
rect 6736 18785 6745 18819
rect 6745 18785 6779 18819
rect 6779 18785 6788 18819
rect 6736 18776 6788 18785
rect 8668 18776 8720 18828
rect 7104 18708 7156 18760
rect 9588 18776 9640 18828
rect 10968 18819 11020 18828
rect 10968 18785 10977 18819
rect 10977 18785 11011 18819
rect 11011 18785 11020 18819
rect 10968 18776 11020 18785
rect 12164 18819 12216 18828
rect 12164 18785 12173 18819
rect 12173 18785 12207 18819
rect 12207 18785 12216 18819
rect 12164 18776 12216 18785
rect 12992 18776 13044 18828
rect 14188 18912 14240 18964
rect 13268 18708 13320 18760
rect 13360 18708 13412 18760
rect 14832 18776 14884 18828
rect 4712 18640 4764 18692
rect 8852 18640 8904 18692
rect 8944 18640 8996 18692
rect 13544 18640 13596 18692
rect 17960 18912 18012 18964
rect 18052 18912 18104 18964
rect 18880 18912 18932 18964
rect 17408 18844 17460 18896
rect 18328 18844 18380 18896
rect 21640 18912 21692 18964
rect 20812 18844 20864 18896
rect 16856 18819 16908 18828
rect 16856 18785 16865 18819
rect 16865 18785 16899 18819
rect 16899 18785 16908 18819
rect 16856 18776 16908 18785
rect 17500 18819 17552 18828
rect 17500 18785 17509 18819
rect 17509 18785 17543 18819
rect 17543 18785 17552 18819
rect 17500 18776 17552 18785
rect 17592 18819 17644 18828
rect 17592 18785 17601 18819
rect 17601 18785 17635 18819
rect 17635 18785 17644 18819
rect 17592 18776 17644 18785
rect 19248 18776 19300 18828
rect 20536 18776 20588 18828
rect 23296 18844 23348 18896
rect 20444 18751 20496 18760
rect 20444 18717 20453 18751
rect 20453 18717 20487 18751
rect 20487 18717 20496 18751
rect 20444 18708 20496 18717
rect 20720 18751 20772 18760
rect 20720 18717 20729 18751
rect 20729 18717 20763 18751
rect 20763 18717 20772 18751
rect 20720 18708 20772 18717
rect 23756 18776 23808 18828
rect 21916 18708 21968 18760
rect 20536 18640 20588 18692
rect 4896 18572 4948 18624
rect 5448 18572 5500 18624
rect 7012 18615 7064 18624
rect 7012 18581 7021 18615
rect 7021 18581 7055 18615
rect 7055 18581 7064 18615
rect 7012 18572 7064 18581
rect 8760 18572 8812 18624
rect 12624 18572 12676 18624
rect 13820 18572 13872 18624
rect 17408 18572 17460 18624
rect 19892 18615 19944 18624
rect 19892 18581 19901 18615
rect 19901 18581 19935 18615
rect 19935 18581 19944 18615
rect 19892 18572 19944 18581
rect 22192 18615 22244 18624
rect 22192 18581 22201 18615
rect 22201 18581 22235 18615
rect 22235 18581 22244 18615
rect 22192 18572 22244 18581
rect 22560 18572 22612 18624
rect 3882 18470 3934 18522
rect 3946 18470 3998 18522
rect 4010 18470 4062 18522
rect 4074 18470 4126 18522
rect 4138 18470 4190 18522
rect 10851 18470 10903 18522
rect 10915 18470 10967 18522
rect 10979 18470 11031 18522
rect 11043 18470 11095 18522
rect 11107 18470 11159 18522
rect 17820 18470 17872 18522
rect 17884 18470 17936 18522
rect 17948 18470 18000 18522
rect 18012 18470 18064 18522
rect 18076 18470 18128 18522
rect 24789 18470 24841 18522
rect 24853 18470 24905 18522
rect 24917 18470 24969 18522
rect 24981 18470 25033 18522
rect 25045 18470 25097 18522
rect 3608 18368 3660 18420
rect 1584 18207 1636 18216
rect 1584 18173 1593 18207
rect 1593 18173 1627 18207
rect 1627 18173 1636 18207
rect 1584 18164 1636 18173
rect 2136 18164 2188 18216
rect 5908 18368 5960 18420
rect 8668 18368 8720 18420
rect 4436 18275 4488 18284
rect 4436 18241 4445 18275
rect 4445 18241 4479 18275
rect 4479 18241 4488 18275
rect 4436 18232 4488 18241
rect 4620 18232 4672 18284
rect 5080 18164 5132 18216
rect 6276 18207 6328 18216
rect 6276 18173 6285 18207
rect 6285 18173 6319 18207
rect 6319 18173 6328 18207
rect 6276 18164 6328 18173
rect 6552 18164 6604 18216
rect 7012 18164 7064 18216
rect 5816 18096 5868 18148
rect 8392 18232 8444 18284
rect 9036 18368 9088 18420
rect 11520 18368 11572 18420
rect 12164 18368 12216 18420
rect 13176 18411 13228 18420
rect 13176 18377 13207 18411
rect 13207 18377 13228 18411
rect 13176 18368 13228 18377
rect 13360 18411 13412 18420
rect 13360 18377 13369 18411
rect 13369 18377 13403 18411
rect 13403 18377 13412 18411
rect 13360 18368 13412 18377
rect 13912 18368 13964 18420
rect 17592 18368 17644 18420
rect 19892 18368 19944 18420
rect 17500 18300 17552 18352
rect 8852 18207 8904 18216
rect 8852 18173 8861 18207
rect 8861 18173 8895 18207
rect 8895 18173 8904 18207
rect 8852 18164 8904 18173
rect 14004 18232 14056 18284
rect 16764 18275 16816 18284
rect 16764 18241 16773 18275
rect 16773 18241 16807 18275
rect 16807 18241 16816 18275
rect 16764 18232 16816 18241
rect 9588 18207 9640 18216
rect 9588 18173 9597 18207
rect 9597 18173 9631 18207
rect 9631 18173 9640 18207
rect 9588 18164 9640 18173
rect 9680 18207 9732 18216
rect 9680 18173 9689 18207
rect 9689 18173 9723 18207
rect 9723 18173 9732 18207
rect 9680 18164 9732 18173
rect 12440 18164 12492 18216
rect 6000 18028 6052 18080
rect 7012 18071 7064 18080
rect 7012 18037 7021 18071
rect 7021 18037 7055 18071
rect 7055 18037 7064 18071
rect 7012 18028 7064 18037
rect 8484 18028 8536 18080
rect 8944 18028 8996 18080
rect 12624 18096 12676 18148
rect 12716 18139 12768 18148
rect 12716 18105 12725 18139
rect 12725 18105 12759 18139
rect 12759 18105 12768 18139
rect 12716 18096 12768 18105
rect 12900 18096 12952 18148
rect 13728 18164 13780 18216
rect 17040 18207 17092 18216
rect 17040 18173 17049 18207
rect 17049 18173 17083 18207
rect 17083 18173 17092 18207
rect 17040 18164 17092 18173
rect 9864 18071 9916 18080
rect 9864 18037 9873 18071
rect 9873 18037 9907 18071
rect 9907 18037 9916 18071
rect 9864 18028 9916 18037
rect 16488 18139 16540 18148
rect 16488 18105 16506 18139
rect 16506 18105 16540 18139
rect 16488 18096 16540 18105
rect 18144 18164 18196 18216
rect 18328 18096 18380 18148
rect 14832 18028 14884 18080
rect 15384 18071 15436 18080
rect 15384 18037 15393 18071
rect 15393 18037 15427 18071
rect 15427 18037 15436 18071
rect 15384 18028 15436 18037
rect 19616 18071 19668 18080
rect 19616 18037 19625 18071
rect 19625 18037 19659 18071
rect 19659 18037 19668 18071
rect 19616 18028 19668 18037
rect 7366 17926 7418 17978
rect 7430 17926 7482 17978
rect 7494 17926 7546 17978
rect 7558 17926 7610 17978
rect 7622 17926 7674 17978
rect 14335 17926 14387 17978
rect 14399 17926 14451 17978
rect 14463 17926 14515 17978
rect 14527 17926 14579 17978
rect 14591 17926 14643 17978
rect 21304 17926 21356 17978
rect 21368 17926 21420 17978
rect 21432 17926 21484 17978
rect 21496 17926 21548 17978
rect 21560 17926 21612 17978
rect 28273 17926 28325 17978
rect 28337 17926 28389 17978
rect 28401 17926 28453 17978
rect 28465 17926 28517 17978
rect 28529 17926 28581 17978
rect 7012 17824 7064 17876
rect 9680 17824 9732 17876
rect 13360 17824 13412 17876
rect 13728 17824 13780 17876
rect 13268 17756 13320 17808
rect 3700 17688 3752 17740
rect 5816 17688 5868 17740
rect 6092 17688 6144 17740
rect 6552 17688 6604 17740
rect 7288 17731 7340 17740
rect 7288 17697 7297 17731
rect 7297 17697 7331 17731
rect 7331 17697 7340 17731
rect 7288 17688 7340 17697
rect 8300 17731 8352 17740
rect 8300 17697 8309 17731
rect 8309 17697 8343 17731
rect 8343 17697 8352 17731
rect 8300 17688 8352 17697
rect 8484 17688 8536 17740
rect 10048 17688 10100 17740
rect 1584 17620 1636 17672
rect 11244 17620 11296 17672
rect 8852 17552 8904 17604
rect 9588 17552 9640 17604
rect 12624 17688 12676 17740
rect 13360 17731 13412 17740
rect 13360 17697 13369 17731
rect 13369 17697 13403 17731
rect 13403 17697 13412 17731
rect 13360 17688 13412 17697
rect 13728 17731 13780 17740
rect 13728 17697 13737 17731
rect 13737 17697 13771 17731
rect 13771 17697 13780 17731
rect 13728 17688 13780 17697
rect 12440 17620 12492 17672
rect 13176 17620 13228 17672
rect 4620 17484 4672 17536
rect 6276 17527 6328 17536
rect 6276 17493 6285 17527
rect 6285 17493 6319 17527
rect 6319 17493 6328 17527
rect 6276 17484 6328 17493
rect 8760 17527 8812 17536
rect 8760 17493 8769 17527
rect 8769 17493 8803 17527
rect 8803 17493 8812 17527
rect 8760 17484 8812 17493
rect 11520 17527 11572 17536
rect 11520 17493 11529 17527
rect 11529 17493 11563 17527
rect 11563 17493 11572 17527
rect 11520 17484 11572 17493
rect 12716 17484 12768 17536
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13544 17620 13596 17629
rect 13636 17620 13688 17672
rect 14556 17663 14608 17672
rect 14556 17629 14565 17663
rect 14565 17629 14599 17663
rect 14599 17629 14608 17663
rect 14556 17620 14608 17629
rect 14648 17663 14700 17672
rect 14648 17629 14657 17663
rect 14657 17629 14691 17663
rect 14691 17629 14700 17663
rect 14648 17620 14700 17629
rect 14832 17731 14884 17740
rect 14832 17697 14841 17731
rect 14841 17697 14875 17731
rect 14875 17697 14884 17731
rect 14832 17688 14884 17697
rect 15016 17731 15068 17740
rect 15016 17697 15025 17731
rect 15025 17697 15059 17731
rect 15059 17697 15068 17731
rect 15016 17688 15068 17697
rect 15108 17688 15160 17740
rect 18696 17824 18748 17876
rect 19616 17824 19668 17876
rect 20720 17824 20772 17876
rect 16764 17688 16816 17740
rect 17684 17731 17736 17740
rect 17684 17697 17693 17731
rect 17693 17697 17727 17731
rect 17727 17697 17736 17731
rect 17684 17688 17736 17697
rect 15660 17620 15712 17672
rect 16488 17620 16540 17672
rect 17040 17620 17092 17672
rect 14004 17484 14056 17536
rect 14464 17552 14516 17604
rect 14556 17484 14608 17536
rect 14648 17484 14700 17536
rect 16948 17484 17000 17536
rect 3882 17382 3934 17434
rect 3946 17382 3998 17434
rect 4010 17382 4062 17434
rect 4074 17382 4126 17434
rect 4138 17382 4190 17434
rect 10851 17382 10903 17434
rect 10915 17382 10967 17434
rect 10979 17382 11031 17434
rect 11043 17382 11095 17434
rect 11107 17382 11159 17434
rect 17820 17382 17872 17434
rect 17884 17382 17936 17434
rect 17948 17382 18000 17434
rect 18012 17382 18064 17434
rect 18076 17382 18128 17434
rect 24789 17382 24841 17434
rect 24853 17382 24905 17434
rect 24917 17382 24969 17434
rect 24981 17382 25033 17434
rect 25045 17382 25097 17434
rect 3700 17323 3752 17332
rect 3700 17289 3709 17323
rect 3709 17289 3743 17323
rect 3743 17289 3752 17323
rect 3700 17280 3752 17289
rect 8944 17323 8996 17332
rect 8944 17289 8953 17323
rect 8953 17289 8987 17323
rect 8987 17289 8996 17323
rect 8944 17280 8996 17289
rect 9864 17323 9916 17332
rect 9864 17289 9873 17323
rect 9873 17289 9907 17323
rect 9907 17289 9916 17323
rect 9864 17280 9916 17289
rect 10048 17323 10100 17332
rect 10048 17289 10057 17323
rect 10057 17289 10091 17323
rect 10091 17289 10100 17323
rect 10048 17280 10100 17289
rect 12440 17280 12492 17332
rect 12900 17280 12952 17332
rect 13452 17280 13504 17332
rect 14004 17280 14056 17332
rect 15292 17280 15344 17332
rect 17040 17323 17092 17332
rect 17040 17289 17049 17323
rect 17049 17289 17083 17323
rect 17083 17289 17092 17323
rect 17040 17280 17092 17289
rect 13360 17144 13412 17196
rect 3332 17119 3384 17128
rect 3332 17085 3341 17119
rect 3341 17085 3375 17119
rect 3375 17085 3384 17119
rect 3332 17076 3384 17085
rect 3424 17119 3476 17128
rect 3424 17085 3433 17119
rect 3433 17085 3467 17119
rect 3467 17085 3476 17119
rect 3424 17076 3476 17085
rect 12716 17119 12768 17128
rect 12716 17085 12725 17119
rect 12725 17085 12759 17119
rect 12759 17085 12768 17119
rect 12716 17076 12768 17085
rect 6736 17008 6788 17060
rect 10416 17008 10468 17060
rect 6552 16940 6604 16992
rect 8576 16983 8628 16992
rect 8576 16949 8585 16983
rect 8585 16949 8619 16983
rect 8619 16949 8628 16983
rect 8576 16940 8628 16949
rect 8668 16983 8720 16992
rect 8668 16949 8677 16983
rect 8677 16949 8711 16983
rect 8711 16949 8720 16983
rect 8668 16940 8720 16949
rect 8944 16940 8996 16992
rect 9772 16940 9824 16992
rect 12532 16940 12584 16992
rect 13176 16983 13228 16992
rect 13176 16949 13211 16983
rect 13211 16949 13228 16983
rect 13176 16940 13228 16949
rect 13636 16940 13688 16992
rect 14004 16940 14056 16992
rect 15200 17119 15252 17128
rect 15200 17085 15209 17119
rect 15209 17085 15243 17119
rect 15243 17085 15252 17119
rect 15200 17076 15252 17085
rect 15476 17119 15528 17128
rect 15476 17085 15485 17119
rect 15485 17085 15519 17119
rect 15519 17085 15528 17119
rect 15476 17076 15528 17085
rect 16672 17144 16724 17196
rect 15936 17119 15988 17128
rect 15936 17085 15950 17119
rect 15950 17085 15984 17119
rect 15984 17085 15988 17119
rect 15936 17076 15988 17085
rect 15016 16940 15068 16992
rect 15844 17051 15896 17060
rect 15844 17017 15853 17051
rect 15853 17017 15887 17051
rect 15887 17017 15896 17051
rect 15844 17008 15896 17017
rect 16212 17051 16264 17060
rect 16212 17017 16221 17051
rect 16221 17017 16255 17051
rect 16255 17017 16264 17051
rect 16212 17008 16264 17017
rect 16396 17051 16448 17060
rect 16396 17017 16405 17051
rect 16405 17017 16439 17051
rect 16439 17017 16448 17051
rect 16396 17008 16448 17017
rect 16856 17144 16908 17196
rect 19340 17212 19392 17264
rect 23296 17212 23348 17264
rect 17408 17119 17460 17128
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 18144 17187 18196 17196
rect 18144 17153 18153 17187
rect 18153 17153 18187 17187
rect 18187 17153 18196 17187
rect 18144 17144 18196 17153
rect 18696 17144 18748 17196
rect 18972 17187 19024 17196
rect 18972 17153 18981 17187
rect 18981 17153 19015 17187
rect 19015 17153 19024 17187
rect 18972 17144 19024 17153
rect 17960 17119 18012 17128
rect 17960 17085 17969 17119
rect 17969 17085 18003 17119
rect 18003 17085 18012 17119
rect 17960 17076 18012 17085
rect 17500 16940 17552 16992
rect 18604 17076 18656 17128
rect 20352 17119 20404 17128
rect 20352 17085 20361 17119
rect 20361 17085 20395 17119
rect 20395 17085 20404 17119
rect 20352 17076 20404 17085
rect 18604 16940 18656 16992
rect 20168 16940 20220 16992
rect 7366 16838 7418 16890
rect 7430 16838 7482 16890
rect 7494 16838 7546 16890
rect 7558 16838 7610 16890
rect 7622 16838 7674 16890
rect 14335 16838 14387 16890
rect 14399 16838 14451 16890
rect 14463 16838 14515 16890
rect 14527 16838 14579 16890
rect 14591 16838 14643 16890
rect 21304 16838 21356 16890
rect 21368 16838 21420 16890
rect 21432 16838 21484 16890
rect 21496 16838 21548 16890
rect 21560 16838 21612 16890
rect 28273 16838 28325 16890
rect 28337 16838 28389 16890
rect 28401 16838 28453 16890
rect 28465 16838 28517 16890
rect 28529 16838 28581 16890
rect 3424 16736 3476 16788
rect 4804 16736 4856 16788
rect 4620 16668 4672 16720
rect 2136 16643 2188 16652
rect 2136 16609 2145 16643
rect 2145 16609 2179 16643
rect 2179 16609 2188 16643
rect 2136 16600 2188 16609
rect 4528 16643 4580 16652
rect 4528 16609 4537 16643
rect 4537 16609 4571 16643
rect 4571 16609 4580 16643
rect 4528 16600 4580 16609
rect 4712 16643 4764 16652
rect 4712 16609 4721 16643
rect 4721 16609 4755 16643
rect 4755 16609 4764 16643
rect 4712 16600 4764 16609
rect 5172 16600 5224 16652
rect 6276 16711 6328 16720
rect 6276 16677 6285 16711
rect 6285 16677 6319 16711
rect 6319 16677 6328 16711
rect 6276 16668 6328 16677
rect 6828 16736 6880 16788
rect 5356 16575 5408 16584
rect 5356 16541 5365 16575
rect 5365 16541 5399 16575
rect 5399 16541 5408 16575
rect 5356 16532 5408 16541
rect 6184 16600 6236 16652
rect 7288 16668 7340 16720
rect 6000 16532 6052 16584
rect 6552 16532 6604 16584
rect 6736 16643 6788 16652
rect 6736 16609 6745 16643
rect 6745 16609 6779 16643
rect 6779 16609 6788 16643
rect 6736 16600 6788 16609
rect 6920 16643 6972 16652
rect 6920 16609 6929 16643
rect 6929 16609 6963 16643
rect 6963 16609 6972 16643
rect 6920 16600 6972 16609
rect 7380 16643 7432 16652
rect 7380 16609 7389 16643
rect 7389 16609 7423 16643
rect 7423 16609 7432 16643
rect 7380 16600 7432 16609
rect 8300 16736 8352 16788
rect 8024 16668 8076 16720
rect 8944 16600 8996 16652
rect 9772 16779 9824 16788
rect 9772 16745 9781 16779
rect 9781 16745 9815 16779
rect 9815 16745 9824 16779
rect 9772 16736 9824 16745
rect 10324 16736 10376 16788
rect 11520 16736 11572 16788
rect 12532 16779 12584 16788
rect 12532 16745 12541 16779
rect 12541 16745 12575 16779
rect 12575 16745 12584 16779
rect 12532 16736 12584 16745
rect 13084 16736 13136 16788
rect 9680 16668 9732 16720
rect 9588 16643 9640 16652
rect 9588 16609 9597 16643
rect 9597 16609 9631 16643
rect 9631 16609 9640 16643
rect 9588 16600 9640 16609
rect 11244 16600 11296 16652
rect 14924 16668 14976 16720
rect 15016 16711 15068 16720
rect 15016 16677 15025 16711
rect 15025 16677 15059 16711
rect 15059 16677 15068 16711
rect 15016 16668 15068 16677
rect 15476 16736 15528 16788
rect 17500 16779 17552 16788
rect 17500 16745 17509 16779
rect 17509 16745 17543 16779
rect 17543 16745 17552 16779
rect 17500 16736 17552 16745
rect 17960 16736 18012 16788
rect 18696 16736 18748 16788
rect 15200 16711 15252 16720
rect 15200 16677 15241 16711
rect 15241 16677 15252 16711
rect 15200 16668 15252 16677
rect 15568 16668 15620 16720
rect 16212 16668 16264 16720
rect 16580 16668 16632 16720
rect 15844 16600 15896 16652
rect 15936 16643 15988 16652
rect 15936 16609 15945 16643
rect 15945 16609 15979 16643
rect 15979 16609 15988 16643
rect 15936 16600 15988 16609
rect 16396 16600 16448 16652
rect 6092 16507 6144 16516
rect 6092 16473 6101 16507
rect 6101 16473 6135 16507
rect 6135 16473 6144 16507
rect 6092 16464 6144 16473
rect 6368 16464 6420 16516
rect 13452 16532 13504 16584
rect 15292 16532 15344 16584
rect 7104 16464 7156 16516
rect 8668 16464 8720 16516
rect 1768 16396 1820 16448
rect 4712 16396 4764 16448
rect 10692 16396 10744 16448
rect 12992 16439 13044 16448
rect 12992 16405 13001 16439
rect 13001 16405 13035 16439
rect 13035 16405 13044 16439
rect 12992 16396 13044 16405
rect 13084 16396 13136 16448
rect 13360 16396 13412 16448
rect 16580 16464 16632 16516
rect 17224 16575 17276 16584
rect 17224 16541 17233 16575
rect 17233 16541 17267 16575
rect 17267 16541 17276 16575
rect 17224 16532 17276 16541
rect 17500 16532 17552 16584
rect 18696 16600 18748 16652
rect 19892 16600 19944 16652
rect 20168 16643 20220 16652
rect 20168 16609 20177 16643
rect 20177 16609 20211 16643
rect 20211 16609 20220 16643
rect 20168 16600 20220 16609
rect 17316 16464 17368 16516
rect 15936 16439 15988 16448
rect 15936 16405 15945 16439
rect 15945 16405 15979 16439
rect 15979 16405 15988 16439
rect 15936 16396 15988 16405
rect 17592 16396 17644 16448
rect 19432 16532 19484 16584
rect 18604 16439 18656 16448
rect 18604 16405 18613 16439
rect 18613 16405 18647 16439
rect 18647 16405 18656 16439
rect 18604 16396 18656 16405
rect 20076 16439 20128 16448
rect 20076 16405 20085 16439
rect 20085 16405 20119 16439
rect 20119 16405 20128 16439
rect 20076 16396 20128 16405
rect 3882 16294 3934 16346
rect 3946 16294 3998 16346
rect 4010 16294 4062 16346
rect 4074 16294 4126 16346
rect 4138 16294 4190 16346
rect 10851 16294 10903 16346
rect 10915 16294 10967 16346
rect 10979 16294 11031 16346
rect 11043 16294 11095 16346
rect 11107 16294 11159 16346
rect 17820 16294 17872 16346
rect 17884 16294 17936 16346
rect 17948 16294 18000 16346
rect 18012 16294 18064 16346
rect 18076 16294 18128 16346
rect 24789 16294 24841 16346
rect 24853 16294 24905 16346
rect 24917 16294 24969 16346
rect 24981 16294 25033 16346
rect 25045 16294 25097 16346
rect 4528 16192 4580 16244
rect 6736 16192 6788 16244
rect 6828 16235 6880 16244
rect 6828 16201 6837 16235
rect 6837 16201 6871 16235
rect 6871 16201 6880 16235
rect 6828 16192 6880 16201
rect 6920 16192 6972 16244
rect 7380 16192 7432 16244
rect 9588 16192 9640 16244
rect 15292 16235 15344 16244
rect 15292 16201 15301 16235
rect 15301 16201 15335 16235
rect 15335 16201 15344 16235
rect 15292 16192 15344 16201
rect 4436 16124 4488 16176
rect 3240 16056 3292 16108
rect 1584 15988 1636 16040
rect 1768 16031 1820 16040
rect 1768 15997 1802 16031
rect 1802 15997 1820 16031
rect 1768 15988 1820 15997
rect 3792 15988 3844 16040
rect 4252 15895 4304 15904
rect 4252 15861 4261 15895
rect 4261 15861 4295 15895
rect 4295 15861 4304 15895
rect 4252 15852 4304 15861
rect 4804 16031 4856 16040
rect 4804 15997 4813 16031
rect 4813 15997 4847 16031
rect 4847 15997 4856 16031
rect 4804 15988 4856 15997
rect 5356 15988 5408 16040
rect 6368 15988 6420 16040
rect 8668 16124 8720 16176
rect 4620 15963 4672 15972
rect 4620 15929 4629 15963
rect 4629 15929 4663 15963
rect 4663 15929 4672 15963
rect 4620 15920 4672 15929
rect 5724 15920 5776 15972
rect 6092 15920 6144 15972
rect 6552 15920 6604 15972
rect 7104 15920 7156 15972
rect 8576 15988 8628 16040
rect 8760 15920 8812 15972
rect 8944 16031 8996 16040
rect 8944 15997 8953 16031
rect 8953 15997 8987 16031
rect 8987 15997 8996 16031
rect 8944 15988 8996 15997
rect 11888 16056 11940 16108
rect 14832 16056 14884 16108
rect 10692 15988 10744 16040
rect 11244 16031 11296 16040
rect 11244 15997 11253 16031
rect 11253 15997 11287 16031
rect 11287 15997 11296 16031
rect 11244 15988 11296 15997
rect 11612 16031 11664 16040
rect 11612 15997 11621 16031
rect 11621 15997 11655 16031
rect 11655 15997 11664 16031
rect 11612 15988 11664 15997
rect 12992 15988 13044 16040
rect 13176 16031 13228 16040
rect 13176 15997 13185 16031
rect 13185 15997 13219 16031
rect 13219 15997 13228 16031
rect 13176 15988 13228 15997
rect 13268 15988 13320 16040
rect 14004 16031 14056 16040
rect 14004 15997 14013 16031
rect 14013 15997 14047 16031
rect 14047 15997 14056 16031
rect 14004 15988 14056 15997
rect 13544 15920 13596 15972
rect 15568 15988 15620 16040
rect 15752 16167 15804 16176
rect 15752 16133 15761 16167
rect 15761 16133 15795 16167
rect 15795 16133 15804 16167
rect 15752 16124 15804 16133
rect 17408 16192 17460 16244
rect 17960 16235 18012 16244
rect 17960 16201 17969 16235
rect 17969 16201 18003 16235
rect 18003 16201 18012 16235
rect 17960 16192 18012 16201
rect 18788 16192 18840 16244
rect 20536 16167 20588 16176
rect 20536 16133 20545 16167
rect 20545 16133 20579 16167
rect 20579 16133 20588 16167
rect 20536 16124 20588 16133
rect 16580 15988 16632 16040
rect 17040 16031 17092 16040
rect 17040 15997 17049 16031
rect 17049 15997 17083 16031
rect 17083 15997 17092 16031
rect 17040 15988 17092 15997
rect 17132 16031 17184 16040
rect 17132 15997 17141 16031
rect 17141 15997 17175 16031
rect 17175 15997 17184 16031
rect 17132 15988 17184 15997
rect 4712 15852 4764 15904
rect 7288 15852 7340 15904
rect 9864 15895 9916 15904
rect 9864 15861 9873 15895
rect 9873 15861 9907 15895
rect 9907 15861 9916 15895
rect 9864 15852 9916 15861
rect 11428 15895 11480 15904
rect 11428 15861 11437 15895
rect 11437 15861 11471 15895
rect 11471 15861 11480 15895
rect 11428 15852 11480 15861
rect 12808 15852 12860 15904
rect 13084 15852 13136 15904
rect 13636 15895 13688 15904
rect 13636 15861 13645 15895
rect 13645 15861 13679 15895
rect 13679 15861 13688 15895
rect 13636 15852 13688 15861
rect 15016 15852 15068 15904
rect 17500 15988 17552 16040
rect 17592 15852 17644 15904
rect 22100 16056 22152 16108
rect 22928 16056 22980 16108
rect 17868 16031 17920 16040
rect 17868 15997 17877 16031
rect 17877 15997 17911 16031
rect 17911 15997 17920 16031
rect 17868 15988 17920 15997
rect 18512 15988 18564 16040
rect 20168 15920 20220 15972
rect 17776 15852 17828 15904
rect 7366 15750 7418 15802
rect 7430 15750 7482 15802
rect 7494 15750 7546 15802
rect 7558 15750 7610 15802
rect 7622 15750 7674 15802
rect 14335 15750 14387 15802
rect 14399 15750 14451 15802
rect 14463 15750 14515 15802
rect 14527 15750 14579 15802
rect 14591 15750 14643 15802
rect 21304 15750 21356 15802
rect 21368 15750 21420 15802
rect 21432 15750 21484 15802
rect 21496 15750 21548 15802
rect 21560 15750 21612 15802
rect 28273 15750 28325 15802
rect 28337 15750 28389 15802
rect 28401 15750 28453 15802
rect 28465 15750 28517 15802
rect 28529 15750 28581 15802
rect 2136 15691 2188 15700
rect 2136 15657 2145 15691
rect 2145 15657 2179 15691
rect 2179 15657 2188 15691
rect 2136 15648 2188 15657
rect 4252 15648 4304 15700
rect 6460 15648 6512 15700
rect 13176 15648 13228 15700
rect 13636 15648 13688 15700
rect 17316 15648 17368 15700
rect 17960 15648 18012 15700
rect 20076 15648 20128 15700
rect 20168 15691 20220 15700
rect 20168 15657 20177 15691
rect 20177 15657 20211 15691
rect 20211 15657 20220 15691
rect 20168 15648 20220 15657
rect 20536 15648 20588 15700
rect 4528 15512 4580 15564
rect 5448 15512 5500 15564
rect 6092 15555 6144 15564
rect 6092 15521 6125 15555
rect 6125 15521 6144 15555
rect 6092 15512 6144 15521
rect 2412 15444 2464 15496
rect 5172 15487 5224 15496
rect 5172 15453 5181 15487
rect 5181 15453 5215 15487
rect 5215 15453 5224 15487
rect 6368 15512 6420 15564
rect 7472 15512 7524 15564
rect 13452 15555 13504 15564
rect 13452 15521 13461 15555
rect 13461 15521 13495 15555
rect 13495 15521 13504 15555
rect 13452 15512 13504 15521
rect 5172 15444 5224 15453
rect 8576 15487 8628 15496
rect 8576 15453 8585 15487
rect 8585 15453 8619 15487
rect 8619 15453 8628 15487
rect 8576 15444 8628 15453
rect 8668 15444 8720 15496
rect 14188 15444 14240 15496
rect 3792 15376 3844 15428
rect 9680 15376 9732 15428
rect 10692 15376 10744 15428
rect 17040 15555 17092 15564
rect 17040 15521 17050 15555
rect 17050 15521 17084 15555
rect 17084 15521 17092 15555
rect 17040 15512 17092 15521
rect 17224 15555 17276 15564
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 18144 15444 18196 15496
rect 18696 15487 18748 15496
rect 18696 15453 18705 15487
rect 18705 15453 18739 15487
rect 18739 15453 18748 15487
rect 18696 15444 18748 15453
rect 19064 15555 19116 15564
rect 19064 15521 19073 15555
rect 19073 15521 19107 15555
rect 19107 15521 19116 15555
rect 19064 15512 19116 15521
rect 19340 15512 19392 15564
rect 19892 15555 19944 15564
rect 19892 15521 19901 15555
rect 19901 15521 19935 15555
rect 19935 15521 19944 15555
rect 19892 15512 19944 15521
rect 19984 15512 20036 15564
rect 20628 15555 20680 15564
rect 20628 15521 20637 15555
rect 20637 15521 20671 15555
rect 20671 15521 20680 15555
rect 20628 15512 20680 15521
rect 20996 15580 21048 15632
rect 22468 15580 22520 15632
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 22928 15512 22980 15564
rect 3332 15308 3384 15360
rect 5816 15308 5868 15360
rect 11980 15308 12032 15360
rect 17316 15308 17368 15360
rect 19064 15308 19116 15360
rect 20260 15308 20312 15360
rect 20352 15351 20404 15360
rect 20352 15317 20361 15351
rect 20361 15317 20395 15351
rect 20395 15317 20404 15351
rect 20352 15308 20404 15317
rect 21640 15351 21692 15360
rect 21640 15317 21649 15351
rect 21649 15317 21683 15351
rect 21683 15317 21692 15351
rect 21640 15308 21692 15317
rect 3882 15206 3934 15258
rect 3946 15206 3998 15258
rect 4010 15206 4062 15258
rect 4074 15206 4126 15258
rect 4138 15206 4190 15258
rect 10851 15206 10903 15258
rect 10915 15206 10967 15258
rect 10979 15206 11031 15258
rect 11043 15206 11095 15258
rect 11107 15206 11159 15258
rect 17820 15206 17872 15258
rect 17884 15206 17936 15258
rect 17948 15206 18000 15258
rect 18012 15206 18064 15258
rect 18076 15206 18128 15258
rect 24789 15206 24841 15258
rect 24853 15206 24905 15258
rect 24917 15206 24969 15258
rect 24981 15206 25033 15258
rect 25045 15206 25097 15258
rect 4436 15104 4488 15156
rect 7472 15147 7524 15156
rect 7472 15113 7481 15147
rect 7481 15113 7515 15147
rect 7515 15113 7524 15147
rect 7472 15104 7524 15113
rect 8576 15104 8628 15156
rect 3148 15036 3200 15088
rect 3056 14900 3108 14952
rect 3700 14943 3752 14952
rect 3700 14909 3709 14943
rect 3709 14909 3743 14943
rect 3743 14909 3752 14943
rect 3700 14900 3752 14909
rect 3884 14943 3936 14952
rect 3884 14909 3893 14943
rect 3893 14909 3927 14943
rect 3927 14909 3936 14943
rect 3884 14900 3936 14909
rect 4528 14900 4580 14952
rect 5172 14900 5224 14952
rect 5908 14943 5960 14952
rect 5908 14909 5917 14943
rect 5917 14909 5951 14943
rect 5951 14909 5960 14943
rect 5908 14900 5960 14909
rect 8944 14968 8996 15020
rect 9772 15011 9824 15020
rect 9772 14977 9781 15011
rect 9781 14977 9815 15011
rect 9815 14977 9824 15011
rect 9772 14968 9824 14977
rect 6276 14832 6328 14884
rect 6368 14832 6420 14884
rect 9588 14900 9640 14952
rect 9956 14900 10008 14952
rect 10692 15036 10744 15088
rect 11336 14968 11388 15020
rect 12072 15147 12124 15156
rect 12072 15113 12081 15147
rect 12081 15113 12115 15147
rect 12115 15113 12124 15147
rect 12072 15104 12124 15113
rect 19984 15147 20036 15156
rect 19984 15113 19993 15147
rect 19993 15113 20027 15147
rect 20027 15113 20036 15147
rect 19984 15104 20036 15113
rect 21272 15104 21324 15156
rect 13912 15036 13964 15088
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 3424 14764 3476 14816
rect 6092 14764 6144 14816
rect 7748 14764 7800 14816
rect 8760 14764 8812 14816
rect 8944 14764 8996 14816
rect 9680 14764 9732 14816
rect 10324 14807 10376 14816
rect 10324 14773 10333 14807
rect 10333 14773 10367 14807
rect 10367 14773 10376 14807
rect 10324 14764 10376 14773
rect 10600 14807 10652 14816
rect 10600 14773 10609 14807
rect 10609 14773 10643 14807
rect 10643 14773 10652 14807
rect 10600 14764 10652 14773
rect 10692 14764 10744 14816
rect 11520 14764 11572 14816
rect 11704 14943 11756 14952
rect 11704 14909 11713 14943
rect 11713 14909 11747 14943
rect 11747 14909 11756 14943
rect 11704 14900 11756 14909
rect 11980 14900 12032 14952
rect 12348 14943 12400 14952
rect 12348 14909 12357 14943
rect 12357 14909 12391 14943
rect 12391 14909 12400 14943
rect 12348 14900 12400 14909
rect 13820 14875 13872 14884
rect 13820 14841 13829 14875
rect 13829 14841 13863 14875
rect 13863 14841 13872 14875
rect 13820 14832 13872 14841
rect 14096 14900 14148 14952
rect 14832 14900 14884 14952
rect 15016 14900 15068 14952
rect 15660 14943 15712 14952
rect 15660 14909 15669 14943
rect 15669 14909 15703 14943
rect 15703 14909 15712 14943
rect 15660 14900 15712 14909
rect 17224 15036 17276 15088
rect 18788 15036 18840 15088
rect 18328 14968 18380 15020
rect 16120 14832 16172 14884
rect 17040 14832 17092 14884
rect 20260 15036 20312 15088
rect 20628 14968 20680 15020
rect 20444 14943 20496 14952
rect 20444 14909 20453 14943
rect 20453 14909 20487 14943
rect 20487 14909 20496 14943
rect 20444 14900 20496 14909
rect 20996 14943 21048 14952
rect 20996 14909 21005 14943
rect 21005 14909 21039 14943
rect 21039 14909 21048 14943
rect 20996 14900 21048 14909
rect 20628 14832 20680 14884
rect 11704 14764 11756 14816
rect 13912 14807 13964 14816
rect 13912 14773 13921 14807
rect 13921 14773 13955 14807
rect 13955 14773 13964 14807
rect 13912 14764 13964 14773
rect 14004 14764 14056 14816
rect 14188 14764 14240 14816
rect 18328 14807 18380 14816
rect 18328 14773 18337 14807
rect 18337 14773 18371 14807
rect 18371 14773 18380 14807
rect 18328 14764 18380 14773
rect 21916 14943 21968 14952
rect 21916 14909 21925 14943
rect 21925 14909 21959 14943
rect 21959 14909 21968 14943
rect 21916 14900 21968 14909
rect 22192 14900 22244 14952
rect 21640 14832 21692 14884
rect 7366 14662 7418 14714
rect 7430 14662 7482 14714
rect 7494 14662 7546 14714
rect 7558 14662 7610 14714
rect 7622 14662 7674 14714
rect 14335 14662 14387 14714
rect 14399 14662 14451 14714
rect 14463 14662 14515 14714
rect 14527 14662 14579 14714
rect 14591 14662 14643 14714
rect 21304 14662 21356 14714
rect 21368 14662 21420 14714
rect 21432 14662 21484 14714
rect 21496 14662 21548 14714
rect 21560 14662 21612 14714
rect 28273 14662 28325 14714
rect 28337 14662 28389 14714
rect 28401 14662 28453 14714
rect 28465 14662 28517 14714
rect 28529 14662 28581 14714
rect 3148 14560 3200 14612
rect 3424 14560 3476 14612
rect 6276 14603 6328 14612
rect 6276 14569 6285 14603
rect 6285 14569 6319 14603
rect 6319 14569 6328 14603
rect 6276 14560 6328 14569
rect 9864 14560 9916 14612
rect 10600 14560 10652 14612
rect 11336 14560 11388 14612
rect 12348 14560 12400 14612
rect 13820 14560 13872 14612
rect 14004 14560 14056 14612
rect 15568 14603 15620 14612
rect 15568 14569 15577 14603
rect 15577 14569 15611 14603
rect 15611 14569 15620 14603
rect 15568 14560 15620 14569
rect 16120 14603 16172 14612
rect 16120 14569 16129 14603
rect 16129 14569 16163 14603
rect 16163 14569 16172 14603
rect 16120 14560 16172 14569
rect 17316 14603 17368 14612
rect 17316 14569 17325 14603
rect 17325 14569 17359 14603
rect 17359 14569 17368 14603
rect 17316 14560 17368 14569
rect 5448 14492 5500 14544
rect 3240 14356 3292 14408
rect 3792 14467 3844 14476
rect 3792 14433 3801 14467
rect 3801 14433 3835 14467
rect 3835 14433 3844 14467
rect 3792 14424 3844 14433
rect 6000 14467 6052 14476
rect 6000 14433 6009 14467
rect 6009 14433 6043 14467
rect 6043 14433 6052 14467
rect 6000 14424 6052 14433
rect 7748 14424 7800 14476
rect 8668 14467 8720 14476
rect 8668 14433 8677 14467
rect 8677 14433 8711 14467
rect 8711 14433 8720 14467
rect 8668 14424 8720 14433
rect 10692 14492 10744 14544
rect 11704 14492 11756 14544
rect 12808 14535 12860 14544
rect 12808 14501 12842 14535
rect 12842 14501 12860 14535
rect 12808 14492 12860 14501
rect 11336 14467 11388 14476
rect 11336 14433 11370 14467
rect 11370 14433 11388 14467
rect 11336 14424 11388 14433
rect 14096 14424 14148 14476
rect 14740 14467 14792 14476
rect 14740 14433 14749 14467
rect 14749 14433 14783 14467
rect 14783 14433 14792 14467
rect 14740 14424 14792 14433
rect 4620 14356 4672 14408
rect 5816 14399 5868 14408
rect 5816 14365 5825 14399
rect 5825 14365 5859 14399
rect 5859 14365 5868 14399
rect 5816 14356 5868 14365
rect 8116 14356 8168 14408
rect 8944 14399 8996 14408
rect 8944 14365 8953 14399
rect 8953 14365 8987 14399
rect 8987 14365 8996 14399
rect 8944 14356 8996 14365
rect 9956 14356 10008 14408
rect 9680 14288 9732 14340
rect 10140 14288 10192 14340
rect 10508 14220 10560 14272
rect 10692 14220 10744 14272
rect 11244 14220 11296 14272
rect 14004 14399 14056 14408
rect 14004 14365 14013 14399
rect 14013 14365 14047 14399
rect 14047 14365 14056 14399
rect 14004 14356 14056 14365
rect 16948 14467 17000 14476
rect 16948 14433 16957 14467
rect 16957 14433 16991 14467
rect 16991 14433 17000 14467
rect 16948 14424 17000 14433
rect 18972 14492 19024 14544
rect 19064 14424 19116 14476
rect 21640 14424 21692 14476
rect 14924 14288 14976 14340
rect 18788 14288 18840 14340
rect 15016 14220 15068 14272
rect 15844 14220 15896 14272
rect 19340 14263 19392 14272
rect 19340 14229 19349 14263
rect 19349 14229 19383 14263
rect 19383 14229 19392 14263
rect 19340 14220 19392 14229
rect 22284 14220 22336 14272
rect 3882 14118 3934 14170
rect 3946 14118 3998 14170
rect 4010 14118 4062 14170
rect 4074 14118 4126 14170
rect 4138 14118 4190 14170
rect 10851 14118 10903 14170
rect 10915 14118 10967 14170
rect 10979 14118 11031 14170
rect 11043 14118 11095 14170
rect 11107 14118 11159 14170
rect 17820 14118 17872 14170
rect 17884 14118 17936 14170
rect 17948 14118 18000 14170
rect 18012 14118 18064 14170
rect 18076 14118 18128 14170
rect 24789 14118 24841 14170
rect 24853 14118 24905 14170
rect 24917 14118 24969 14170
rect 24981 14118 25033 14170
rect 25045 14118 25097 14170
rect 6000 14059 6052 14068
rect 6000 14025 6009 14059
rect 6009 14025 6043 14059
rect 6043 14025 6052 14059
rect 6000 14016 6052 14025
rect 7748 14016 7800 14068
rect 8944 14059 8996 14068
rect 8944 14025 8953 14059
rect 8953 14025 8987 14059
rect 8987 14025 8996 14059
rect 8944 14016 8996 14025
rect 11336 14016 11388 14068
rect 19340 14016 19392 14068
rect 2044 13855 2096 13864
rect 2044 13821 2053 13855
rect 2053 13821 2087 13855
rect 2087 13821 2096 13855
rect 2044 13812 2096 13821
rect 3240 13744 3292 13796
rect 4068 13812 4120 13864
rect 4528 13812 4580 13864
rect 4804 13812 4856 13864
rect 5724 13855 5776 13864
rect 5724 13821 5733 13855
rect 5733 13821 5767 13855
rect 5767 13821 5776 13855
rect 5724 13812 5776 13821
rect 10508 13948 10560 14000
rect 5080 13744 5132 13796
rect 5632 13787 5684 13796
rect 5632 13753 5641 13787
rect 5641 13753 5675 13787
rect 5675 13753 5684 13787
rect 5632 13744 5684 13753
rect 1768 13676 1820 13728
rect 4160 13719 4212 13728
rect 4160 13685 4169 13719
rect 4169 13685 4203 13719
rect 4203 13685 4212 13719
rect 4160 13676 4212 13685
rect 4528 13676 4580 13728
rect 4712 13676 4764 13728
rect 7196 13744 7248 13796
rect 11428 13880 11480 13932
rect 17224 13880 17276 13932
rect 18972 13880 19024 13932
rect 9864 13812 9916 13864
rect 10692 13812 10744 13864
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 18328 13812 18380 13864
rect 19064 13855 19116 13864
rect 19064 13821 19073 13855
rect 19073 13821 19107 13855
rect 19107 13821 19116 13855
rect 19064 13812 19116 13821
rect 19432 13812 19484 13864
rect 19524 13855 19576 13864
rect 19524 13821 19533 13855
rect 19533 13821 19567 13855
rect 19567 13821 19576 13855
rect 19524 13812 19576 13821
rect 19892 13855 19944 13864
rect 19892 13821 19901 13855
rect 19901 13821 19935 13855
rect 19935 13821 19944 13855
rect 19892 13812 19944 13821
rect 20352 13812 20404 13864
rect 20628 13812 20680 13864
rect 7288 13719 7340 13728
rect 7288 13685 7297 13719
rect 7297 13685 7331 13719
rect 7331 13685 7340 13719
rect 7288 13676 7340 13685
rect 7748 13676 7800 13728
rect 13452 13676 13504 13728
rect 13728 13719 13780 13728
rect 13728 13685 13737 13719
rect 13737 13685 13771 13719
rect 13771 13685 13780 13719
rect 13728 13676 13780 13685
rect 18880 13676 18932 13728
rect 19432 13719 19484 13728
rect 19432 13685 19441 13719
rect 19441 13685 19475 13719
rect 19475 13685 19484 13719
rect 19432 13676 19484 13685
rect 19984 13676 20036 13728
rect 20260 13676 20312 13728
rect 22008 13744 22060 13796
rect 22284 13787 22336 13796
rect 22284 13753 22302 13787
rect 22302 13753 22336 13787
rect 22284 13744 22336 13753
rect 21088 13719 21140 13728
rect 21088 13685 21097 13719
rect 21097 13685 21131 13719
rect 21131 13685 21140 13719
rect 21088 13676 21140 13685
rect 7366 13574 7418 13626
rect 7430 13574 7482 13626
rect 7494 13574 7546 13626
rect 7558 13574 7610 13626
rect 7622 13574 7674 13626
rect 14335 13574 14387 13626
rect 14399 13574 14451 13626
rect 14463 13574 14515 13626
rect 14527 13574 14579 13626
rect 14591 13574 14643 13626
rect 21304 13574 21356 13626
rect 21368 13574 21420 13626
rect 21432 13574 21484 13626
rect 21496 13574 21548 13626
rect 21560 13574 21612 13626
rect 28273 13574 28325 13626
rect 28337 13574 28389 13626
rect 28401 13574 28453 13626
rect 28465 13574 28517 13626
rect 28529 13574 28581 13626
rect 1584 13404 1636 13456
rect 5908 13472 5960 13524
rect 3056 13404 3108 13456
rect 1768 13379 1820 13388
rect 1768 13345 1802 13379
rect 1802 13345 1820 13379
rect 1768 13336 1820 13345
rect 4068 13404 4120 13456
rect 4160 13404 4212 13456
rect 5080 13404 5132 13456
rect 3240 13311 3292 13320
rect 3240 13277 3249 13311
rect 3249 13277 3283 13311
rect 3283 13277 3292 13311
rect 3240 13268 3292 13277
rect 4528 13379 4580 13388
rect 4528 13345 4537 13379
rect 4537 13345 4571 13379
rect 4571 13345 4580 13379
rect 4528 13336 4580 13345
rect 4712 13379 4764 13388
rect 4712 13345 4721 13379
rect 4721 13345 4755 13379
rect 4755 13345 4764 13379
rect 4712 13336 4764 13345
rect 4896 13379 4948 13388
rect 4896 13345 4905 13379
rect 4905 13345 4939 13379
rect 4939 13345 4948 13379
rect 7748 13472 7800 13524
rect 10324 13472 10376 13524
rect 10416 13472 10468 13524
rect 8208 13404 8260 13456
rect 11244 13404 11296 13456
rect 11428 13447 11480 13456
rect 11428 13413 11437 13447
rect 11437 13413 11471 13447
rect 11471 13413 11480 13447
rect 11428 13404 11480 13413
rect 14188 13472 14240 13524
rect 13636 13404 13688 13456
rect 13820 13404 13872 13456
rect 14740 13404 14792 13456
rect 4896 13336 4948 13345
rect 9864 13379 9916 13388
rect 9864 13345 9873 13379
rect 9873 13345 9907 13379
rect 9907 13345 9916 13379
rect 9864 13336 9916 13345
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 4620 13268 4672 13320
rect 9036 13268 9088 13320
rect 9404 13268 9456 13320
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 3516 13243 3568 13252
rect 3516 13209 3525 13243
rect 3525 13209 3559 13243
rect 3559 13209 3568 13243
rect 3516 13200 3568 13209
rect 3792 13200 3844 13252
rect 14004 13268 14056 13320
rect 13912 13200 13964 13252
rect 14188 13336 14240 13388
rect 14372 13379 14424 13388
rect 14372 13345 14381 13379
rect 14381 13345 14415 13379
rect 14415 13345 14424 13379
rect 14372 13336 14424 13345
rect 16304 13472 16356 13524
rect 15200 13379 15252 13388
rect 3424 13132 3476 13184
rect 9680 13175 9732 13184
rect 9680 13141 9689 13175
rect 9689 13141 9723 13175
rect 9723 13141 9732 13175
rect 9680 13132 9732 13141
rect 10416 13175 10468 13184
rect 10416 13141 10425 13175
rect 10425 13141 10459 13175
rect 10459 13141 10468 13175
rect 10416 13132 10468 13141
rect 11704 13175 11756 13184
rect 11704 13141 11713 13175
rect 11713 13141 11747 13175
rect 11747 13141 11756 13175
rect 11704 13132 11756 13141
rect 12900 13132 12952 13184
rect 12992 13132 13044 13184
rect 13544 13175 13596 13184
rect 13544 13141 13553 13175
rect 13553 13141 13587 13175
rect 13587 13141 13596 13175
rect 13544 13132 13596 13141
rect 15200 13345 15209 13379
rect 15209 13345 15243 13379
rect 15243 13345 15252 13379
rect 15200 13336 15252 13345
rect 15568 13404 15620 13456
rect 15844 13379 15896 13388
rect 15844 13345 15853 13379
rect 15853 13345 15887 13379
rect 15887 13345 15896 13379
rect 15844 13336 15896 13345
rect 16212 13336 16264 13388
rect 16304 13379 16356 13388
rect 16304 13345 16313 13379
rect 16313 13345 16347 13379
rect 16347 13345 16356 13379
rect 16304 13336 16356 13345
rect 17684 13404 17736 13456
rect 19340 13472 19392 13524
rect 19524 13515 19576 13524
rect 19524 13481 19533 13515
rect 19533 13481 19567 13515
rect 19567 13481 19576 13515
rect 19524 13472 19576 13481
rect 19892 13472 19944 13524
rect 21088 13472 21140 13524
rect 21640 13515 21692 13524
rect 21640 13481 21649 13515
rect 21649 13481 21683 13515
rect 21683 13481 21692 13515
rect 21640 13472 21692 13481
rect 18788 13404 18840 13456
rect 19432 13336 19484 13388
rect 14556 13200 14608 13252
rect 14832 13132 14884 13184
rect 15016 13132 15068 13184
rect 15568 13175 15620 13184
rect 15568 13141 15577 13175
rect 15577 13141 15611 13175
rect 15611 13141 15620 13175
rect 15568 13132 15620 13141
rect 16120 13175 16172 13184
rect 16120 13141 16129 13175
rect 16129 13141 16163 13175
rect 16163 13141 16172 13175
rect 16120 13132 16172 13141
rect 18052 13311 18104 13320
rect 18052 13277 18061 13311
rect 18061 13277 18095 13311
rect 18095 13277 18104 13311
rect 18052 13268 18104 13277
rect 18604 13311 18656 13320
rect 18604 13277 18613 13311
rect 18613 13277 18647 13311
rect 18647 13277 18656 13311
rect 18604 13268 18656 13277
rect 16764 13200 16816 13252
rect 17040 13132 17092 13184
rect 18880 13311 18932 13320
rect 18880 13277 18889 13311
rect 18889 13277 18923 13311
rect 18923 13277 18932 13311
rect 18880 13268 18932 13277
rect 18972 13200 19024 13252
rect 20352 13268 20404 13320
rect 21916 13268 21968 13320
rect 19616 13175 19668 13184
rect 19616 13141 19625 13175
rect 19625 13141 19659 13175
rect 19659 13141 19668 13175
rect 19616 13132 19668 13141
rect 3882 13030 3934 13082
rect 3946 13030 3998 13082
rect 4010 13030 4062 13082
rect 4074 13030 4126 13082
rect 4138 13030 4190 13082
rect 10851 13030 10903 13082
rect 10915 13030 10967 13082
rect 10979 13030 11031 13082
rect 11043 13030 11095 13082
rect 11107 13030 11159 13082
rect 17820 13030 17872 13082
rect 17884 13030 17936 13082
rect 17948 13030 18000 13082
rect 18012 13030 18064 13082
rect 18076 13030 18128 13082
rect 24789 13030 24841 13082
rect 24853 13030 24905 13082
rect 24917 13030 24969 13082
rect 24981 13030 25033 13082
rect 25045 13030 25097 13082
rect 2044 12971 2096 12980
rect 2044 12937 2053 12971
rect 2053 12937 2087 12971
rect 2087 12937 2096 12971
rect 2044 12928 2096 12937
rect 3424 12928 3476 12980
rect 3516 12928 3568 12980
rect 4712 12928 4764 12980
rect 5632 12928 5684 12980
rect 7748 12928 7800 12980
rect 9036 12971 9088 12980
rect 9036 12937 9045 12971
rect 9045 12937 9079 12971
rect 9079 12937 9088 12971
rect 9036 12928 9088 12937
rect 9772 12928 9824 12980
rect 10508 12928 10560 12980
rect 10416 12860 10468 12912
rect 11888 12928 11940 12980
rect 2412 12767 2464 12776
rect 2412 12733 2421 12767
rect 2421 12733 2455 12767
rect 2455 12733 2464 12767
rect 2412 12724 2464 12733
rect 3792 12767 3844 12776
rect 3792 12733 3801 12767
rect 3801 12733 3835 12767
rect 3835 12733 3844 12767
rect 3792 12724 3844 12733
rect 6092 12724 6144 12776
rect 7196 12792 7248 12844
rect 7288 12724 7340 12776
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 8668 12767 8720 12776
rect 8668 12733 8677 12767
rect 8677 12733 8711 12767
rect 8711 12733 8720 12767
rect 8668 12724 8720 12733
rect 8944 12724 8996 12776
rect 9772 12767 9824 12776
rect 9772 12733 9781 12767
rect 9781 12733 9815 12767
rect 9815 12733 9824 12767
rect 9772 12724 9824 12733
rect 10140 12792 10192 12844
rect 10784 12792 10836 12844
rect 11244 12835 11296 12844
rect 11244 12801 11253 12835
rect 11253 12801 11287 12835
rect 11287 12801 11296 12835
rect 11244 12792 11296 12801
rect 10232 12724 10284 12776
rect 7104 12631 7156 12640
rect 7104 12597 7113 12631
rect 7113 12597 7147 12631
rect 7147 12597 7156 12631
rect 7104 12588 7156 12597
rect 9864 12699 9916 12708
rect 9864 12665 9873 12699
rect 9873 12665 9907 12699
rect 9907 12665 9916 12699
rect 9864 12656 9916 12665
rect 10324 12656 10376 12708
rect 11888 12656 11940 12708
rect 12992 12971 13044 12980
rect 12992 12937 13001 12971
rect 13001 12937 13035 12971
rect 13035 12937 13044 12971
rect 12992 12928 13044 12937
rect 13544 12928 13596 12980
rect 14740 12860 14792 12912
rect 12900 12792 12952 12844
rect 15200 12792 15252 12844
rect 16120 12835 16172 12844
rect 16120 12801 16129 12835
rect 16129 12801 16163 12835
rect 16163 12801 16172 12835
rect 16120 12792 16172 12801
rect 13452 12656 13504 12708
rect 13728 12699 13780 12708
rect 13728 12665 13755 12699
rect 13755 12665 13780 12699
rect 13728 12656 13780 12665
rect 14372 12724 14424 12776
rect 15016 12767 15068 12776
rect 15016 12733 15025 12767
rect 15025 12733 15059 12767
rect 15059 12733 15068 12767
rect 15016 12724 15068 12733
rect 15292 12767 15344 12776
rect 15292 12733 15301 12767
rect 15301 12733 15335 12767
rect 15335 12733 15344 12767
rect 15292 12724 15344 12733
rect 14004 12656 14056 12708
rect 14832 12699 14884 12708
rect 14832 12665 14841 12699
rect 14841 12665 14875 12699
rect 14875 12665 14884 12699
rect 16304 12724 16356 12776
rect 17040 12767 17092 12776
rect 17040 12733 17049 12767
rect 17049 12733 17083 12767
rect 17083 12733 17092 12767
rect 17040 12724 17092 12733
rect 17684 12928 17736 12980
rect 17224 12792 17276 12844
rect 17592 12860 17644 12912
rect 19984 12860 20036 12912
rect 14832 12656 14884 12665
rect 10232 12588 10284 12640
rect 10600 12631 10652 12640
rect 10600 12597 10609 12631
rect 10609 12597 10643 12631
rect 10643 12597 10652 12631
rect 10600 12588 10652 12597
rect 10784 12631 10836 12640
rect 10784 12597 10811 12631
rect 10811 12597 10836 12631
rect 10784 12588 10836 12597
rect 12808 12631 12860 12640
rect 12808 12597 12817 12631
rect 12817 12597 12851 12631
rect 12851 12597 12860 12631
rect 12808 12588 12860 12597
rect 13084 12588 13136 12640
rect 13544 12631 13596 12640
rect 13544 12597 13553 12631
rect 13553 12597 13587 12631
rect 13587 12597 13596 12631
rect 13544 12588 13596 12597
rect 15108 12588 15160 12640
rect 15200 12631 15252 12640
rect 15200 12597 15209 12631
rect 15209 12597 15243 12631
rect 15243 12597 15252 12631
rect 15200 12588 15252 12597
rect 19708 12656 19760 12708
rect 20628 12656 20680 12708
rect 16764 12588 16816 12640
rect 17224 12588 17276 12640
rect 20352 12588 20404 12640
rect 7366 12486 7418 12538
rect 7430 12486 7482 12538
rect 7494 12486 7546 12538
rect 7558 12486 7610 12538
rect 7622 12486 7674 12538
rect 14335 12486 14387 12538
rect 14399 12486 14451 12538
rect 14463 12486 14515 12538
rect 14527 12486 14579 12538
rect 14591 12486 14643 12538
rect 21304 12486 21356 12538
rect 21368 12486 21420 12538
rect 21432 12486 21484 12538
rect 21496 12486 21548 12538
rect 21560 12486 21612 12538
rect 28273 12486 28325 12538
rect 28337 12486 28389 12538
rect 28401 12486 28453 12538
rect 28465 12486 28517 12538
rect 28529 12486 28581 12538
rect 4620 12384 4672 12436
rect 4344 12316 4396 12368
rect 5448 12291 5500 12300
rect 5448 12257 5457 12291
rect 5457 12257 5491 12291
rect 5491 12257 5500 12291
rect 5448 12248 5500 12257
rect 5724 12248 5776 12300
rect 6184 12291 6236 12300
rect 6184 12257 6193 12291
rect 6193 12257 6227 12291
rect 6227 12257 6236 12291
rect 6184 12248 6236 12257
rect 7104 12316 7156 12368
rect 7656 12359 7708 12368
rect 7656 12325 7665 12359
rect 7665 12325 7699 12359
rect 7699 12325 7708 12359
rect 7656 12316 7708 12325
rect 7196 12223 7248 12232
rect 7196 12189 7205 12223
rect 7205 12189 7239 12223
rect 7239 12189 7248 12223
rect 7196 12180 7248 12189
rect 8668 12316 8720 12368
rect 9772 12384 9824 12436
rect 11980 12384 12032 12436
rect 12164 12384 12216 12436
rect 13084 12384 13136 12436
rect 5816 12087 5868 12096
rect 5816 12053 5825 12087
rect 5825 12053 5859 12087
rect 5859 12053 5868 12087
rect 5816 12044 5868 12053
rect 6828 12087 6880 12096
rect 6828 12053 6837 12087
rect 6837 12053 6871 12087
rect 6871 12053 6880 12087
rect 6828 12044 6880 12053
rect 7656 12112 7708 12164
rect 10508 12248 10560 12300
rect 9864 12112 9916 12164
rect 13360 12316 13412 12368
rect 16120 12316 16172 12368
rect 12808 12248 12860 12300
rect 18604 12248 18656 12300
rect 19156 12248 19208 12300
rect 19248 12291 19300 12300
rect 19248 12257 19257 12291
rect 19257 12257 19291 12291
rect 19291 12257 19300 12291
rect 19248 12248 19300 12257
rect 19708 12248 19760 12300
rect 11888 12180 11940 12232
rect 13544 12180 13596 12232
rect 19984 12291 20036 12300
rect 19984 12257 19993 12291
rect 19993 12257 20027 12291
rect 20027 12257 20036 12291
rect 19984 12248 20036 12257
rect 20352 12291 20404 12300
rect 20352 12257 20361 12291
rect 20361 12257 20395 12291
rect 20395 12257 20404 12291
rect 20352 12248 20404 12257
rect 13084 12112 13136 12164
rect 13268 12112 13320 12164
rect 19616 12112 19668 12164
rect 8024 12087 8076 12096
rect 8024 12053 8033 12087
rect 8033 12053 8067 12087
rect 8067 12053 8076 12087
rect 8024 12044 8076 12053
rect 8944 12087 8996 12096
rect 8944 12053 8953 12087
rect 8953 12053 8987 12087
rect 8987 12053 8996 12087
rect 8944 12044 8996 12053
rect 9588 12044 9640 12096
rect 11520 12087 11572 12096
rect 11520 12053 11529 12087
rect 11529 12053 11563 12087
rect 11563 12053 11572 12087
rect 11520 12044 11572 12053
rect 12164 12044 12216 12096
rect 13728 12044 13780 12096
rect 14924 12044 14976 12096
rect 16396 12044 16448 12096
rect 20904 12087 20956 12096
rect 20904 12053 20913 12087
rect 20913 12053 20947 12087
rect 20947 12053 20956 12087
rect 20904 12044 20956 12053
rect 3882 11942 3934 11994
rect 3946 11942 3998 11994
rect 4010 11942 4062 11994
rect 4074 11942 4126 11994
rect 4138 11942 4190 11994
rect 10851 11942 10903 11994
rect 10915 11942 10967 11994
rect 10979 11942 11031 11994
rect 11043 11942 11095 11994
rect 11107 11942 11159 11994
rect 17820 11942 17872 11994
rect 17884 11942 17936 11994
rect 17948 11942 18000 11994
rect 18012 11942 18064 11994
rect 18076 11942 18128 11994
rect 24789 11942 24841 11994
rect 24853 11942 24905 11994
rect 24917 11942 24969 11994
rect 24981 11942 25033 11994
rect 25045 11942 25097 11994
rect 3792 11883 3844 11892
rect 3792 11849 3801 11883
rect 3801 11849 3835 11883
rect 3835 11849 3844 11883
rect 3792 11840 3844 11849
rect 5816 11840 5868 11892
rect 6828 11840 6880 11892
rect 5908 11636 5960 11688
rect 6644 11636 6696 11688
rect 8024 11840 8076 11892
rect 9312 11840 9364 11892
rect 9680 11840 9732 11892
rect 10600 11840 10652 11892
rect 11520 11840 11572 11892
rect 9588 11772 9640 11824
rect 9404 11747 9456 11756
rect 7196 11568 7248 11620
rect 8116 11636 8168 11688
rect 9404 11713 9413 11747
rect 9413 11713 9447 11747
rect 9447 11713 9456 11747
rect 9404 11704 9456 11713
rect 9864 11772 9916 11824
rect 9864 11636 9916 11688
rect 9772 11568 9824 11620
rect 13452 11704 13504 11756
rect 13084 11611 13136 11620
rect 6736 11543 6788 11552
rect 6736 11509 6745 11543
rect 6745 11509 6779 11543
rect 6779 11509 6788 11543
rect 6736 11500 6788 11509
rect 7012 11500 7064 11552
rect 9220 11543 9272 11552
rect 9220 11509 9229 11543
rect 9229 11509 9263 11543
rect 9263 11509 9272 11543
rect 9220 11500 9272 11509
rect 10140 11500 10192 11552
rect 10416 11500 10468 11552
rect 11612 11500 11664 11552
rect 13084 11577 13093 11611
rect 13093 11577 13127 11611
rect 13127 11577 13136 11611
rect 13084 11568 13136 11577
rect 13360 11679 13412 11688
rect 13360 11645 13369 11679
rect 13369 11645 13403 11679
rect 13403 11645 13412 11679
rect 13360 11636 13412 11645
rect 14924 11840 14976 11892
rect 14096 11815 14148 11824
rect 14096 11781 14105 11815
rect 14105 11781 14139 11815
rect 14139 11781 14148 11815
rect 14096 11772 14148 11781
rect 14740 11636 14792 11688
rect 15200 11772 15252 11824
rect 18144 11840 18196 11892
rect 15384 11636 15436 11688
rect 19248 11772 19300 11824
rect 19156 11704 19208 11756
rect 22008 11840 22060 11892
rect 18788 11636 18840 11688
rect 20904 11679 20956 11688
rect 20904 11645 20922 11679
rect 20922 11645 20956 11679
rect 20904 11636 20956 11645
rect 14188 11568 14240 11620
rect 15292 11611 15344 11620
rect 15292 11577 15301 11611
rect 15301 11577 15335 11611
rect 15335 11577 15344 11611
rect 15292 11568 15344 11577
rect 13268 11500 13320 11552
rect 13544 11543 13596 11552
rect 13544 11509 13553 11543
rect 13553 11509 13587 11543
rect 13587 11509 13596 11543
rect 13544 11500 13596 11509
rect 15384 11543 15436 11552
rect 15384 11509 15393 11543
rect 15393 11509 15427 11543
rect 15427 11509 15436 11543
rect 15384 11500 15436 11509
rect 15568 11543 15620 11552
rect 15568 11509 15577 11543
rect 15577 11509 15611 11543
rect 15611 11509 15620 11543
rect 15568 11500 15620 11509
rect 16212 11543 16264 11552
rect 16212 11509 16221 11543
rect 16221 11509 16255 11543
rect 16255 11509 16264 11543
rect 16212 11500 16264 11509
rect 7366 11398 7418 11450
rect 7430 11398 7482 11450
rect 7494 11398 7546 11450
rect 7558 11398 7610 11450
rect 7622 11398 7674 11450
rect 14335 11398 14387 11450
rect 14399 11398 14451 11450
rect 14463 11398 14515 11450
rect 14527 11398 14579 11450
rect 14591 11398 14643 11450
rect 21304 11398 21356 11450
rect 21368 11398 21420 11450
rect 21432 11398 21484 11450
rect 21496 11398 21548 11450
rect 21560 11398 21612 11450
rect 28273 11398 28325 11450
rect 28337 11398 28389 11450
rect 28401 11398 28453 11450
rect 28465 11398 28517 11450
rect 28529 11398 28581 11450
rect 6184 11296 6236 11348
rect 8944 11296 8996 11348
rect 9220 11296 9272 11348
rect 6736 11203 6788 11212
rect 6736 11169 6745 11203
rect 6745 11169 6779 11203
rect 6779 11169 6788 11203
rect 6736 11160 6788 11169
rect 7380 10999 7432 11008
rect 7380 10965 7389 10999
rect 7389 10965 7423 10999
rect 7423 10965 7432 10999
rect 7380 10956 7432 10965
rect 8208 11135 8260 11144
rect 8208 11101 8217 11135
rect 8217 11101 8251 11135
rect 8251 11101 8260 11135
rect 8208 11092 8260 11101
rect 8760 11160 8812 11212
rect 9128 11228 9180 11280
rect 10140 11271 10192 11280
rect 10140 11237 10149 11271
rect 10149 11237 10183 11271
rect 10183 11237 10192 11271
rect 10140 11228 10192 11237
rect 11704 11296 11756 11348
rect 13360 11296 13412 11348
rect 14188 11296 14240 11348
rect 9312 11092 9364 11144
rect 9220 11024 9272 11076
rect 10416 11203 10468 11212
rect 10416 11169 10425 11203
rect 10425 11169 10459 11203
rect 10459 11169 10468 11203
rect 10416 11160 10468 11169
rect 11796 11160 11848 11212
rect 11244 11092 11296 11144
rect 14096 11228 14148 11280
rect 14832 11296 14884 11348
rect 15292 11296 15344 11348
rect 15568 11296 15620 11348
rect 16212 11296 16264 11348
rect 15384 11228 15436 11280
rect 14832 11203 14884 11212
rect 14832 11169 14841 11203
rect 14841 11169 14875 11203
rect 14875 11169 14884 11203
rect 14832 11160 14884 11169
rect 15016 11203 15068 11212
rect 15016 11169 15025 11203
rect 15025 11169 15059 11203
rect 15059 11169 15068 11203
rect 15016 11160 15068 11169
rect 16396 11271 16448 11280
rect 16396 11237 16405 11271
rect 16405 11237 16439 11271
rect 16439 11237 16448 11271
rect 16396 11228 16448 11237
rect 10508 11024 10560 11076
rect 11336 11024 11388 11076
rect 14832 11024 14884 11076
rect 16856 11092 16908 11144
rect 10140 10999 10192 11008
rect 10140 10965 10149 10999
rect 10149 10965 10183 10999
rect 10183 10965 10192 10999
rect 10140 10956 10192 10965
rect 16120 10956 16172 11008
rect 18144 11160 18196 11212
rect 16580 10999 16632 11008
rect 16580 10965 16589 10999
rect 16589 10965 16623 10999
rect 16623 10965 16632 10999
rect 16580 10956 16632 10965
rect 3882 10854 3934 10906
rect 3946 10854 3998 10906
rect 4010 10854 4062 10906
rect 4074 10854 4126 10906
rect 4138 10854 4190 10906
rect 10851 10854 10903 10906
rect 10915 10854 10967 10906
rect 10979 10854 11031 10906
rect 11043 10854 11095 10906
rect 11107 10854 11159 10906
rect 17820 10854 17872 10906
rect 17884 10854 17936 10906
rect 17948 10854 18000 10906
rect 18012 10854 18064 10906
rect 18076 10854 18128 10906
rect 24789 10854 24841 10906
rect 24853 10854 24905 10906
rect 24917 10854 24969 10906
rect 24981 10854 25033 10906
rect 25045 10854 25097 10906
rect 7012 10752 7064 10804
rect 11336 10752 11388 10804
rect 11796 10752 11848 10804
rect 16856 10752 16908 10804
rect 11612 10616 11664 10668
rect 16580 10616 16632 10668
rect 6644 10548 6696 10600
rect 7380 10523 7432 10532
rect 7380 10489 7398 10523
rect 7398 10489 7432 10523
rect 7380 10480 7432 10489
rect 11244 10548 11296 10600
rect 17592 10591 17644 10600
rect 17592 10557 17601 10591
rect 17601 10557 17635 10591
rect 17635 10557 17644 10591
rect 17592 10548 17644 10557
rect 10140 10523 10192 10532
rect 10140 10489 10174 10523
rect 10174 10489 10192 10523
rect 10140 10480 10192 10489
rect 7840 10412 7892 10464
rect 7366 10310 7418 10362
rect 7430 10310 7482 10362
rect 7494 10310 7546 10362
rect 7558 10310 7610 10362
rect 7622 10310 7674 10362
rect 14335 10310 14387 10362
rect 14399 10310 14451 10362
rect 14463 10310 14515 10362
rect 14527 10310 14579 10362
rect 14591 10310 14643 10362
rect 21304 10310 21356 10362
rect 21368 10310 21420 10362
rect 21432 10310 21484 10362
rect 21496 10310 21548 10362
rect 21560 10310 21612 10362
rect 28273 10310 28325 10362
rect 28337 10310 28389 10362
rect 28401 10310 28453 10362
rect 28465 10310 28517 10362
rect 28529 10310 28581 10362
rect 9220 10251 9272 10260
rect 9220 10217 9229 10251
rect 9229 10217 9263 10251
rect 9263 10217 9272 10251
rect 9220 10208 9272 10217
rect 8208 10140 8260 10192
rect 7840 10115 7892 10124
rect 7840 10081 7849 10115
rect 7849 10081 7883 10115
rect 7883 10081 7892 10115
rect 7840 10072 7892 10081
rect 3882 9766 3934 9818
rect 3946 9766 3998 9818
rect 4010 9766 4062 9818
rect 4074 9766 4126 9818
rect 4138 9766 4190 9818
rect 10851 9766 10903 9818
rect 10915 9766 10967 9818
rect 10979 9766 11031 9818
rect 11043 9766 11095 9818
rect 11107 9766 11159 9818
rect 17820 9766 17872 9818
rect 17884 9766 17936 9818
rect 17948 9766 18000 9818
rect 18012 9766 18064 9818
rect 18076 9766 18128 9818
rect 24789 9766 24841 9818
rect 24853 9766 24905 9818
rect 24917 9766 24969 9818
rect 24981 9766 25033 9818
rect 25045 9766 25097 9818
rect 7366 9222 7418 9274
rect 7430 9222 7482 9274
rect 7494 9222 7546 9274
rect 7558 9222 7610 9274
rect 7622 9222 7674 9274
rect 14335 9222 14387 9274
rect 14399 9222 14451 9274
rect 14463 9222 14515 9274
rect 14527 9222 14579 9274
rect 14591 9222 14643 9274
rect 21304 9222 21356 9274
rect 21368 9222 21420 9274
rect 21432 9222 21484 9274
rect 21496 9222 21548 9274
rect 21560 9222 21612 9274
rect 28273 9222 28325 9274
rect 28337 9222 28389 9274
rect 28401 9222 28453 9274
rect 28465 9222 28517 9274
rect 28529 9222 28581 9274
rect 3882 8678 3934 8730
rect 3946 8678 3998 8730
rect 4010 8678 4062 8730
rect 4074 8678 4126 8730
rect 4138 8678 4190 8730
rect 10851 8678 10903 8730
rect 10915 8678 10967 8730
rect 10979 8678 11031 8730
rect 11043 8678 11095 8730
rect 11107 8678 11159 8730
rect 17820 8678 17872 8730
rect 17884 8678 17936 8730
rect 17948 8678 18000 8730
rect 18012 8678 18064 8730
rect 18076 8678 18128 8730
rect 24789 8678 24841 8730
rect 24853 8678 24905 8730
rect 24917 8678 24969 8730
rect 24981 8678 25033 8730
rect 25045 8678 25097 8730
rect 7366 8134 7418 8186
rect 7430 8134 7482 8186
rect 7494 8134 7546 8186
rect 7558 8134 7610 8186
rect 7622 8134 7674 8186
rect 14335 8134 14387 8186
rect 14399 8134 14451 8186
rect 14463 8134 14515 8186
rect 14527 8134 14579 8186
rect 14591 8134 14643 8186
rect 21304 8134 21356 8186
rect 21368 8134 21420 8186
rect 21432 8134 21484 8186
rect 21496 8134 21548 8186
rect 21560 8134 21612 8186
rect 28273 8134 28325 8186
rect 28337 8134 28389 8186
rect 28401 8134 28453 8186
rect 28465 8134 28517 8186
rect 28529 8134 28581 8186
rect 3882 7590 3934 7642
rect 3946 7590 3998 7642
rect 4010 7590 4062 7642
rect 4074 7590 4126 7642
rect 4138 7590 4190 7642
rect 10851 7590 10903 7642
rect 10915 7590 10967 7642
rect 10979 7590 11031 7642
rect 11043 7590 11095 7642
rect 11107 7590 11159 7642
rect 17820 7590 17872 7642
rect 17884 7590 17936 7642
rect 17948 7590 18000 7642
rect 18012 7590 18064 7642
rect 18076 7590 18128 7642
rect 24789 7590 24841 7642
rect 24853 7590 24905 7642
rect 24917 7590 24969 7642
rect 24981 7590 25033 7642
rect 25045 7590 25097 7642
rect 7366 7046 7418 7098
rect 7430 7046 7482 7098
rect 7494 7046 7546 7098
rect 7558 7046 7610 7098
rect 7622 7046 7674 7098
rect 14335 7046 14387 7098
rect 14399 7046 14451 7098
rect 14463 7046 14515 7098
rect 14527 7046 14579 7098
rect 14591 7046 14643 7098
rect 21304 7046 21356 7098
rect 21368 7046 21420 7098
rect 21432 7046 21484 7098
rect 21496 7046 21548 7098
rect 21560 7046 21612 7098
rect 28273 7046 28325 7098
rect 28337 7046 28389 7098
rect 28401 7046 28453 7098
rect 28465 7046 28517 7098
rect 28529 7046 28581 7098
rect 3882 6502 3934 6554
rect 3946 6502 3998 6554
rect 4010 6502 4062 6554
rect 4074 6502 4126 6554
rect 4138 6502 4190 6554
rect 10851 6502 10903 6554
rect 10915 6502 10967 6554
rect 10979 6502 11031 6554
rect 11043 6502 11095 6554
rect 11107 6502 11159 6554
rect 17820 6502 17872 6554
rect 17884 6502 17936 6554
rect 17948 6502 18000 6554
rect 18012 6502 18064 6554
rect 18076 6502 18128 6554
rect 24789 6502 24841 6554
rect 24853 6502 24905 6554
rect 24917 6502 24969 6554
rect 24981 6502 25033 6554
rect 25045 6502 25097 6554
rect 7366 5958 7418 6010
rect 7430 5958 7482 6010
rect 7494 5958 7546 6010
rect 7558 5958 7610 6010
rect 7622 5958 7674 6010
rect 14335 5958 14387 6010
rect 14399 5958 14451 6010
rect 14463 5958 14515 6010
rect 14527 5958 14579 6010
rect 14591 5958 14643 6010
rect 21304 5958 21356 6010
rect 21368 5958 21420 6010
rect 21432 5958 21484 6010
rect 21496 5958 21548 6010
rect 21560 5958 21612 6010
rect 28273 5958 28325 6010
rect 28337 5958 28389 6010
rect 28401 5958 28453 6010
rect 28465 5958 28517 6010
rect 28529 5958 28581 6010
rect 3882 5414 3934 5466
rect 3946 5414 3998 5466
rect 4010 5414 4062 5466
rect 4074 5414 4126 5466
rect 4138 5414 4190 5466
rect 10851 5414 10903 5466
rect 10915 5414 10967 5466
rect 10979 5414 11031 5466
rect 11043 5414 11095 5466
rect 11107 5414 11159 5466
rect 17820 5414 17872 5466
rect 17884 5414 17936 5466
rect 17948 5414 18000 5466
rect 18012 5414 18064 5466
rect 18076 5414 18128 5466
rect 24789 5414 24841 5466
rect 24853 5414 24905 5466
rect 24917 5414 24969 5466
rect 24981 5414 25033 5466
rect 25045 5414 25097 5466
rect 7366 4870 7418 4922
rect 7430 4870 7482 4922
rect 7494 4870 7546 4922
rect 7558 4870 7610 4922
rect 7622 4870 7674 4922
rect 14335 4870 14387 4922
rect 14399 4870 14451 4922
rect 14463 4870 14515 4922
rect 14527 4870 14579 4922
rect 14591 4870 14643 4922
rect 21304 4870 21356 4922
rect 21368 4870 21420 4922
rect 21432 4870 21484 4922
rect 21496 4870 21548 4922
rect 21560 4870 21612 4922
rect 28273 4870 28325 4922
rect 28337 4870 28389 4922
rect 28401 4870 28453 4922
rect 28465 4870 28517 4922
rect 28529 4870 28581 4922
rect 3882 4326 3934 4378
rect 3946 4326 3998 4378
rect 4010 4326 4062 4378
rect 4074 4326 4126 4378
rect 4138 4326 4190 4378
rect 10851 4326 10903 4378
rect 10915 4326 10967 4378
rect 10979 4326 11031 4378
rect 11043 4326 11095 4378
rect 11107 4326 11159 4378
rect 17820 4326 17872 4378
rect 17884 4326 17936 4378
rect 17948 4326 18000 4378
rect 18012 4326 18064 4378
rect 18076 4326 18128 4378
rect 24789 4326 24841 4378
rect 24853 4326 24905 4378
rect 24917 4326 24969 4378
rect 24981 4326 25033 4378
rect 25045 4326 25097 4378
rect 7366 3782 7418 3834
rect 7430 3782 7482 3834
rect 7494 3782 7546 3834
rect 7558 3782 7610 3834
rect 7622 3782 7674 3834
rect 14335 3782 14387 3834
rect 14399 3782 14451 3834
rect 14463 3782 14515 3834
rect 14527 3782 14579 3834
rect 14591 3782 14643 3834
rect 21304 3782 21356 3834
rect 21368 3782 21420 3834
rect 21432 3782 21484 3834
rect 21496 3782 21548 3834
rect 21560 3782 21612 3834
rect 28273 3782 28325 3834
rect 28337 3782 28389 3834
rect 28401 3782 28453 3834
rect 28465 3782 28517 3834
rect 28529 3782 28581 3834
rect 3882 3238 3934 3290
rect 3946 3238 3998 3290
rect 4010 3238 4062 3290
rect 4074 3238 4126 3290
rect 4138 3238 4190 3290
rect 10851 3238 10903 3290
rect 10915 3238 10967 3290
rect 10979 3238 11031 3290
rect 11043 3238 11095 3290
rect 11107 3238 11159 3290
rect 17820 3238 17872 3290
rect 17884 3238 17936 3290
rect 17948 3238 18000 3290
rect 18012 3238 18064 3290
rect 18076 3238 18128 3290
rect 24789 3238 24841 3290
rect 24853 3238 24905 3290
rect 24917 3238 24969 3290
rect 24981 3238 25033 3290
rect 25045 3238 25097 3290
rect 7366 2694 7418 2746
rect 7430 2694 7482 2746
rect 7494 2694 7546 2746
rect 7558 2694 7610 2746
rect 7622 2694 7674 2746
rect 14335 2694 14387 2746
rect 14399 2694 14451 2746
rect 14463 2694 14515 2746
rect 14527 2694 14579 2746
rect 14591 2694 14643 2746
rect 21304 2694 21356 2746
rect 21368 2694 21420 2746
rect 21432 2694 21484 2746
rect 21496 2694 21548 2746
rect 21560 2694 21612 2746
rect 28273 2694 28325 2746
rect 28337 2694 28389 2746
rect 28401 2694 28453 2746
rect 28465 2694 28517 2746
rect 28529 2694 28581 2746
rect 3882 2150 3934 2202
rect 3946 2150 3998 2202
rect 4010 2150 4062 2202
rect 4074 2150 4126 2202
rect 4138 2150 4190 2202
rect 10851 2150 10903 2202
rect 10915 2150 10967 2202
rect 10979 2150 11031 2202
rect 11043 2150 11095 2202
rect 11107 2150 11159 2202
rect 17820 2150 17872 2202
rect 17884 2150 17936 2202
rect 17948 2150 18000 2202
rect 18012 2150 18064 2202
rect 18076 2150 18128 2202
rect 24789 2150 24841 2202
rect 24853 2150 24905 2202
rect 24917 2150 24969 2202
rect 24981 2150 25033 2202
rect 25045 2150 25097 2202
rect 7366 1606 7418 1658
rect 7430 1606 7482 1658
rect 7494 1606 7546 1658
rect 7558 1606 7610 1658
rect 7622 1606 7674 1658
rect 14335 1606 14387 1658
rect 14399 1606 14451 1658
rect 14463 1606 14515 1658
rect 14527 1606 14579 1658
rect 14591 1606 14643 1658
rect 21304 1606 21356 1658
rect 21368 1606 21420 1658
rect 21432 1606 21484 1658
rect 21496 1606 21548 1658
rect 21560 1606 21612 1658
rect 28273 1606 28325 1658
rect 28337 1606 28389 1658
rect 28401 1606 28453 1658
rect 28465 1606 28517 1658
rect 28529 1606 28581 1658
rect 3882 1062 3934 1114
rect 3946 1062 3998 1114
rect 4010 1062 4062 1114
rect 4074 1062 4126 1114
rect 4138 1062 4190 1114
rect 10851 1062 10903 1114
rect 10915 1062 10967 1114
rect 10979 1062 11031 1114
rect 11043 1062 11095 1114
rect 11107 1062 11159 1114
rect 17820 1062 17872 1114
rect 17884 1062 17936 1114
rect 17948 1062 18000 1114
rect 18012 1062 18064 1114
rect 18076 1062 18128 1114
rect 24789 1062 24841 1114
rect 24853 1062 24905 1114
rect 24917 1062 24969 1114
rect 24981 1062 25033 1114
rect 25045 1062 25097 1114
rect 7366 518 7418 570
rect 7430 518 7482 570
rect 7494 518 7546 570
rect 7558 518 7610 570
rect 7622 518 7674 570
rect 14335 518 14387 570
rect 14399 518 14451 570
rect 14463 518 14515 570
rect 14527 518 14579 570
rect 14591 518 14643 570
rect 21304 518 21356 570
rect 21368 518 21420 570
rect 21432 518 21484 570
rect 21496 518 21548 570
rect 21560 518 21612 570
rect 28273 518 28325 570
rect 28337 518 28389 570
rect 28401 518 28453 570
rect 28465 518 28517 570
rect 28529 518 28581 570
<< metal2 >>
rect 1306 28600 1362 29000
rect 3330 28600 3386 29000
rect 5354 28600 5410 29000
rect 7378 28600 7434 29000
rect 9402 28600 9458 29000
rect 11426 28600 11482 29000
rect 13450 28600 13506 29000
rect 15474 28600 15530 29000
rect 17498 28600 17554 29000
rect 19522 28600 19578 29000
rect 21546 28600 21602 29000
rect 23570 28600 23626 29000
rect 25594 28600 25650 29000
rect 27618 28600 27674 29000
rect 1320 27606 1348 28600
rect 3344 27606 3372 28600
rect 3882 28316 4190 28325
rect 3882 28314 3888 28316
rect 3944 28314 3968 28316
rect 4024 28314 4048 28316
rect 4104 28314 4128 28316
rect 4184 28314 4190 28316
rect 3944 28262 3946 28314
rect 4126 28262 4128 28314
rect 3882 28260 3888 28262
rect 3944 28260 3968 28262
rect 4024 28260 4048 28262
rect 4104 28260 4128 28262
rect 4184 28260 4190 28262
rect 3882 28251 4190 28260
rect 5368 27606 5396 28600
rect 7392 27962 7420 28600
rect 7300 27934 7420 27962
rect 1308 27600 1360 27606
rect 1308 27542 1360 27548
rect 3332 27600 3384 27606
rect 3332 27542 3384 27548
rect 5356 27600 5408 27606
rect 5356 27542 5408 27548
rect 2228 27532 2280 27538
rect 2228 27474 2280 27480
rect 2596 27532 2648 27538
rect 2596 27474 2648 27480
rect 4896 27532 4948 27538
rect 4896 27474 4948 27480
rect 5540 27532 5592 27538
rect 5540 27474 5592 27480
rect 5908 27532 5960 27538
rect 5908 27474 5960 27480
rect 7012 27532 7064 27538
rect 7012 27474 7064 27480
rect 1400 25832 1452 25838
rect 1400 25774 1452 25780
rect 1308 24268 1360 24274
rect 1308 24210 1360 24216
rect 1124 24064 1176 24070
rect 1124 24006 1176 24012
rect 1136 23594 1164 24006
rect 1124 23588 1176 23594
rect 1124 23530 1176 23536
rect 1216 23520 1268 23526
rect 1216 23462 1268 23468
rect 1228 22094 1256 23462
rect 1320 23322 1348 24210
rect 1412 24206 1440 25774
rect 2136 24268 2188 24274
rect 2136 24210 2188 24216
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1412 23662 1440 24142
rect 2148 23866 2176 24210
rect 2136 23860 2188 23866
rect 2136 23802 2188 23808
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1308 23316 1360 23322
rect 1308 23258 1360 23264
rect 1768 23248 1820 23254
rect 1768 23190 1820 23196
rect 2136 23248 2188 23254
rect 2136 23190 2188 23196
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1136 22066 1256 22094
rect 1492 22092 1544 22098
rect 1136 21486 1164 22066
rect 1492 22034 1544 22040
rect 1124 21480 1176 21486
rect 1124 21422 1176 21428
rect 1136 19922 1164 21422
rect 1504 20806 1532 22034
rect 1688 21010 1716 22918
rect 1780 22778 1808 23190
rect 2148 22778 2176 23190
rect 2240 23089 2268 27474
rect 2320 27464 2372 27470
rect 2320 27406 2372 27412
rect 2332 25838 2360 27406
rect 2608 27130 2636 27474
rect 4344 27464 4396 27470
rect 4344 27406 4396 27412
rect 3700 27328 3752 27334
rect 3700 27270 3752 27276
rect 2596 27124 2648 27130
rect 2596 27066 2648 27072
rect 3712 27062 3740 27270
rect 3882 27228 4190 27237
rect 3882 27226 3888 27228
rect 3944 27226 3968 27228
rect 4024 27226 4048 27228
rect 4104 27226 4128 27228
rect 4184 27226 4190 27228
rect 3944 27174 3946 27226
rect 4126 27174 4128 27226
rect 3882 27172 3888 27174
rect 3944 27172 3968 27174
rect 4024 27172 4048 27174
rect 4104 27172 4128 27174
rect 4184 27172 4190 27174
rect 3882 27163 4190 27172
rect 3700 27056 3752 27062
rect 3752 27004 3832 27010
rect 3700 26998 3832 27004
rect 3712 26982 3832 26998
rect 3700 26920 3752 26926
rect 3700 26862 3752 26868
rect 2320 25832 2372 25838
rect 2320 25774 2372 25780
rect 2412 25764 2464 25770
rect 2412 25706 2464 25712
rect 2424 25498 2452 25706
rect 3148 25696 3200 25702
rect 3148 25638 3200 25644
rect 3160 25498 3188 25638
rect 3712 25498 3740 26862
rect 2412 25492 2464 25498
rect 2412 25434 2464 25440
rect 3148 25492 3200 25498
rect 3700 25492 3752 25498
rect 3200 25452 3372 25480
rect 3148 25434 3200 25440
rect 3344 25362 3372 25452
rect 3700 25434 3752 25440
rect 3332 25356 3384 25362
rect 3332 25298 3384 25304
rect 3804 25294 3832 26982
rect 4356 26790 4384 27406
rect 4436 27328 4488 27334
rect 4436 27270 4488 27276
rect 4252 26784 4304 26790
rect 4252 26726 4304 26732
rect 4344 26784 4396 26790
rect 4344 26726 4396 26732
rect 3882 26140 4190 26149
rect 3882 26138 3888 26140
rect 3944 26138 3968 26140
rect 4024 26138 4048 26140
rect 4104 26138 4128 26140
rect 4184 26138 4190 26140
rect 3944 26086 3946 26138
rect 4126 26086 4128 26138
rect 3882 26084 3888 26086
rect 3944 26084 3968 26086
rect 4024 26084 4048 26086
rect 4104 26084 4128 26086
rect 4184 26084 4190 26086
rect 3882 26075 4190 26084
rect 3792 25288 3844 25294
rect 3792 25230 3844 25236
rect 3804 24886 3832 25230
rect 4264 25140 4292 26726
rect 4356 25498 4384 26726
rect 4448 26246 4476 27270
rect 4528 27124 4580 27130
rect 4528 27066 4580 27072
rect 4540 26382 4568 27066
rect 4908 27062 4936 27474
rect 4988 27328 5040 27334
rect 4988 27270 5040 27276
rect 4896 27056 4948 27062
rect 4896 26998 4948 27004
rect 5000 26586 5028 27270
rect 4988 26580 5040 26586
rect 4988 26522 5040 26528
rect 4528 26376 4580 26382
rect 4528 26318 4580 26324
rect 4436 26240 4488 26246
rect 4436 26182 4488 26188
rect 4344 25492 4396 25498
rect 4344 25434 4396 25440
rect 4344 25152 4396 25158
rect 4264 25112 4344 25140
rect 4344 25094 4396 25100
rect 3882 25052 4190 25061
rect 3882 25050 3888 25052
rect 3944 25050 3968 25052
rect 4024 25050 4048 25052
rect 4104 25050 4128 25052
rect 4184 25050 4190 25052
rect 3944 24998 3946 25050
rect 4126 24998 4128 25050
rect 3882 24996 3888 24998
rect 3944 24996 3968 24998
rect 4024 24996 4048 24998
rect 4104 24996 4128 24998
rect 4184 24996 4190 24998
rect 3882 24987 4190 24996
rect 3792 24880 3844 24886
rect 3792 24822 3844 24828
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3700 24268 3752 24274
rect 3700 24210 3752 24216
rect 2872 23656 2924 23662
rect 2872 23598 2924 23604
rect 2412 23520 2464 23526
rect 2412 23462 2464 23468
rect 2424 23118 2452 23462
rect 2412 23112 2464 23118
rect 2226 23080 2282 23089
rect 2412 23054 2464 23060
rect 2226 23015 2282 23024
rect 1768 22772 1820 22778
rect 1768 22714 1820 22720
rect 2136 22772 2188 22778
rect 2136 22714 2188 22720
rect 2424 22574 2452 23054
rect 2884 23050 2912 23598
rect 3528 23322 3556 24210
rect 3712 23866 3740 24210
rect 4252 24064 4304 24070
rect 4252 24006 4304 24012
rect 3882 23964 4190 23973
rect 3882 23962 3888 23964
rect 3944 23962 3968 23964
rect 4024 23962 4048 23964
rect 4104 23962 4128 23964
rect 4184 23962 4190 23964
rect 3944 23910 3946 23962
rect 4126 23910 4128 23962
rect 3882 23908 3888 23910
rect 3944 23908 3968 23910
rect 4024 23908 4048 23910
rect 4104 23908 4128 23910
rect 4184 23908 4190 23910
rect 3882 23899 4190 23908
rect 4264 23866 4292 24006
rect 3700 23860 3752 23866
rect 3700 23802 3752 23808
rect 4252 23860 4304 23866
rect 4252 23802 4304 23808
rect 4252 23656 4304 23662
rect 4356 23644 4384 25094
rect 4304 23616 4384 23644
rect 4252 23598 4304 23604
rect 3700 23588 3752 23594
rect 3700 23530 3752 23536
rect 3608 23520 3660 23526
rect 3608 23462 3660 23468
rect 3516 23316 3568 23322
rect 3516 23258 3568 23264
rect 3240 23248 3292 23254
rect 3240 23190 3292 23196
rect 2872 23044 2924 23050
rect 2872 22986 2924 22992
rect 3252 22778 3280 23190
rect 3240 22772 3292 22778
rect 3240 22714 3292 22720
rect 2412 22568 2464 22574
rect 2412 22510 2464 22516
rect 3424 22568 3476 22574
rect 3424 22510 3476 22516
rect 3436 22438 3464 22510
rect 3620 22506 3648 23462
rect 3712 22778 3740 23530
rect 4540 23254 4568 26318
rect 4712 25764 4764 25770
rect 4712 25706 4764 25712
rect 4724 25498 4752 25706
rect 4712 25492 4764 25498
rect 4712 25434 4764 25440
rect 4896 25356 4948 25362
rect 4896 25298 4948 25304
rect 5448 25356 5500 25362
rect 5448 25298 5500 25304
rect 4908 23866 4936 25298
rect 5460 25158 5488 25298
rect 5356 25152 5408 25158
rect 5356 25094 5408 25100
rect 5448 25152 5500 25158
rect 5448 25094 5500 25100
rect 5368 24410 5396 25094
rect 5356 24404 5408 24410
rect 5356 24346 5408 24352
rect 5356 24200 5408 24206
rect 5356 24142 5408 24148
rect 5368 24070 5396 24142
rect 5264 24064 5316 24070
rect 5264 24006 5316 24012
rect 5356 24064 5408 24070
rect 5356 24006 5408 24012
rect 4896 23860 4948 23866
rect 4896 23802 4948 23808
rect 5276 23662 5304 24006
rect 5264 23656 5316 23662
rect 5264 23598 5316 23604
rect 4528 23248 4580 23254
rect 4528 23190 4580 23196
rect 4436 23180 4488 23186
rect 4436 23122 4488 23128
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 3792 22976 3844 22982
rect 3792 22918 3844 22924
rect 3804 22778 3832 22918
rect 3882 22876 4190 22885
rect 3882 22874 3888 22876
rect 3944 22874 3968 22876
rect 4024 22874 4048 22876
rect 4104 22874 4128 22876
rect 4184 22874 4190 22876
rect 3944 22822 3946 22874
rect 4126 22822 4128 22874
rect 3882 22820 3888 22822
rect 3944 22820 3968 22822
rect 4024 22820 4048 22822
rect 4104 22820 4128 22822
rect 4184 22820 4190 22822
rect 3882 22811 4190 22820
rect 3700 22772 3752 22778
rect 3700 22714 3752 22720
rect 3792 22772 3844 22778
rect 3792 22714 3844 22720
rect 4342 22536 4398 22545
rect 3608 22500 3660 22506
rect 4342 22471 4344 22480
rect 3608 22442 3660 22448
rect 4396 22471 4398 22480
rect 4344 22442 4396 22448
rect 3424 22432 3476 22438
rect 3424 22374 3476 22380
rect 1860 22092 1912 22098
rect 1860 22034 1912 22040
rect 1768 21888 1820 21894
rect 1768 21830 1820 21836
rect 1780 21486 1808 21830
rect 1768 21480 1820 21486
rect 1768 21422 1820 21428
rect 1872 21146 1900 22034
rect 3436 22030 3464 22374
rect 3424 22024 3476 22030
rect 3424 21966 3476 21972
rect 2044 21888 2096 21894
rect 2044 21830 2096 21836
rect 2412 21888 2464 21894
rect 2412 21830 2464 21836
rect 1860 21140 1912 21146
rect 1860 21082 1912 21088
rect 2056 21010 2084 21830
rect 2424 21690 2452 21830
rect 3882 21788 4190 21797
rect 3882 21786 3888 21788
rect 3944 21786 3968 21788
rect 4024 21786 4048 21788
rect 4104 21786 4128 21788
rect 4184 21786 4190 21788
rect 3944 21734 3946 21786
rect 4126 21734 4128 21786
rect 3882 21732 3888 21734
rect 3944 21732 3968 21734
rect 4024 21732 4048 21734
rect 4104 21732 4128 21734
rect 4184 21732 4190 21734
rect 3882 21723 4190 21732
rect 2412 21684 2464 21690
rect 2412 21626 2464 21632
rect 3056 21412 3108 21418
rect 3056 21354 3108 21360
rect 2872 21344 2924 21350
rect 2872 21286 2924 21292
rect 2884 21010 2912 21286
rect 3068 21146 3096 21354
rect 3332 21344 3384 21350
rect 3332 21286 3384 21292
rect 3056 21140 3108 21146
rect 3056 21082 3108 21088
rect 1676 21004 1728 21010
rect 1676 20946 1728 20952
rect 2044 21004 2096 21010
rect 2044 20946 2096 20952
rect 2872 21004 2924 21010
rect 2872 20946 2924 20952
rect 1492 20800 1544 20806
rect 1492 20742 1544 20748
rect 1124 19916 1176 19922
rect 1124 19858 1176 19864
rect 1504 19718 1532 20742
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 19990 1624 20198
rect 1584 19984 1636 19990
rect 1584 19926 1636 19932
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1504 19446 1532 19654
rect 1688 19514 1716 20946
rect 3344 20874 3372 21286
rect 3332 20868 3384 20874
rect 3332 20810 3384 20816
rect 3700 20800 3752 20806
rect 3700 20742 3752 20748
rect 1952 20392 2004 20398
rect 1952 20334 2004 20340
rect 1964 19514 1992 20334
rect 3608 19984 3660 19990
rect 3608 19926 3660 19932
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 1676 19508 1728 19514
rect 1676 19450 1728 19456
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1492 19440 1544 19446
rect 1492 19382 1544 19388
rect 2884 19242 2912 19654
rect 3620 19417 3648 19926
rect 3712 19514 3740 20742
rect 3882 20700 4190 20709
rect 3882 20698 3888 20700
rect 3944 20698 3968 20700
rect 4024 20698 4048 20700
rect 4104 20698 4128 20700
rect 4184 20698 4190 20700
rect 3944 20646 3946 20698
rect 4126 20646 4128 20698
rect 3882 20644 3888 20646
rect 3944 20644 3968 20646
rect 4024 20644 4048 20646
rect 4104 20644 4128 20646
rect 4184 20644 4190 20646
rect 3882 20635 4190 20644
rect 3792 19780 3844 19786
rect 3792 19722 3844 19728
rect 3700 19508 3752 19514
rect 3700 19450 3752 19456
rect 3606 19408 3662 19417
rect 3606 19343 3608 19352
rect 3660 19343 3662 19352
rect 3608 19314 3660 19320
rect 2872 19236 2924 19242
rect 2872 19178 2924 19184
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2148 18222 2176 19110
rect 3620 18834 3648 19314
rect 3804 19310 3832 19722
rect 3882 19612 4190 19621
rect 3882 19610 3888 19612
rect 3944 19610 3968 19612
rect 4024 19610 4048 19612
rect 4104 19610 4128 19612
rect 4184 19610 4190 19612
rect 3944 19558 3946 19610
rect 4126 19558 4128 19610
rect 3882 19556 3888 19558
rect 3944 19556 3968 19558
rect 4024 19556 4048 19558
rect 4104 19556 4128 19558
rect 4184 19556 4190 19558
rect 3882 19547 4190 19556
rect 3792 19304 3844 19310
rect 3792 19246 3844 19252
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3988 18970 4016 19246
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3620 18426 3648 18770
rect 3882 18524 4190 18533
rect 3882 18522 3888 18524
rect 3944 18522 3968 18524
rect 4024 18522 4048 18524
rect 4104 18522 4128 18524
rect 4184 18522 4190 18524
rect 3944 18470 3946 18522
rect 4126 18470 4128 18522
rect 3882 18468 3888 18470
rect 3944 18468 3968 18470
rect 4024 18468 4048 18470
rect 4104 18468 4128 18470
rect 4184 18468 4190 18470
rect 3882 18459 4190 18468
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 1584 18216 1636 18222
rect 1584 18158 1636 18164
rect 2136 18216 2188 18222
rect 2136 18158 2188 18164
rect 1596 17678 1624 18158
rect 3700 17740 3752 17746
rect 3700 17682 3752 17688
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1596 16046 1624 17614
rect 3712 17338 3740 17682
rect 3882 17436 4190 17445
rect 3882 17434 3888 17436
rect 3944 17434 3968 17436
rect 4024 17434 4048 17436
rect 4104 17434 4128 17436
rect 4184 17434 4190 17436
rect 3944 17382 3946 17434
rect 4126 17382 4128 17434
rect 3882 17380 3888 17382
rect 3944 17380 3968 17382
rect 4024 17380 4048 17382
rect 4104 17380 4128 17382
rect 4184 17380 4190 17382
rect 3882 17371 4190 17380
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1780 16046 1808 16390
rect 1584 16040 1636 16046
rect 1584 15982 1636 15988
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1596 13462 1624 15982
rect 2148 15706 2176 16594
rect 3240 16108 3292 16114
rect 3240 16050 3292 16056
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1584 13456 1636 13462
rect 1584 13398 1636 13404
rect 1780 13394 1808 13670
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 2056 12986 2084 13806
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 2424 12782 2452 15438
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 3068 13462 3096 14894
rect 3160 14618 3188 15030
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3252 14414 3280 16050
rect 3344 15366 3372 17070
rect 3436 16794 3464 17070
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3882 16348 4190 16357
rect 3882 16346 3888 16348
rect 3944 16346 3968 16348
rect 4024 16346 4048 16348
rect 4104 16346 4128 16348
rect 4184 16346 4190 16348
rect 3944 16294 3946 16346
rect 4126 16294 4128 16346
rect 3882 16292 3888 16294
rect 3944 16292 3968 16294
rect 4024 16292 4048 16294
rect 4104 16292 4128 16294
rect 4184 16292 4190 16294
rect 3882 16283 4190 16292
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3804 15434 3832 15982
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 4264 15706 4292 15846
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 3792 15428 3844 15434
rect 3792 15370 3844 15376
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3804 15042 3832 15370
rect 3882 15260 4190 15269
rect 3882 15258 3888 15260
rect 3944 15258 3968 15260
rect 4024 15258 4048 15260
rect 4104 15258 4128 15260
rect 4184 15258 4190 15260
rect 3944 15206 3946 15258
rect 4126 15206 4128 15258
rect 3882 15204 3888 15206
rect 3944 15204 3968 15206
rect 4024 15204 4048 15206
rect 4104 15204 4128 15206
rect 4184 15204 4190 15206
rect 3882 15195 4190 15204
rect 3804 15014 3924 15042
rect 3896 14958 3924 15014
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3436 14618 3464 14758
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3712 14498 3740 14894
rect 3712 14482 3832 14498
rect 3712 14476 3844 14482
rect 3712 14470 3792 14476
rect 3792 14418 3844 14424
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 3252 13326 3280 13738
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3804 13258 3832 14418
rect 3882 14172 4190 14181
rect 3882 14170 3888 14172
rect 3944 14170 3968 14172
rect 4024 14170 4048 14172
rect 4104 14170 4128 14172
rect 4184 14170 4190 14172
rect 3944 14118 3946 14170
rect 4126 14118 4128 14170
rect 3882 14116 3888 14118
rect 3944 14116 3968 14118
rect 4024 14116 4048 14118
rect 4104 14116 4128 14118
rect 4184 14116 4190 14118
rect 3882 14107 4190 14116
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 4080 13462 4108 13806
rect 4160 13728 4212 13734
rect 4160 13670 4212 13676
rect 4172 13462 4200 13670
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 4160 13456 4212 13462
rect 4160 13398 4212 13404
rect 3516 13252 3568 13258
rect 3516 13194 3568 13200
rect 3792 13252 3844 13258
rect 3792 13194 3844 13200
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3436 12986 3464 13126
rect 3528 12986 3556 13194
rect 3882 13084 4190 13093
rect 3882 13082 3888 13084
rect 3944 13082 3968 13084
rect 4024 13082 4048 13084
rect 4104 13082 4128 13084
rect 4184 13082 4190 13084
rect 3944 13030 3946 13082
rect 4126 13030 4128 13082
rect 3882 13028 3888 13030
rect 3944 13028 3968 13030
rect 4024 13028 4048 13030
rect 4104 13028 4128 13030
rect 4184 13028 4190 13030
rect 3882 13019 4190 13028
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3804 12434 3832 12718
rect 4356 12434 4384 22442
rect 4448 22166 4476 23122
rect 4528 22976 4580 22982
rect 4528 22918 4580 22924
rect 4540 22778 4568 22918
rect 4528 22772 4580 22778
rect 4528 22714 4580 22720
rect 4632 22438 4660 23122
rect 4896 22568 4948 22574
rect 4896 22510 4948 22516
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4908 22234 4936 22510
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 4436 22160 4488 22166
rect 4436 22102 4488 22108
rect 5172 21616 5224 21622
rect 5172 21558 5224 21564
rect 4804 21344 4856 21350
rect 4804 21286 4856 21292
rect 4816 21010 4844 21286
rect 4804 21004 4856 21010
rect 4804 20946 4856 20952
rect 4988 21004 5040 21010
rect 4988 20946 5040 20952
rect 4816 19922 4844 20946
rect 5000 20262 5028 20946
rect 5080 20936 5132 20942
rect 5080 20878 5132 20884
rect 4988 20256 5040 20262
rect 4988 20198 5040 20204
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 4436 19712 4488 19718
rect 4436 19654 4488 19660
rect 4528 19712 4580 19718
rect 4528 19654 4580 19660
rect 4448 19514 4476 19654
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4540 18970 4568 19654
rect 4528 18964 4580 18970
rect 4528 18906 4580 18912
rect 4712 18692 4764 18698
rect 4712 18634 4764 18640
rect 4436 18284 4488 18290
rect 4436 18226 4488 18232
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4448 16182 4476 18226
rect 4632 17542 4660 18226
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4632 16726 4660 17478
rect 4620 16720 4672 16726
rect 4620 16662 4672 16668
rect 4724 16658 4752 18634
rect 4816 16794 4844 19858
rect 5000 19854 5028 20198
rect 5092 19854 5120 20878
rect 4988 19848 5040 19854
rect 4988 19790 5040 19796
rect 5080 19848 5132 19854
rect 5080 19790 5132 19796
rect 5092 19242 5120 19790
rect 4896 19236 4948 19242
rect 4896 19178 4948 19184
rect 5080 19236 5132 19242
rect 5080 19178 5132 19184
rect 4908 18970 4936 19178
rect 4896 18964 4948 18970
rect 4896 18906 4948 18912
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4540 16250 4568 16594
rect 4724 16538 4752 16594
rect 4724 16510 4844 16538
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4436 16176 4488 16182
rect 4436 16118 4488 16124
rect 4448 15162 4476 16118
rect 4620 15972 4672 15978
rect 4620 15914 4672 15920
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4540 14958 4568 15506
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 4540 13870 4568 14894
rect 4632 14414 4660 15914
rect 4724 15910 4752 16390
rect 4816 16046 4844 16510
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4528 13864 4580 13870
rect 4528 13806 4580 13812
rect 4724 13734 4752 15846
rect 4816 13870 4844 15982
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4540 13394 4568 13670
rect 4908 13394 4936 18566
rect 5092 18222 5120 19178
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5184 16776 5212 21558
rect 5276 21146 5304 23598
rect 5368 23186 5396 24006
rect 5356 23180 5408 23186
rect 5356 23122 5408 23128
rect 5356 22568 5408 22574
rect 5354 22536 5356 22545
rect 5408 22536 5410 22545
rect 5354 22471 5410 22480
rect 5356 22160 5408 22166
rect 5356 22102 5408 22108
rect 5368 21622 5396 22102
rect 5552 22094 5580 27474
rect 5920 26382 5948 27474
rect 6092 27464 6144 27470
rect 6092 27406 6144 27412
rect 6000 27328 6052 27334
rect 6000 27270 6052 27276
rect 6012 26926 6040 27270
rect 6000 26920 6052 26926
rect 6000 26862 6052 26868
rect 6104 26586 6132 27406
rect 6920 27396 6972 27402
rect 6920 27338 6972 27344
rect 6276 26920 6328 26926
rect 6276 26862 6328 26868
rect 6092 26580 6144 26586
rect 6092 26522 6144 26528
rect 5908 26376 5960 26382
rect 5908 26318 5960 26324
rect 6000 26036 6052 26042
rect 6000 25978 6052 25984
rect 6012 25702 6040 25978
rect 6288 25838 6316 26862
rect 6828 26444 6880 26450
rect 6828 26386 6880 26392
rect 6552 26376 6604 26382
rect 6552 26318 6604 26324
rect 6368 26308 6420 26314
rect 6368 26250 6420 26256
rect 6276 25832 6328 25838
rect 6276 25774 6328 25780
rect 6000 25696 6052 25702
rect 6000 25638 6052 25644
rect 5908 24676 5960 24682
rect 5908 24618 5960 24624
rect 5920 24206 5948 24618
rect 5908 24200 5960 24206
rect 5908 24142 5960 24148
rect 6012 24154 6040 25638
rect 6012 24138 6224 24154
rect 6012 24132 6236 24138
rect 6012 24126 6184 24132
rect 6012 24070 6040 24126
rect 6184 24074 6236 24080
rect 5816 24064 5868 24070
rect 5816 24006 5868 24012
rect 6000 24064 6052 24070
rect 6000 24006 6052 24012
rect 6092 24064 6144 24070
rect 6092 24006 6144 24012
rect 5828 23866 5856 24006
rect 6104 23866 6132 24006
rect 5816 23860 5868 23866
rect 5816 23802 5868 23808
rect 6092 23860 6144 23866
rect 6092 23802 6144 23808
rect 6196 22778 6224 24074
rect 6000 22772 6052 22778
rect 6000 22714 6052 22720
rect 6184 22772 6236 22778
rect 6184 22714 6236 22720
rect 6012 22438 6040 22714
rect 5816 22432 5868 22438
rect 6000 22432 6052 22438
rect 5816 22374 5868 22380
rect 5920 22392 6000 22420
rect 5828 22234 5856 22374
rect 5816 22228 5868 22234
rect 5816 22170 5868 22176
rect 5552 22066 5764 22094
rect 5356 21616 5408 21622
rect 5356 21558 5408 21564
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5356 21480 5408 21486
rect 5356 21422 5408 21428
rect 5264 21140 5316 21146
rect 5264 21082 5316 21088
rect 5368 20330 5396 21422
rect 5552 21146 5580 21490
rect 5540 21140 5592 21146
rect 5540 21082 5592 21088
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 5356 20324 5408 20330
rect 5356 20266 5408 20272
rect 5460 19310 5488 20946
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5552 19718 5580 20878
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 5644 20398 5672 20742
rect 5736 20505 5764 22066
rect 5816 21412 5868 21418
rect 5816 21354 5868 21360
rect 5828 20602 5856 21354
rect 5816 20596 5868 20602
rect 5816 20538 5868 20544
rect 5722 20496 5778 20505
rect 5722 20431 5778 20440
rect 5632 20392 5684 20398
rect 5632 20334 5684 20340
rect 5724 20324 5776 20330
rect 5724 20266 5776 20272
rect 5736 19854 5764 20266
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5736 19514 5764 19790
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5460 18630 5488 18906
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 5920 18426 5948 22392
rect 6000 22374 6052 22380
rect 6288 21010 6316 25774
rect 6380 25702 6408 26250
rect 6564 26042 6592 26318
rect 6552 26036 6604 26042
rect 6552 25978 6604 25984
rect 6736 25968 6788 25974
rect 6736 25910 6788 25916
rect 6368 25696 6420 25702
rect 6368 25638 6420 25644
rect 6644 25288 6696 25294
rect 6644 25230 6696 25236
rect 6656 24954 6684 25230
rect 6644 24948 6696 24954
rect 6644 24890 6696 24896
rect 6368 24268 6420 24274
rect 6368 24210 6420 24216
rect 6380 22642 6408 24210
rect 6460 24064 6512 24070
rect 6460 24006 6512 24012
rect 6472 23662 6500 24006
rect 6460 23656 6512 23662
rect 6460 23598 6512 23604
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6552 22704 6604 22710
rect 6552 22646 6604 22652
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 6460 22636 6512 22642
rect 6460 22578 6512 22584
rect 6472 22234 6500 22578
rect 6460 22228 6512 22234
rect 6460 22170 6512 22176
rect 6460 21956 6512 21962
rect 6460 21898 6512 21904
rect 6276 21004 6328 21010
rect 6276 20946 6328 20952
rect 6092 20868 6144 20874
rect 6092 20810 6144 20816
rect 6000 20800 6052 20806
rect 6000 20742 6052 20748
rect 6012 20398 6040 20742
rect 6104 20466 6132 20810
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 6000 20392 6052 20398
rect 6000 20334 6052 20340
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 6104 19174 6132 20198
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6196 19417 6224 19858
rect 6472 19718 6500 21898
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6472 19514 6500 19654
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6182 19408 6238 19417
rect 6182 19343 6184 19352
rect 6236 19343 6238 19352
rect 6184 19314 6236 19320
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 6564 18222 6592 22646
rect 6656 22488 6684 23122
rect 6748 23118 6776 25910
rect 6840 25770 6868 26386
rect 6828 25764 6880 25770
rect 6828 25706 6880 25712
rect 6736 23112 6788 23118
rect 6736 23054 6788 23060
rect 6932 22778 6960 27338
rect 7024 25974 7052 27474
rect 7300 27402 7328 27934
rect 7366 27772 7674 27781
rect 7366 27770 7372 27772
rect 7428 27770 7452 27772
rect 7508 27770 7532 27772
rect 7588 27770 7612 27772
rect 7668 27770 7674 27772
rect 7428 27718 7430 27770
rect 7610 27718 7612 27770
rect 7366 27716 7372 27718
rect 7428 27716 7452 27718
rect 7508 27716 7532 27718
rect 7588 27716 7612 27718
rect 7668 27716 7674 27718
rect 7366 27707 7674 27716
rect 7932 27532 7984 27538
rect 7932 27474 7984 27480
rect 8944 27532 8996 27538
rect 8944 27474 8996 27480
rect 7840 27464 7892 27470
rect 7840 27406 7892 27412
rect 7288 27396 7340 27402
rect 7288 27338 7340 27344
rect 7472 27328 7524 27334
rect 7472 27270 7524 27276
rect 7288 26852 7340 26858
rect 7288 26794 7340 26800
rect 7300 26586 7328 26794
rect 7484 26790 7512 27270
rect 7852 27130 7880 27406
rect 7840 27124 7892 27130
rect 7840 27066 7892 27072
rect 7748 27056 7800 27062
rect 7748 26998 7800 27004
rect 7472 26784 7524 26790
rect 7472 26726 7524 26732
rect 7366 26684 7674 26693
rect 7366 26682 7372 26684
rect 7428 26682 7452 26684
rect 7508 26682 7532 26684
rect 7588 26682 7612 26684
rect 7668 26682 7674 26684
rect 7428 26630 7430 26682
rect 7610 26630 7612 26682
rect 7366 26628 7372 26630
rect 7428 26628 7452 26630
rect 7508 26628 7532 26630
rect 7588 26628 7612 26630
rect 7668 26628 7674 26630
rect 7366 26619 7674 26628
rect 7760 26586 7788 26998
rect 7288 26580 7340 26586
rect 7288 26522 7340 26528
rect 7564 26580 7616 26586
rect 7564 26522 7616 26528
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7576 26450 7604 26522
rect 7564 26444 7616 26450
rect 7564 26386 7616 26392
rect 7840 26444 7892 26450
rect 7944 26432 7972 27474
rect 8760 26920 8812 26926
rect 7892 26404 7972 26432
rect 7840 26386 7892 26392
rect 7944 26042 7972 26404
rect 8588 26880 8760 26908
rect 7932 26036 7984 26042
rect 7932 25978 7984 25984
rect 7012 25968 7064 25974
rect 7012 25910 7064 25916
rect 7024 24954 7052 25910
rect 7932 25832 7984 25838
rect 7932 25774 7984 25780
rect 7748 25764 7800 25770
rect 7748 25706 7800 25712
rect 7366 25596 7674 25605
rect 7366 25594 7372 25596
rect 7428 25594 7452 25596
rect 7508 25594 7532 25596
rect 7588 25594 7612 25596
rect 7668 25594 7674 25596
rect 7428 25542 7430 25594
rect 7610 25542 7612 25594
rect 7366 25540 7372 25542
rect 7428 25540 7452 25542
rect 7508 25540 7532 25542
rect 7588 25540 7612 25542
rect 7668 25540 7674 25542
rect 7366 25531 7674 25540
rect 7012 24948 7064 24954
rect 7012 24890 7064 24896
rect 7288 24608 7340 24614
rect 7288 24550 7340 24556
rect 7300 24138 7328 24550
rect 7366 24508 7674 24517
rect 7366 24506 7372 24508
rect 7428 24506 7452 24508
rect 7508 24506 7532 24508
rect 7588 24506 7612 24508
rect 7668 24506 7674 24508
rect 7428 24454 7430 24506
rect 7610 24454 7612 24506
rect 7366 24452 7372 24454
rect 7428 24452 7452 24454
rect 7508 24452 7532 24454
rect 7588 24452 7612 24454
rect 7668 24452 7674 24454
rect 7366 24443 7674 24452
rect 7760 24410 7788 25706
rect 7944 25498 7972 25774
rect 7932 25492 7984 25498
rect 7932 25434 7984 25440
rect 8300 25356 8352 25362
rect 8300 25298 8352 25304
rect 7748 24404 7800 24410
rect 7748 24346 7800 24352
rect 7748 24268 7800 24274
rect 7800 24228 7880 24256
rect 7748 24210 7800 24216
rect 7288 24132 7340 24138
rect 7288 24074 7340 24080
rect 7300 23866 7328 24074
rect 7748 24064 7800 24070
rect 7748 24006 7800 24012
rect 7288 23860 7340 23866
rect 7288 23802 7340 23808
rect 7366 23420 7674 23429
rect 7366 23418 7372 23420
rect 7428 23418 7452 23420
rect 7508 23418 7532 23420
rect 7588 23418 7612 23420
rect 7668 23418 7674 23420
rect 7428 23366 7430 23418
rect 7610 23366 7612 23418
rect 7366 23364 7372 23366
rect 7428 23364 7452 23366
rect 7508 23364 7532 23366
rect 7588 23364 7612 23366
rect 7668 23364 7674 23366
rect 7366 23355 7674 23364
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 7760 22506 7788 24006
rect 7852 23594 7880 24228
rect 7840 23588 7892 23594
rect 7840 23530 7892 23536
rect 7852 23186 7880 23530
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 8312 23118 8340 25298
rect 8300 23112 8352 23118
rect 8300 23054 8352 23060
rect 8024 22568 8076 22574
rect 8024 22510 8076 22516
rect 6736 22500 6788 22506
rect 6656 22460 6736 22488
rect 6656 21894 6684 22460
rect 6736 22442 6788 22448
rect 7748 22500 7800 22506
rect 7748 22442 7800 22448
rect 7366 22332 7674 22341
rect 7366 22330 7372 22332
rect 7428 22330 7452 22332
rect 7508 22330 7532 22332
rect 7588 22330 7612 22332
rect 7668 22330 7674 22332
rect 7428 22278 7430 22330
rect 7610 22278 7612 22330
rect 7366 22276 7372 22278
rect 7428 22276 7452 22278
rect 7508 22276 7532 22278
rect 7588 22276 7612 22278
rect 7668 22276 7674 22278
rect 7366 22267 7674 22276
rect 6736 22092 6788 22098
rect 6736 22034 6788 22040
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6656 19718 6684 21830
rect 6748 21350 6776 22034
rect 7746 21992 7802 22001
rect 7746 21927 7802 21936
rect 6920 21684 6972 21690
rect 6920 21626 6972 21632
rect 6736 21344 6788 21350
rect 6736 21286 6788 21292
rect 6748 20534 6776 21286
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6736 20528 6788 20534
rect 6736 20470 6788 20476
rect 6736 20324 6788 20330
rect 6736 20266 6788 20272
rect 6748 19922 6776 20266
rect 6736 19916 6788 19922
rect 6736 19858 6788 19864
rect 6644 19712 6696 19718
rect 6644 19654 6696 19660
rect 6656 19174 6684 19654
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6748 18834 6776 19858
rect 6840 19310 6868 20538
rect 6932 20398 6960 21626
rect 7760 21486 7788 21927
rect 8036 21554 8064 22510
rect 8300 22500 8352 22506
rect 8300 22442 8352 22448
rect 8312 21894 8340 22442
rect 8484 22092 8536 22098
rect 8484 22034 8536 22040
rect 8300 21888 8352 21894
rect 8300 21830 8352 21836
rect 8312 21690 8340 21830
rect 8300 21684 8352 21690
rect 8300 21626 8352 21632
rect 8024 21548 8076 21554
rect 8024 21490 8076 21496
rect 7012 21480 7064 21486
rect 7012 21422 7064 21428
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 7748 21480 7800 21486
rect 7748 21422 7800 21428
rect 8392 21480 8444 21486
rect 8392 21422 8444 21428
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 7024 20262 7052 21422
rect 7116 20398 7144 21422
rect 7366 21244 7674 21253
rect 7366 21242 7372 21244
rect 7428 21242 7452 21244
rect 7508 21242 7532 21244
rect 7588 21242 7612 21244
rect 7668 21242 7674 21244
rect 7428 21190 7430 21242
rect 7610 21190 7612 21242
rect 7366 21188 7372 21190
rect 7428 21188 7452 21190
rect 7508 21188 7532 21190
rect 7588 21188 7612 21190
rect 7668 21188 7674 21190
rect 7366 21179 7674 21188
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 7196 20460 7248 20466
rect 7196 20402 7248 20408
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 7116 20074 7144 20334
rect 7208 20262 7236 20402
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7024 20058 7144 20074
rect 7012 20052 7144 20058
rect 7064 20046 7144 20052
rect 7012 19994 7064 20000
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 6932 19514 6960 19858
rect 7300 19854 7328 20402
rect 7366 20156 7674 20165
rect 7366 20154 7372 20156
rect 7428 20154 7452 20156
rect 7508 20154 7532 20156
rect 7588 20154 7612 20156
rect 7668 20154 7674 20156
rect 7428 20102 7430 20154
rect 7610 20102 7612 20154
rect 7366 20100 7372 20102
rect 7428 20100 7452 20102
rect 7508 20100 7532 20102
rect 7588 20100 7612 20102
rect 7668 20100 7674 20102
rect 7366 20091 7674 20100
rect 7380 19984 7432 19990
rect 7380 19926 7432 19932
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 6920 19508 6972 19514
rect 6920 19450 6972 19456
rect 7392 19446 7420 19926
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 8024 19712 8076 19718
rect 8024 19654 8076 19660
rect 7380 19440 7432 19446
rect 7380 19382 7432 19388
rect 8036 19378 8064 19654
rect 8128 19514 8156 19858
rect 8220 19514 8248 20946
rect 8404 20466 8432 21422
rect 8496 20466 8524 22034
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 8588 19990 8616 26880
rect 8760 26862 8812 26868
rect 8668 25832 8720 25838
rect 8668 25774 8720 25780
rect 8680 25498 8708 25774
rect 8760 25696 8812 25702
rect 8760 25638 8812 25644
rect 8772 25498 8800 25638
rect 8956 25498 8984 27474
rect 9416 27130 9444 28600
rect 10851 28316 11159 28325
rect 10851 28314 10857 28316
rect 10913 28314 10937 28316
rect 10993 28314 11017 28316
rect 11073 28314 11097 28316
rect 11153 28314 11159 28316
rect 10913 28262 10915 28314
rect 11095 28262 11097 28314
rect 10851 28260 10857 28262
rect 10913 28260 10937 28262
rect 10993 28260 11017 28262
rect 11073 28260 11097 28262
rect 11153 28260 11159 28262
rect 10851 28251 11159 28260
rect 11440 28218 11468 28600
rect 11428 28212 11480 28218
rect 11428 28154 11480 28160
rect 11152 28008 11204 28014
rect 11152 27950 11204 27956
rect 9496 27532 9548 27538
rect 9496 27474 9548 27480
rect 9956 27532 10008 27538
rect 9956 27474 10008 27480
rect 9404 27124 9456 27130
rect 9404 27066 9456 27072
rect 8668 25492 8720 25498
rect 8668 25434 8720 25440
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 8944 25492 8996 25498
rect 8944 25434 8996 25440
rect 8668 25288 8720 25294
rect 8668 25230 8720 25236
rect 8680 24410 8708 25230
rect 9508 24750 9536 27474
rect 9588 25152 9640 25158
rect 9588 25094 9640 25100
rect 9600 24750 9628 25094
rect 9864 24948 9916 24954
rect 9864 24890 9916 24896
rect 9496 24744 9548 24750
rect 9496 24686 9548 24692
rect 9588 24744 9640 24750
rect 9588 24686 9640 24692
rect 8668 24404 8720 24410
rect 8668 24346 8720 24352
rect 9220 24404 9272 24410
rect 9220 24346 9272 24352
rect 9036 24064 9088 24070
rect 9036 24006 9088 24012
rect 9048 23866 9076 24006
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 9128 23860 9180 23866
rect 9128 23802 9180 23808
rect 9140 23746 9168 23802
rect 9232 23798 9260 24346
rect 8864 23718 9168 23746
rect 9220 23792 9272 23798
rect 9220 23734 9272 23740
rect 8864 23526 8892 23718
rect 9232 23662 9260 23734
rect 9036 23656 9088 23662
rect 9036 23598 9088 23604
rect 9220 23656 9272 23662
rect 9220 23598 9272 23604
rect 9404 23656 9456 23662
rect 9404 23598 9456 23604
rect 8852 23520 8904 23526
rect 8852 23462 8904 23468
rect 8944 23520 8996 23526
rect 8944 23462 8996 23468
rect 8760 23248 8812 23254
rect 8760 23190 8812 23196
rect 8668 23180 8720 23186
rect 8668 23122 8720 23128
rect 8680 22094 8708 23122
rect 8772 22760 8800 23190
rect 8956 22982 8984 23462
rect 9048 23254 9076 23598
rect 9036 23248 9088 23254
rect 9036 23190 9088 23196
rect 8944 22976 8996 22982
rect 8944 22918 8996 22924
rect 8944 22772 8996 22778
rect 8772 22732 8944 22760
rect 8944 22714 8996 22720
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8772 22438 8800 22578
rect 8760 22432 8812 22438
rect 8760 22374 8812 22380
rect 8944 22432 8996 22438
rect 8944 22374 8996 22380
rect 8956 22234 8984 22374
rect 8944 22228 8996 22234
rect 8944 22170 8996 22176
rect 9232 22094 9260 23598
rect 9416 23322 9444 23598
rect 9404 23316 9456 23322
rect 9404 23258 9456 23264
rect 9508 23186 9536 24686
rect 9600 24138 9628 24686
rect 9588 24132 9640 24138
rect 9588 24074 9640 24080
rect 9772 24064 9824 24070
rect 9772 24006 9824 24012
rect 9784 23730 9812 24006
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 9692 23254 9720 23462
rect 9680 23248 9732 23254
rect 9680 23190 9732 23196
rect 9496 23180 9548 23186
rect 9496 23122 9548 23128
rect 8680 22066 8800 22094
rect 8668 21888 8720 21894
rect 8668 21830 8720 21836
rect 8680 21486 8708 21830
rect 8668 21480 8720 21486
rect 8668 21422 8720 21428
rect 8576 19984 8628 19990
rect 8576 19926 8628 19932
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 7366 19068 7674 19077
rect 7366 19066 7372 19068
rect 7428 19066 7452 19068
rect 7508 19066 7532 19068
rect 7588 19066 7612 19068
rect 7668 19066 7674 19068
rect 7428 19014 7430 19066
rect 7610 19014 7612 19066
rect 7366 19012 7372 19014
rect 7428 19012 7452 19014
rect 7508 19012 7532 19014
rect 7588 19012 7612 19014
rect 7668 19012 7674 19014
rect 7366 19003 7674 19012
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 7024 18222 7052 18566
rect 6276 18216 6328 18222
rect 6276 18158 6328 18164
rect 6552 18216 6604 18222
rect 7012 18216 7064 18222
rect 6552 18158 6604 18164
rect 6932 18176 7012 18204
rect 5816 18148 5868 18154
rect 5816 18090 5868 18096
rect 5828 17746 5856 18090
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 5816 17740 5868 17746
rect 5816 17682 5868 17688
rect 5092 16748 5212 16776
rect 5092 13802 5120 16748
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 5184 15502 5212 16594
rect 6012 16590 6040 18022
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 5368 16046 5396 16526
rect 6104 16522 6132 17682
rect 6288 17542 6316 18158
rect 6564 17746 6592 18158
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6276 17536 6328 17542
rect 6276 17478 6328 17484
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6276 16720 6328 16726
rect 6328 16680 6500 16708
rect 6276 16662 6328 16668
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6196 16538 6224 16594
rect 6196 16522 6408 16538
rect 6092 16516 6144 16522
rect 6196 16516 6420 16522
rect 6196 16510 6368 16516
rect 6092 16458 6144 16464
rect 6368 16458 6420 16464
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 5724 15972 5776 15978
rect 5724 15914 5776 15920
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 5184 14958 5212 15438
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5460 14550 5488 15506
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 5736 13870 5764 15914
rect 6104 15570 6132 15914
rect 6380 15570 6408 15982
rect 6472 15706 6500 16680
rect 6564 16590 6592 16934
rect 6748 16658 6776 17002
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6564 15978 6592 16526
rect 6748 16250 6776 16594
rect 6840 16250 6868 16730
rect 6932 16658 6960 18176
rect 7012 18158 7064 18164
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 7024 17882 7052 18022
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 6932 16250 6960 16594
rect 7116 16522 7144 18702
rect 7366 17980 7674 17989
rect 7366 17978 7372 17980
rect 7428 17978 7452 17980
rect 7508 17978 7532 17980
rect 7588 17978 7612 17980
rect 7668 17978 7674 17980
rect 7428 17926 7430 17978
rect 7610 17926 7612 17978
rect 7366 17924 7372 17926
rect 7428 17924 7452 17926
rect 7508 17924 7532 17926
rect 7588 17924 7612 17926
rect 7668 17924 7674 17926
rect 7366 17915 7674 17924
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7300 16726 7328 17682
rect 7366 16892 7674 16901
rect 7366 16890 7372 16892
rect 7428 16890 7452 16892
rect 7508 16890 7532 16892
rect 7588 16890 7612 16892
rect 7668 16890 7674 16892
rect 7428 16838 7430 16890
rect 7610 16838 7612 16890
rect 7366 16836 7372 16838
rect 7428 16836 7452 16838
rect 7508 16836 7532 16838
rect 7588 16836 7612 16838
rect 7668 16836 7674 16838
rect 7366 16827 7674 16836
rect 8036 16726 8064 19314
rect 7288 16720 7340 16726
rect 7288 16662 7340 16668
rect 8024 16720 8076 16726
rect 8024 16662 8076 16668
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7104 16516 7156 16522
rect 7104 16458 7156 16464
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 7116 15978 7144 16458
rect 7392 16250 7420 16594
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 6552 15972 6604 15978
rect 6552 15914 6604 15920
rect 7104 15972 7156 15978
rect 7104 15914 7156 15920
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 7300 15586 7328 15846
rect 7366 15804 7674 15813
rect 7366 15802 7372 15804
rect 7428 15802 7452 15804
rect 7508 15802 7532 15804
rect 7588 15802 7612 15804
rect 7668 15802 7674 15804
rect 7428 15750 7430 15802
rect 7610 15750 7612 15802
rect 7366 15748 7372 15750
rect 7428 15748 7452 15750
rect 7508 15748 7532 15750
rect 7588 15748 7612 15750
rect 7668 15748 7674 15750
rect 7366 15739 7674 15748
rect 7300 15570 7512 15586
rect 6092 15564 6144 15570
rect 6092 15506 6144 15512
rect 6368 15564 6420 15570
rect 7300 15564 7524 15570
rect 7300 15558 7472 15564
rect 6368 15506 6420 15512
rect 7472 15506 7524 15512
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5828 14414 5856 15302
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 5632 13796 5684 13802
rect 5632 13738 5684 13744
rect 5092 13462 5120 13738
rect 5080 13456 5132 13462
rect 5080 13398 5132 13404
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4632 12442 4660 13262
rect 4724 12986 4752 13330
rect 5644 12986 5672 13738
rect 5920 13530 5948 14894
rect 6380 14890 6408 15506
rect 7484 15162 7512 15506
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 6276 14884 6328 14890
rect 6276 14826 6328 14832
rect 6368 14884 6420 14890
rect 6368 14826 6420 14832
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 6012 14074 6040 14418
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 3804 12406 4384 12434
rect 3804 11898 3832 12406
rect 4356 12374 4384 12406
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4344 12368 4396 12374
rect 4344 12310 4396 12316
rect 5448 12300 5500 12306
rect 5724 12300 5776 12306
rect 5500 12260 5724 12288
rect 5448 12242 5500 12248
rect 5724 12242 5776 12248
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 3882 11996 4190 12005
rect 3882 11994 3888 11996
rect 3944 11994 3968 11996
rect 4024 11994 4048 11996
rect 4104 11994 4128 11996
rect 4184 11994 4190 11996
rect 3944 11942 3946 11994
rect 4126 11942 4128 11994
rect 3882 11940 3888 11942
rect 3944 11940 3968 11942
rect 4024 11940 4048 11942
rect 4104 11940 4128 11942
rect 4184 11940 4190 11942
rect 3882 11931 4190 11940
rect 5828 11898 5856 12038
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5920 11694 5948 13466
rect 6104 12782 6132 14758
rect 6288 14618 6316 14826
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7366 14716 7674 14725
rect 7366 14714 7372 14716
rect 7428 14714 7452 14716
rect 7508 14714 7532 14716
rect 7588 14714 7612 14716
rect 7668 14714 7674 14716
rect 7428 14662 7430 14714
rect 7610 14662 7612 14714
rect 7366 14660 7372 14662
rect 7428 14660 7452 14662
rect 7508 14660 7532 14662
rect 7588 14660 7612 14662
rect 7668 14660 7674 14662
rect 7366 14651 7674 14660
rect 6276 14612 6328 14618
rect 6276 14554 6328 14560
rect 7760 14482 7788 14758
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7760 14074 7788 14418
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7208 12850 7236 13738
rect 7288 13728 7340 13734
rect 7288 13670 7340 13676
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7300 12782 7328 13670
rect 7366 13628 7674 13637
rect 7366 13626 7372 13628
rect 7428 13626 7452 13628
rect 7508 13626 7532 13628
rect 7588 13626 7612 13628
rect 7668 13626 7674 13628
rect 7428 13574 7430 13626
rect 7610 13574 7612 13626
rect 7366 13572 7372 13574
rect 7428 13572 7452 13574
rect 7508 13572 7532 13574
rect 7588 13572 7612 13574
rect 7668 13572 7674 13574
rect 7366 13563 7674 13572
rect 7760 13530 7788 13670
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7116 12374 7144 12582
rect 7366 12540 7674 12549
rect 7366 12538 7372 12540
rect 7428 12538 7452 12540
rect 7508 12538 7532 12540
rect 7588 12538 7612 12540
rect 7668 12538 7674 12540
rect 7428 12486 7430 12538
rect 7610 12486 7612 12538
rect 7366 12484 7372 12486
rect 7428 12484 7452 12486
rect 7508 12484 7532 12486
rect 7588 12484 7612 12486
rect 7668 12484 7674 12486
rect 7366 12475 7674 12484
rect 7760 12434 7788 12922
rect 7668 12406 7788 12434
rect 7668 12374 7696 12406
rect 7104 12368 7156 12374
rect 7104 12310 7156 12316
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 6196 11354 6224 12242
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6840 11898 6868 12038
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 3882 10908 4190 10917
rect 3882 10906 3888 10908
rect 3944 10906 3968 10908
rect 4024 10906 4048 10908
rect 4104 10906 4128 10908
rect 4184 10906 4190 10908
rect 3944 10854 3946 10906
rect 4126 10854 4128 10906
rect 3882 10852 3888 10854
rect 3944 10852 3968 10854
rect 4024 10852 4048 10854
rect 4104 10852 4128 10854
rect 4184 10852 4190 10854
rect 3882 10843 4190 10852
rect 6656 10606 6684 11630
rect 7208 11626 7236 12174
rect 7668 12170 7696 12310
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11898 8064 12038
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 8128 11694 8156 14350
rect 8220 13462 8248 19450
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8404 18290 8432 19110
rect 8680 18834 8708 19110
rect 8772 18970 8800 22066
rect 8956 22066 9260 22094
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8956 18850 8984 22066
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9048 21486 9076 21830
rect 9324 21690 9352 21830
rect 9312 21684 9364 21690
rect 9312 21626 9364 21632
rect 9324 21554 9352 21626
rect 9312 21548 9364 21554
rect 9312 21490 9364 21496
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 9048 20058 9076 21422
rect 9508 21146 9536 23122
rect 9876 22778 9904 24890
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 9680 22568 9732 22574
rect 9680 22510 9732 22516
rect 9692 22166 9720 22510
rect 9680 22160 9732 22166
rect 9680 22102 9732 22108
rect 9588 22092 9640 22098
rect 9588 22034 9640 22040
rect 9600 21690 9628 22034
rect 9588 21684 9640 21690
rect 9588 21626 9640 21632
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9496 21140 9548 21146
rect 9496 21082 9548 21088
rect 9600 20466 9628 21286
rect 9692 21078 9720 22102
rect 9968 21962 9996 27474
rect 11164 27402 11192 27950
rect 11244 27532 11296 27538
rect 11244 27474 11296 27480
rect 13268 27532 13320 27538
rect 13268 27474 13320 27480
rect 11152 27396 11204 27402
rect 11152 27338 11204 27344
rect 10692 27328 10744 27334
rect 10692 27270 10744 27276
rect 10704 27130 10732 27270
rect 10851 27228 11159 27237
rect 10851 27226 10857 27228
rect 10913 27226 10937 27228
rect 10993 27226 11017 27228
rect 11073 27226 11097 27228
rect 11153 27226 11159 27228
rect 10913 27174 10915 27226
rect 11095 27174 11097 27226
rect 10851 27172 10857 27174
rect 10913 27172 10937 27174
rect 10993 27172 11017 27174
rect 11073 27172 11097 27174
rect 11153 27172 11159 27174
rect 10851 27163 11159 27172
rect 10692 27124 10744 27130
rect 10692 27066 10744 27072
rect 11152 26988 11204 26994
rect 11152 26930 11204 26936
rect 11164 26586 11192 26930
rect 11152 26580 11204 26586
rect 11152 26522 11204 26528
rect 10048 26444 10100 26450
rect 10048 26386 10100 26392
rect 10060 22982 10088 26386
rect 10851 26140 11159 26149
rect 10851 26138 10857 26140
rect 10913 26138 10937 26140
rect 10993 26138 11017 26140
rect 11073 26138 11097 26140
rect 11153 26138 11159 26140
rect 10913 26086 10915 26138
rect 11095 26086 11097 26138
rect 10851 26084 10857 26086
rect 10913 26084 10937 26086
rect 10993 26084 11017 26086
rect 11073 26084 11097 26086
rect 11153 26084 11159 26086
rect 10851 26075 11159 26084
rect 10851 25052 11159 25061
rect 10851 25050 10857 25052
rect 10913 25050 10937 25052
rect 10993 25050 11017 25052
rect 11073 25050 11097 25052
rect 11153 25050 11159 25052
rect 10913 24998 10915 25050
rect 11095 24998 11097 25050
rect 10851 24996 10857 24998
rect 10913 24996 10937 24998
rect 10993 24996 11017 24998
rect 11073 24996 11097 24998
rect 11153 24996 11159 24998
rect 10851 24987 11159 24996
rect 11060 24744 11112 24750
rect 11060 24686 11112 24692
rect 10600 24676 10652 24682
rect 10600 24618 10652 24624
rect 10784 24676 10836 24682
rect 10784 24618 10836 24624
rect 10416 24608 10468 24614
rect 10416 24550 10468 24556
rect 10428 24410 10456 24550
rect 10612 24410 10640 24618
rect 10796 24410 10824 24618
rect 10968 24608 11020 24614
rect 10968 24550 11020 24556
rect 10416 24404 10468 24410
rect 10416 24346 10468 24352
rect 10600 24404 10652 24410
rect 10600 24346 10652 24352
rect 10784 24404 10836 24410
rect 10784 24346 10836 24352
rect 10980 24206 11008 24550
rect 11072 24206 11100 24686
rect 11152 24404 11204 24410
rect 11152 24346 11204 24352
rect 11164 24206 11192 24346
rect 10968 24200 11020 24206
rect 10968 24142 11020 24148
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 11152 24200 11204 24206
rect 11152 24142 11204 24148
rect 10692 24064 10744 24070
rect 10692 24006 10744 24012
rect 10704 23322 10732 24006
rect 10851 23964 11159 23973
rect 10851 23962 10857 23964
rect 10913 23962 10937 23964
rect 10993 23962 11017 23964
rect 11073 23962 11097 23964
rect 11153 23962 11159 23964
rect 10913 23910 10915 23962
rect 11095 23910 11097 23962
rect 10851 23908 10857 23910
rect 10913 23908 10937 23910
rect 10993 23908 11017 23910
rect 11073 23908 11097 23910
rect 11153 23908 11159 23910
rect 10851 23899 11159 23908
rect 10692 23316 10744 23322
rect 10692 23258 10744 23264
rect 10048 22976 10100 22982
rect 10048 22918 10100 22924
rect 10692 22976 10744 22982
rect 10692 22918 10744 22924
rect 10416 22772 10468 22778
rect 10416 22714 10468 22720
rect 9956 21956 10008 21962
rect 9956 21898 10008 21904
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9876 21554 9904 21830
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9680 21072 9732 21078
rect 9680 21014 9732 21020
rect 9588 20460 9640 20466
rect 9588 20402 9640 20408
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 9324 20058 9352 20334
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 9312 20052 9364 20058
rect 9312 19994 9364 20000
rect 9600 19446 9628 20402
rect 9784 19922 9812 21082
rect 10060 20942 10088 21422
rect 10232 21412 10284 21418
rect 10232 21354 10284 21360
rect 10244 21010 10272 21354
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 10336 21146 10364 21286
rect 10324 21140 10376 21146
rect 10324 21082 10376 21088
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 9864 20936 9916 20942
rect 9862 20904 9864 20913
rect 9956 20936 10008 20942
rect 9916 20904 9918 20913
rect 9956 20878 10008 20884
rect 10048 20936 10100 20942
rect 10048 20878 10100 20884
rect 9862 20839 9918 20848
rect 9968 20602 9996 20878
rect 9956 20596 10008 20602
rect 10008 20556 10088 20584
rect 9956 20538 10008 20544
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9956 19916 10008 19922
rect 9956 19858 10008 19864
rect 9968 19446 9996 19858
rect 10060 19446 10088 20556
rect 10244 19718 10272 20946
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 9588 19440 9640 19446
rect 9588 19382 9640 19388
rect 9956 19440 10008 19446
rect 9956 19382 10008 19388
rect 10048 19440 10100 19446
rect 10048 19382 10100 19388
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 9048 18902 9076 19110
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8864 18822 8984 18850
rect 9036 18896 9088 18902
rect 9036 18838 9088 18844
rect 8680 18426 8708 18770
rect 8864 18698 8892 18822
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8944 18692 8996 18698
rect 8944 18634 8996 18640
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8496 17746 8524 18022
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 8312 16794 8340 17682
rect 8680 17354 8708 18362
rect 8772 17542 8800 18566
rect 8852 18216 8904 18222
rect 8852 18158 8904 18164
rect 8864 17610 8892 18158
rect 8956 18086 8984 18634
rect 9048 18426 9076 18838
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9600 18222 9628 18770
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 8944 18080 8996 18086
rect 8944 18022 8996 18028
rect 8852 17604 8904 17610
rect 8852 17546 8904 17552
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8680 17326 8800 17354
rect 8956 17338 8984 18022
rect 9600 17610 9628 18158
rect 9692 17882 9720 18158
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9588 17604 9640 17610
rect 9588 17546 9640 17552
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8588 16046 8616 16934
rect 8680 16522 8708 16934
rect 8668 16516 8720 16522
rect 8668 16458 8720 16464
rect 8680 16182 8708 16458
rect 8668 16176 8720 16182
rect 8668 16118 8720 16124
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8680 15502 8708 16118
rect 8772 15978 8800 17326
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 9784 17082 9812 19246
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9876 17338 9904 18022
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9692 17054 9812 17082
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 8956 16658 8984 16934
rect 9692 16726 9720 17054
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9784 16794 9812 16934
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9680 16720 9732 16726
rect 9680 16662 9732 16668
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 8956 16046 8984 16594
rect 9600 16250 9628 16594
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8588 15162 8616 15438
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8680 14482 8708 15438
rect 8772 14822 8800 15914
rect 8956 15026 8984 15982
rect 9692 15434 9720 16662
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 8944 15020 8996 15026
rect 9692 15008 9720 15370
rect 9772 15020 9824 15026
rect 9692 14980 9772 15008
rect 8944 14962 8996 14968
rect 9772 14962 9824 14968
rect 9588 14952 9640 14958
rect 9640 14900 9812 14906
rect 9588 14894 9812 14900
rect 9600 14878 9812 14894
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8772 12850 8800 14758
rect 8956 14414 8984 14758
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 8956 14074 8984 14350
rect 9692 14346 9720 14758
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8680 12374 8708 12718
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6748 11218 6776 11494
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 7024 10810 7052 11494
rect 7366 11452 7674 11461
rect 7366 11450 7372 11452
rect 7428 11450 7452 11452
rect 7508 11450 7532 11452
rect 7588 11450 7612 11452
rect 7668 11450 7674 11452
rect 7428 11398 7430 11450
rect 7610 11398 7612 11450
rect 7366 11396 7372 11398
rect 7428 11396 7452 11398
rect 7508 11396 7532 11398
rect 7588 11396 7612 11398
rect 7668 11396 7674 11398
rect 7366 11387 7674 11396
rect 8772 11218 8800 12786
rect 8956 12782 8984 14010
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9048 12986 9076 13262
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8956 12102 8984 12718
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9232 11354 9260 11494
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 8956 11234 8984 11290
rect 9128 11280 9180 11286
rect 8956 11228 9128 11234
rect 8956 11222 9180 11228
rect 8760 11212 8812 11218
rect 8956 11206 9168 11222
rect 8760 11154 8812 11160
rect 9324 11150 9352 11834
rect 9416 11762 9444 13262
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9600 11830 9628 12038
rect 9692 11898 9720 13126
rect 9784 12986 9812 14878
rect 9876 14618 9904 15846
rect 9968 14958 9996 19246
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 10060 17338 10088 17682
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 10336 16794 10364 19654
rect 10428 17066 10456 22714
rect 10704 22574 10732 22918
rect 10851 22876 11159 22885
rect 10851 22874 10857 22876
rect 10913 22874 10937 22876
rect 10993 22874 11017 22876
rect 11073 22874 11097 22876
rect 11153 22874 11159 22876
rect 10913 22822 10915 22874
rect 11095 22822 11097 22874
rect 10851 22820 10857 22822
rect 10913 22820 10937 22822
rect 10993 22820 11017 22822
rect 11073 22820 11097 22822
rect 11153 22820 11159 22822
rect 10851 22811 11159 22820
rect 10692 22568 10744 22574
rect 10692 22510 10744 22516
rect 10600 22160 10652 22166
rect 10652 22108 11100 22114
rect 10600 22102 11100 22108
rect 10612 22098 11100 22102
rect 10508 22092 10560 22098
rect 10612 22092 11112 22098
rect 11256 22094 11284 27474
rect 13280 27130 13308 27474
rect 13464 27334 13492 28600
rect 14335 27772 14643 27781
rect 14335 27770 14341 27772
rect 14397 27770 14421 27772
rect 14477 27770 14501 27772
rect 14557 27770 14581 27772
rect 14637 27770 14643 27772
rect 14397 27718 14399 27770
rect 14579 27718 14581 27770
rect 14335 27716 14341 27718
rect 14397 27716 14421 27718
rect 14477 27716 14501 27718
rect 14557 27716 14581 27718
rect 14637 27716 14643 27718
rect 14335 27707 14643 27716
rect 15488 27606 15516 28600
rect 17512 28014 17540 28600
rect 17820 28316 18128 28325
rect 17820 28314 17826 28316
rect 17882 28314 17906 28316
rect 17962 28314 17986 28316
rect 18042 28314 18066 28316
rect 18122 28314 18128 28316
rect 17882 28262 17884 28314
rect 18064 28262 18066 28314
rect 17820 28260 17826 28262
rect 17882 28260 17906 28262
rect 17962 28260 17986 28262
rect 18042 28260 18066 28262
rect 18122 28260 18128 28262
rect 17820 28251 18128 28260
rect 19536 28218 19564 28600
rect 19524 28212 19576 28218
rect 19524 28154 19576 28160
rect 21560 28014 21588 28600
rect 23584 28014 23612 28600
rect 24789 28316 25097 28325
rect 24789 28314 24795 28316
rect 24851 28314 24875 28316
rect 24931 28314 24955 28316
rect 25011 28314 25035 28316
rect 25091 28314 25097 28316
rect 24851 28262 24853 28314
rect 25033 28262 25035 28314
rect 24789 28260 24795 28262
rect 24851 28260 24875 28262
rect 24931 28260 24955 28262
rect 25011 28260 25035 28262
rect 25091 28260 25097 28262
rect 24789 28251 25097 28260
rect 25608 28014 25636 28600
rect 15660 28008 15712 28014
rect 15660 27950 15712 27956
rect 17500 28008 17552 28014
rect 17500 27950 17552 27956
rect 19248 28008 19300 28014
rect 19248 27950 19300 27956
rect 21548 28008 21600 28014
rect 21548 27950 21600 27956
rect 23572 28008 23624 28014
rect 23572 27950 23624 27956
rect 25596 28008 25648 28014
rect 25596 27950 25648 27956
rect 15672 27674 15700 27950
rect 16212 27872 16264 27878
rect 16212 27814 16264 27820
rect 18144 27872 18196 27878
rect 18144 27814 18196 27820
rect 15660 27668 15712 27674
rect 15660 27610 15712 27616
rect 15016 27600 15068 27606
rect 15016 27542 15068 27548
rect 15476 27600 15528 27606
rect 15476 27542 15528 27548
rect 14188 27396 14240 27402
rect 14188 27338 14240 27344
rect 13452 27328 13504 27334
rect 13452 27270 13504 27276
rect 13268 27124 13320 27130
rect 13268 27066 13320 27072
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 12808 26920 12860 26926
rect 12808 26862 12860 26868
rect 11428 26784 11480 26790
rect 11428 26726 11480 26732
rect 11980 26784 12032 26790
rect 11980 26726 12032 26732
rect 11336 25968 11388 25974
rect 11336 25910 11388 25916
rect 11348 23322 11376 25910
rect 11336 23316 11388 23322
rect 11336 23258 11388 23264
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 10612 22086 11060 22092
rect 10508 22034 10560 22040
rect 11060 22034 11112 22040
rect 11164 22066 11284 22094
rect 11348 22094 11376 23054
rect 11440 22778 11468 26726
rect 11992 26586 12020 26726
rect 11980 26580 12032 26586
rect 11980 26522 12032 26528
rect 12256 26444 12308 26450
rect 12256 26386 12308 26392
rect 12348 26444 12400 26450
rect 12348 26386 12400 26392
rect 11612 26308 11664 26314
rect 11612 26250 11664 26256
rect 11796 26308 11848 26314
rect 11796 26250 11848 26256
rect 11624 25430 11652 26250
rect 11612 25424 11664 25430
rect 11612 25366 11664 25372
rect 11624 24274 11652 25366
rect 11704 24880 11756 24886
rect 11704 24822 11756 24828
rect 11716 24614 11744 24822
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11612 24268 11664 24274
rect 11612 24210 11664 24216
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11532 22094 11560 23802
rect 11624 23526 11652 24210
rect 11716 24138 11744 24550
rect 11808 24274 11836 26250
rect 12268 25838 12296 26386
rect 12256 25832 12308 25838
rect 12256 25774 12308 25780
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 11900 24954 11928 25638
rect 12268 25498 12296 25774
rect 12256 25492 12308 25498
rect 12256 25434 12308 25440
rect 11888 24948 11940 24954
rect 11888 24890 11940 24896
rect 12360 24818 12388 26386
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 11796 24268 11848 24274
rect 11796 24210 11848 24216
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 11704 24132 11756 24138
rect 11704 24074 11756 24080
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11612 23520 11664 23526
rect 11612 23462 11664 23468
rect 11808 23186 11836 24006
rect 11888 23316 11940 23322
rect 11888 23258 11940 23264
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 11704 23112 11756 23118
rect 11704 23054 11756 23060
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 11624 22710 11652 22918
rect 11612 22704 11664 22710
rect 11612 22646 11664 22652
rect 11716 22506 11744 23054
rect 11808 22778 11836 23122
rect 11900 22778 11928 23258
rect 11796 22772 11848 22778
rect 11796 22714 11848 22720
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 11704 22500 11756 22506
rect 11704 22442 11756 22448
rect 11348 22066 11468 22094
rect 11532 22066 11652 22094
rect 10520 21486 10548 22034
rect 11164 21962 11192 22066
rect 11152 21956 11204 21962
rect 11152 21898 11204 21904
rect 11440 21894 11468 22066
rect 11428 21888 11480 21894
rect 11428 21830 11480 21836
rect 10851 21788 11159 21797
rect 10851 21786 10857 21788
rect 10913 21786 10937 21788
rect 10993 21786 11017 21788
rect 11073 21786 11097 21788
rect 11153 21786 11159 21788
rect 10913 21734 10915 21786
rect 11095 21734 11097 21786
rect 10851 21732 10857 21734
rect 10913 21732 10937 21734
rect 10993 21732 11017 21734
rect 11073 21732 11097 21734
rect 11153 21732 11159 21734
rect 10851 21723 11159 21732
rect 10508 21480 10560 21486
rect 10508 21422 10560 21428
rect 11244 20868 11296 20874
rect 11244 20810 11296 20816
rect 10851 20700 11159 20709
rect 10851 20698 10857 20700
rect 10913 20698 10937 20700
rect 10993 20698 11017 20700
rect 11073 20698 11097 20700
rect 11153 20698 11159 20700
rect 10913 20646 10915 20698
rect 11095 20646 11097 20698
rect 10851 20644 10857 20646
rect 10913 20644 10937 20646
rect 10993 20644 11017 20646
rect 11073 20644 11097 20646
rect 11153 20644 11159 20646
rect 10851 20635 11159 20644
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11072 20505 11100 20538
rect 11058 20496 11114 20505
rect 11058 20431 11114 20440
rect 11256 20398 11284 20810
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 11440 20330 11468 21830
rect 11624 21570 11652 22066
rect 11532 21542 11652 21570
rect 11532 21078 11560 21542
rect 11610 21448 11666 21457
rect 11610 21383 11666 21392
rect 11520 21072 11572 21078
rect 11520 21014 11572 21020
rect 11428 20324 11480 20330
rect 11428 20266 11480 20272
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 11348 20058 11376 20198
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 10851 19612 11159 19621
rect 10851 19610 10857 19612
rect 10913 19610 10937 19612
rect 10993 19610 11017 19612
rect 11073 19610 11097 19612
rect 11153 19610 11159 19612
rect 10913 19558 10915 19610
rect 11095 19558 11097 19610
rect 10851 19556 10857 19558
rect 10913 19556 10937 19558
rect 10993 19556 11017 19558
rect 11073 19556 11097 19558
rect 11153 19556 11159 19558
rect 10851 19547 11159 19556
rect 11256 19378 11284 19654
rect 11244 19372 11296 19378
rect 11244 19314 11296 19320
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10980 18834 11008 19110
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10851 18524 11159 18533
rect 10851 18522 10857 18524
rect 10913 18522 10937 18524
rect 10993 18522 11017 18524
rect 11073 18522 11097 18524
rect 11153 18522 11159 18524
rect 10913 18470 10915 18522
rect 11095 18470 11097 18522
rect 10851 18468 10857 18470
rect 10913 18468 10937 18470
rect 10993 18468 11017 18470
rect 11073 18468 11097 18470
rect 11153 18468 11159 18470
rect 10851 18459 11159 18468
rect 11532 18426 11560 21014
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 10851 17436 11159 17445
rect 10851 17434 10857 17436
rect 10913 17434 10937 17436
rect 10993 17434 11017 17436
rect 11073 17434 11097 17436
rect 11153 17434 11159 17436
rect 10913 17382 10915 17434
rect 11095 17382 11097 17434
rect 10851 17380 10857 17382
rect 10913 17380 10937 17382
rect 10993 17380 11017 17382
rect 11073 17380 11097 17382
rect 11153 17380 11159 17382
rect 10851 17371 11159 17380
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 11256 16658 11284 17614
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11532 16794 11560 17478
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10704 16046 10732 16390
rect 10851 16348 11159 16357
rect 10851 16346 10857 16348
rect 10913 16346 10937 16348
rect 10993 16346 11017 16348
rect 11073 16346 11097 16348
rect 11153 16346 11159 16348
rect 10913 16294 10915 16346
rect 11095 16294 11097 16346
rect 10851 16292 10857 16294
rect 10913 16292 10937 16294
rect 10993 16292 11017 16294
rect 11073 16292 11097 16294
rect 11153 16292 11159 16294
rect 10851 16283 11159 16292
rect 11256 16046 11284 16594
rect 11624 16046 11652 21383
rect 11716 20942 11744 22442
rect 11980 21956 12032 21962
rect 11980 21898 12032 21904
rect 11888 21616 11940 21622
rect 11888 21558 11940 21564
rect 11900 21457 11928 21558
rect 11886 21448 11942 21457
rect 11886 21383 11942 21392
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11704 20936 11756 20942
rect 11704 20878 11756 20884
rect 11808 18970 11836 21286
rect 11992 21078 12020 21898
rect 12084 21554 12112 24142
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 12268 23186 12296 23462
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 12256 23180 12308 23186
rect 12256 23122 12308 23128
rect 12348 23180 12400 23186
rect 12348 23122 12400 23128
rect 12176 22778 12204 23122
rect 12164 22772 12216 22778
rect 12164 22714 12216 22720
rect 12268 22166 12296 23122
rect 12360 22953 12388 23122
rect 12346 22944 12402 22953
rect 12346 22879 12402 22888
rect 12256 22160 12308 22166
rect 12256 22102 12308 22108
rect 12452 22030 12480 26862
rect 12624 26784 12676 26790
rect 12624 26726 12676 26732
rect 12636 26450 12664 26726
rect 12820 26586 12848 26862
rect 13912 26784 13964 26790
rect 13912 26726 13964 26732
rect 12808 26580 12860 26586
rect 12808 26522 12860 26528
rect 13924 26518 13952 26726
rect 14200 26586 14228 27338
rect 14832 27328 14884 27334
rect 14832 27270 14884 27276
rect 14740 26920 14792 26926
rect 14740 26862 14792 26868
rect 14335 26684 14643 26693
rect 14335 26682 14341 26684
rect 14397 26682 14421 26684
rect 14477 26682 14501 26684
rect 14557 26682 14581 26684
rect 14637 26682 14643 26684
rect 14397 26630 14399 26682
rect 14579 26630 14581 26682
rect 14335 26628 14341 26630
rect 14397 26628 14421 26630
rect 14477 26628 14501 26630
rect 14557 26628 14581 26630
rect 14637 26628 14643 26630
rect 14335 26619 14643 26628
rect 14752 26586 14780 26862
rect 14188 26580 14240 26586
rect 14188 26522 14240 26528
rect 14740 26580 14792 26586
rect 14740 26522 14792 26528
rect 13912 26512 13964 26518
rect 13912 26454 13964 26460
rect 12532 26444 12584 26450
rect 12532 26386 12584 26392
rect 12624 26444 12676 26450
rect 12624 26386 12676 26392
rect 12544 26042 12572 26386
rect 13084 26308 13136 26314
rect 13084 26250 13136 26256
rect 13096 26042 13124 26250
rect 12532 26036 12584 26042
rect 12532 25978 12584 25984
rect 13084 26036 13136 26042
rect 13084 25978 13136 25984
rect 13924 25974 13952 26454
rect 14004 26240 14056 26246
rect 14004 26182 14056 26188
rect 13912 25968 13964 25974
rect 13912 25910 13964 25916
rect 14016 25838 14044 26182
rect 14004 25832 14056 25838
rect 14004 25774 14056 25780
rect 12624 25764 12676 25770
rect 12624 25706 12676 25712
rect 12716 25764 12768 25770
rect 12716 25706 12768 25712
rect 12532 25288 12584 25294
rect 12532 25230 12584 25236
rect 12544 24954 12572 25230
rect 12532 24948 12584 24954
rect 12532 24890 12584 24896
rect 12636 24750 12664 25706
rect 12728 25158 12756 25706
rect 14200 25480 14228 26522
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 14335 25596 14643 25605
rect 14335 25594 14341 25596
rect 14397 25594 14421 25596
rect 14477 25594 14501 25596
rect 14557 25594 14581 25596
rect 14637 25594 14643 25596
rect 14397 25542 14399 25594
rect 14579 25542 14581 25594
rect 14335 25540 14341 25542
rect 14397 25540 14421 25542
rect 14477 25540 14501 25542
rect 14557 25540 14581 25542
rect 14637 25540 14643 25542
rect 14335 25531 14643 25540
rect 14372 25492 14424 25498
rect 14200 25452 14372 25480
rect 14004 25424 14056 25430
rect 13726 25392 13782 25401
rect 14004 25366 14056 25372
rect 13726 25327 13728 25336
rect 13780 25327 13782 25336
rect 13728 25298 13780 25304
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 13084 25152 13136 25158
rect 13084 25094 13136 25100
rect 12728 24750 12756 25094
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12716 24744 12768 24750
rect 12716 24686 12768 24692
rect 12728 23866 12756 24686
rect 12992 24404 13044 24410
rect 12992 24346 13044 24352
rect 12808 24200 12860 24206
rect 12808 24142 12860 24148
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12532 23520 12584 23526
rect 12532 23462 12584 23468
rect 12544 23186 12572 23462
rect 12532 23180 12584 23186
rect 12532 23122 12584 23128
rect 12624 23044 12676 23050
rect 12624 22986 12676 22992
rect 12636 22778 12664 22986
rect 12624 22772 12676 22778
rect 12624 22714 12676 22720
rect 12728 22642 12756 23802
rect 12820 23594 12848 24142
rect 13004 23730 13032 24346
rect 13096 24274 13124 25094
rect 14016 24750 14044 25366
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 13912 24744 13964 24750
rect 13912 24686 13964 24692
rect 14004 24744 14056 24750
rect 14004 24686 14056 24692
rect 13924 24410 13952 24686
rect 14016 24410 14044 24686
rect 14108 24682 14136 25094
rect 14200 24954 14228 25452
rect 14372 25434 14424 25440
rect 14556 25288 14608 25294
rect 14556 25230 14608 25236
rect 14188 24948 14240 24954
rect 14188 24890 14240 24896
rect 14568 24682 14596 25230
rect 14752 24954 14780 26318
rect 14844 25906 14872 27270
rect 15028 27130 15056 27542
rect 16224 27538 16252 27814
rect 15200 27532 15252 27538
rect 15200 27474 15252 27480
rect 16212 27532 16264 27538
rect 16212 27474 16264 27480
rect 15108 27328 15160 27334
rect 15108 27270 15160 27276
rect 15016 27124 15068 27130
rect 15016 27066 15068 27072
rect 15120 26790 15148 27270
rect 15212 26994 15240 27474
rect 16120 27464 16172 27470
rect 16120 27406 16172 27412
rect 15200 26988 15252 26994
rect 15200 26930 15252 26936
rect 15292 26920 15344 26926
rect 15292 26862 15344 26868
rect 15108 26784 15160 26790
rect 15108 26726 15160 26732
rect 15304 26586 15332 26862
rect 15292 26580 15344 26586
rect 15292 26522 15344 26528
rect 16132 26450 16160 27406
rect 17820 27228 18128 27237
rect 17820 27226 17826 27228
rect 17882 27226 17906 27228
rect 17962 27226 17986 27228
rect 18042 27226 18066 27228
rect 18122 27226 18128 27228
rect 17882 27174 17884 27226
rect 18064 27174 18066 27226
rect 17820 27172 17826 27174
rect 17882 27172 17906 27174
rect 17962 27172 17986 27174
rect 18042 27172 18066 27174
rect 18122 27172 18128 27174
rect 17820 27163 18128 27172
rect 16764 27056 16816 27062
rect 16764 26998 16816 27004
rect 16672 26920 16724 26926
rect 16672 26862 16724 26868
rect 16120 26444 16172 26450
rect 16120 26386 16172 26392
rect 16580 26444 16632 26450
rect 16580 26386 16632 26392
rect 15200 26376 15252 26382
rect 15200 26318 15252 26324
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 14924 25832 14976 25838
rect 14924 25774 14976 25780
rect 14832 25492 14884 25498
rect 14832 25434 14884 25440
rect 14740 24948 14792 24954
rect 14740 24890 14792 24896
rect 14096 24676 14148 24682
rect 14096 24618 14148 24624
rect 14556 24676 14608 24682
rect 14556 24618 14608 24624
rect 13912 24404 13964 24410
rect 13912 24346 13964 24352
rect 14004 24404 14056 24410
rect 14004 24346 14056 24352
rect 13084 24268 13136 24274
rect 13084 24210 13136 24216
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 13096 23662 13124 24210
rect 14108 24206 14136 24618
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 14200 24410 14228 24550
rect 14335 24508 14643 24517
rect 14335 24506 14341 24508
rect 14397 24506 14421 24508
rect 14477 24506 14501 24508
rect 14557 24506 14581 24508
rect 14637 24506 14643 24508
rect 14397 24454 14399 24506
rect 14579 24454 14581 24506
rect 14335 24452 14341 24454
rect 14397 24452 14421 24454
rect 14477 24452 14501 24454
rect 14557 24452 14581 24454
rect 14637 24452 14643 24454
rect 14335 24443 14643 24452
rect 14188 24404 14240 24410
rect 14188 24346 14240 24352
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 14648 24064 14700 24070
rect 14752 24052 14780 24890
rect 14844 24886 14872 25434
rect 14936 25294 14964 25774
rect 14924 25288 14976 25294
rect 14924 25230 14976 25236
rect 14832 24880 14884 24886
rect 14832 24822 14884 24828
rect 14700 24024 14780 24052
rect 14648 24006 14700 24012
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 13084 23656 13136 23662
rect 13084 23598 13136 23604
rect 12808 23588 12860 23594
rect 12808 23530 12860 23536
rect 12992 23588 13044 23594
rect 12992 23530 13044 23536
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12820 22574 12848 23530
rect 13004 23322 13032 23530
rect 12992 23316 13044 23322
rect 12992 23258 13044 23264
rect 13096 23186 13124 23598
rect 13636 23520 13688 23526
rect 13636 23462 13688 23468
rect 12900 23180 12952 23186
rect 12900 23122 12952 23128
rect 13084 23180 13136 23186
rect 13084 23122 13136 23128
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 12808 22568 12860 22574
rect 12808 22510 12860 22516
rect 12912 22438 12940 23122
rect 13174 23080 13230 23089
rect 13174 23015 13176 23024
rect 13228 23015 13230 23024
rect 13176 22986 13228 22992
rect 13372 22506 13400 23122
rect 13648 22982 13676 23462
rect 13832 23322 13860 23666
rect 13820 23316 13872 23322
rect 13820 23258 13872 23264
rect 13726 23080 13782 23089
rect 13726 23015 13782 23024
rect 13740 22982 13768 23015
rect 13636 22976 13688 22982
rect 13636 22918 13688 22924
rect 13728 22976 13780 22982
rect 13728 22918 13780 22924
rect 13648 22710 13676 22918
rect 13636 22704 13688 22710
rect 13636 22646 13688 22652
rect 13360 22500 13412 22506
rect 13360 22442 13412 22448
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 12900 22432 12952 22438
rect 12900 22374 12952 22380
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 12544 21146 12572 22374
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12532 21140 12584 21146
rect 12532 21082 12584 21088
rect 11980 21072 12032 21078
rect 11900 21032 11980 21060
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11900 16114 11928 21032
rect 11980 21014 12032 21020
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 11992 20398 12020 20878
rect 11980 20392 12032 20398
rect 11980 20334 12032 20340
rect 11992 20058 12020 20334
rect 12164 20324 12216 20330
rect 12164 20266 12216 20272
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11980 19236 12032 19242
rect 11980 19178 12032 19184
rect 11992 18970 12020 19178
rect 12176 18986 12204 20266
rect 12348 20256 12400 20262
rect 12348 20198 12400 20204
rect 12360 19334 12388 20198
rect 12544 19718 12572 21082
rect 12636 20466 12664 21966
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12728 20534 12756 21422
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 12820 20602 12848 20946
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 12716 20528 12768 20534
rect 12716 20470 12768 20476
rect 12624 20460 12676 20466
rect 12624 20402 12676 20408
rect 12912 20262 12940 22374
rect 13372 22166 13400 22442
rect 13360 22160 13412 22166
rect 13636 22160 13688 22166
rect 13360 22102 13412 22108
rect 13556 22120 13636 22148
rect 13556 21146 13584 22120
rect 13636 22102 13688 22108
rect 13740 22001 13768 22918
rect 13924 22094 13952 24006
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 14108 23322 14136 23802
rect 14188 23520 14240 23526
rect 14188 23462 14240 23468
rect 14004 23316 14056 23322
rect 14004 23258 14056 23264
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 14016 23050 14044 23258
rect 14004 23044 14056 23050
rect 14004 22986 14056 22992
rect 14016 22710 14044 22986
rect 14200 22794 14228 23462
rect 14335 23420 14643 23429
rect 14335 23418 14341 23420
rect 14397 23418 14421 23420
rect 14477 23418 14501 23420
rect 14557 23418 14581 23420
rect 14637 23418 14643 23420
rect 14397 23366 14399 23418
rect 14579 23366 14581 23418
rect 14335 23364 14341 23366
rect 14397 23364 14421 23366
rect 14477 23364 14501 23366
rect 14557 23364 14581 23366
rect 14637 23364 14643 23366
rect 14335 23355 14643 23364
rect 14832 23180 14884 23186
rect 14832 23122 14884 23128
rect 14740 23112 14792 23118
rect 14740 23054 14792 23060
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14108 22766 14228 22794
rect 14004 22704 14056 22710
rect 14004 22646 14056 22652
rect 13924 22066 14044 22094
rect 13726 21992 13782 22001
rect 13726 21927 13782 21936
rect 14016 21690 14044 22066
rect 14004 21684 14056 21690
rect 14004 21626 14056 21632
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 12992 20392 13044 20398
rect 12992 20334 13044 20340
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 13004 20058 13032 20334
rect 13188 20262 13216 20334
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 12992 20052 13044 20058
rect 13188 20040 13216 20198
rect 13556 20058 13584 21082
rect 13912 21072 13964 21078
rect 13912 21014 13964 21020
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 13648 20058 13676 20334
rect 12992 19994 13044 20000
rect 13096 20012 13216 20040
rect 13268 20052 13320 20058
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12820 19378 12848 19858
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 12808 19372 12860 19378
rect 12360 19306 12664 19334
rect 12808 19314 12860 19320
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 12084 18958 12204 18986
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11612 16040 11664 16046
rect 11664 15988 11836 15994
rect 11612 15982 11836 15988
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10704 15094 10732 15370
rect 10851 15260 11159 15269
rect 10851 15258 10857 15260
rect 10913 15258 10937 15260
rect 10993 15258 11017 15260
rect 11073 15258 11097 15260
rect 11153 15258 11159 15260
rect 10913 15206 10915 15258
rect 11095 15206 11097 15258
rect 10851 15204 10857 15206
rect 10913 15204 10937 15206
rect 10993 15204 11017 15206
rect 11073 15204 11097 15206
rect 11153 15204 11159 15206
rect 10851 15195 11159 15204
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 10322 14920 10378 14929
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9876 13870 9904 14554
rect 9968 14414 9996 14894
rect 10322 14855 10378 14864
rect 10336 14822 10364 14855
rect 10324 14816 10376 14822
rect 10600 14816 10652 14822
rect 10376 14776 10456 14804
rect 10324 14758 10376 14764
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 10152 13394 10180 14282
rect 10428 13530 10456 14776
rect 10600 14758 10652 14764
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10612 14618 10640 14758
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10704 14550 10732 14758
rect 10692 14544 10744 14550
rect 10692 14486 10744 14492
rect 11256 14278 11284 15982
rect 11624 15966 11836 15982
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 11348 14618 11376 14962
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 10520 14006 10548 14214
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10704 13870 10732 14214
rect 10851 14172 11159 14181
rect 10851 14170 10857 14172
rect 10913 14170 10937 14172
rect 10993 14170 11017 14172
rect 11073 14170 11097 14172
rect 11153 14170 11159 14172
rect 10913 14118 10915 14170
rect 11095 14118 11097 14170
rect 10851 14116 10857 14118
rect 10913 14116 10937 14118
rect 10993 14116 11017 14118
rect 11073 14116 11097 14118
rect 11153 14116 11159 14118
rect 10851 14107 11159 14116
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10336 13410 10364 13466
rect 11256 13462 11284 14214
rect 11348 14074 11376 14418
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11440 13938 11468 15846
rect 11808 15026 11836 15966
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11704 14952 11756 14958
rect 11702 14920 11704 14929
rect 11756 14920 11758 14929
rect 11702 14855 11758 14864
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11428 13932 11480 13938
rect 11428 13874 11480 13880
rect 11440 13462 11468 13874
rect 11244 13456 11296 13462
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 10140 13388 10192 13394
rect 10336 13382 10456 13410
rect 11244 13398 11296 13404
rect 11428 13456 11480 13462
rect 11428 13398 11480 13404
rect 10140 13330 10192 13336
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9784 12442 9812 12718
rect 9876 12714 9904 13330
rect 10152 12850 10180 13330
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 10244 12646 10272 12718
rect 10336 12714 10364 13262
rect 10428 13190 10456 13382
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10428 12918 10456 13126
rect 10851 13084 11159 13093
rect 10851 13082 10857 13084
rect 10913 13082 10937 13084
rect 10993 13082 11017 13084
rect 11073 13082 11097 13084
rect 11153 13082 11159 13084
rect 10913 13030 10915 13082
rect 11095 13030 11097 13082
rect 10851 13028 10857 13030
rect 10913 13028 10937 13030
rect 10993 13028 11017 13030
rect 11073 13028 11097 13030
rect 11153 13028 11159 13030
rect 10851 13019 11159 13028
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9784 11626 9812 12378
rect 10520 12306 10548 12922
rect 11256 12850 11284 13398
rect 11532 13172 11560 14758
rect 11716 14550 11744 14758
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11704 13184 11756 13190
rect 11532 13144 11704 13172
rect 11704 13126 11756 13132
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 10796 12646 10824 12786
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9876 11830 9904 12106
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 9876 11694 9904 11766
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10152 11286 10180 11494
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10428 11218 10456 11494
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 7392 10538 7420 10950
rect 7380 10532 7432 10538
rect 7380 10474 7432 10480
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7366 10364 7674 10373
rect 7366 10362 7372 10364
rect 7428 10362 7452 10364
rect 7508 10362 7532 10364
rect 7588 10362 7612 10364
rect 7668 10362 7674 10364
rect 7428 10310 7430 10362
rect 7610 10310 7612 10362
rect 7366 10308 7372 10310
rect 7428 10308 7452 10310
rect 7508 10308 7532 10310
rect 7588 10308 7612 10310
rect 7668 10308 7674 10310
rect 7366 10299 7674 10308
rect 7852 10130 7880 10406
rect 8220 10198 8248 11086
rect 10520 11082 10548 12242
rect 10612 11898 10640 12582
rect 10851 11996 11159 12005
rect 10851 11994 10857 11996
rect 10913 11994 10937 11996
rect 10993 11994 11017 11996
rect 11073 11994 11097 11996
rect 11153 11994 11159 11996
rect 10913 11942 10915 11994
rect 11095 11942 11097 11994
rect 10851 11940 10857 11942
rect 10913 11940 10937 11942
rect 10993 11940 11017 11942
rect 11073 11940 11097 11942
rect 11153 11940 11159 11942
rect 10851 11931 11159 11940
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 11256 11150 11284 12786
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11532 11898 11560 12038
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 9232 10266 9260 11018
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10152 10538 10180 10950
rect 10851 10908 11159 10917
rect 10851 10906 10857 10908
rect 10913 10906 10937 10908
rect 10993 10906 11017 10908
rect 11073 10906 11097 10908
rect 11153 10906 11159 10908
rect 10913 10854 10915 10906
rect 11095 10854 11097 10906
rect 10851 10852 10857 10854
rect 10913 10852 10937 10854
rect 10993 10852 11017 10854
rect 11073 10852 11097 10854
rect 11153 10852 11159 10854
rect 10851 10843 11159 10852
rect 11256 10606 11284 11086
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11348 10810 11376 11018
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11624 10674 11652 11494
rect 11716 11354 11744 13126
rect 11900 12986 11928 16050
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11992 14958 12020 15302
rect 12084 15162 12112 18958
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12176 18426 12204 18770
rect 12636 18630 12664 19306
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12452 17678 12480 18158
rect 12636 18154 12664 18566
rect 12912 18154 12940 19790
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 13004 18970 13032 19654
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 12992 18828 13044 18834
rect 12992 18770 13044 18776
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12716 18148 12768 18154
rect 12716 18090 12768 18096
rect 12900 18148 12952 18154
rect 12900 18090 12952 18096
rect 12636 17746 12664 18090
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12452 17338 12480 17614
rect 12728 17542 12756 18090
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12728 17134 12756 17478
rect 12912 17338 12940 18090
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 12716 17128 12768 17134
rect 13004 17105 13032 18770
rect 12716 17070 12768 17076
rect 12990 17096 13046 17105
rect 12990 17031 13046 17040
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12544 16794 12572 16934
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 13004 16674 13032 17031
rect 13096 16794 13124 20012
rect 13268 19994 13320 20000
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13176 19916 13228 19922
rect 13176 19858 13228 19864
rect 13188 19446 13216 19858
rect 13280 19718 13308 19994
rect 13924 19922 13952 21014
rect 14016 20466 14044 21626
rect 14108 21418 14136 22766
rect 14188 22568 14240 22574
rect 14188 22510 14240 22516
rect 14096 21412 14148 21418
rect 14096 21354 14148 21360
rect 14200 21010 14228 22510
rect 14476 22506 14504 22918
rect 14464 22500 14516 22506
rect 14464 22442 14516 22448
rect 14335 22332 14643 22341
rect 14335 22330 14341 22332
rect 14397 22330 14421 22332
rect 14477 22330 14501 22332
rect 14557 22330 14581 22332
rect 14637 22330 14643 22332
rect 14397 22278 14399 22330
rect 14579 22278 14581 22330
rect 14335 22276 14341 22278
rect 14397 22276 14421 22278
rect 14477 22276 14501 22278
rect 14557 22276 14581 22278
rect 14637 22276 14643 22278
rect 14335 22267 14643 22276
rect 14752 22098 14780 23054
rect 14844 22574 14872 23122
rect 14832 22568 14884 22574
rect 14832 22510 14884 22516
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14335 21244 14643 21253
rect 14335 21242 14341 21244
rect 14397 21242 14421 21244
rect 14477 21242 14501 21244
rect 14557 21242 14581 21244
rect 14637 21242 14643 21244
rect 14397 21190 14399 21242
rect 14579 21190 14581 21242
rect 14335 21188 14341 21190
rect 14397 21188 14421 21190
rect 14477 21188 14501 21190
rect 14557 21188 14581 21190
rect 14637 21188 14643 21190
rect 14335 21179 14643 21188
rect 14188 21004 14240 21010
rect 14188 20946 14240 20952
rect 14752 20806 14780 22034
rect 14832 21412 14884 21418
rect 14832 21354 14884 21360
rect 14844 21146 14872 21354
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 14096 20800 14148 20806
rect 14094 20768 14096 20777
rect 14740 20800 14792 20806
rect 14148 20768 14150 20777
rect 14740 20742 14792 20748
rect 14094 20703 14150 20712
rect 14752 20466 14780 20742
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 14335 20156 14643 20165
rect 14335 20154 14341 20156
rect 14397 20154 14421 20156
rect 14477 20154 14501 20156
rect 14557 20154 14581 20156
rect 14637 20154 14643 20156
rect 14397 20102 14399 20154
rect 14579 20102 14581 20154
rect 14335 20100 14341 20102
rect 14397 20100 14421 20102
rect 14477 20100 14501 20102
rect 14557 20100 14581 20102
rect 14637 20100 14643 20102
rect 14335 20091 14643 20100
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 13912 19916 13964 19922
rect 13912 19858 13964 19864
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 13636 19848 13688 19854
rect 13636 19790 13688 19796
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13268 19712 13320 19718
rect 13268 19654 13320 19660
rect 13176 19440 13228 19446
rect 13176 19382 13228 19388
rect 13188 18902 13216 19382
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13372 18902 13400 19110
rect 13176 18896 13228 18902
rect 13176 18838 13228 18844
rect 13360 18896 13412 18902
rect 13360 18838 13412 18844
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13188 17678 13216 18362
rect 13280 17814 13308 18702
rect 13372 18426 13400 18702
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13372 17882 13400 18362
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13268 17808 13320 17814
rect 13268 17750 13320 17756
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 13188 16998 13216 17614
rect 13176 16992 13228 16998
rect 13176 16934 13228 16940
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 13004 16646 13124 16674
rect 13096 16454 13124 16646
rect 12992 16448 13044 16454
rect 12992 16390 13044 16396
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 13004 16046 13032 16390
rect 13280 16046 13308 17750
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13372 17649 13400 17682
rect 13358 17640 13414 17649
rect 13358 17575 13414 17584
rect 13372 17202 13400 17575
rect 13464 17338 13492 19722
rect 13648 19718 13676 19790
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13556 18698 13584 19314
rect 13544 18692 13596 18698
rect 13544 18634 13596 18640
rect 13556 17678 13584 18634
rect 13648 17678 13676 19654
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13740 18222 13768 19382
rect 13832 18630 13860 19858
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13924 18426 13952 19858
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 14016 18290 14044 19110
rect 14200 18970 14228 19858
rect 14335 19068 14643 19077
rect 14335 19066 14341 19068
rect 14397 19066 14421 19068
rect 14477 19066 14501 19068
rect 14557 19066 14581 19068
rect 14637 19066 14643 19068
rect 14397 19014 14399 19066
rect 14579 19014 14581 19066
rect 14335 19012 14341 19014
rect 14397 19012 14421 19014
rect 14477 19012 14501 19014
rect 14557 19012 14581 19014
rect 14637 19012 14643 19014
rect 14335 19003 14643 19012
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13740 17746 13768 17818
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 13464 16590 13492 17274
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13450 16416 13506 16425
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12360 14618 12388 14894
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12820 14550 12848 15846
rect 13096 15586 13124 15846
rect 13188 15706 13216 15982
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13096 15558 13216 15586
rect 12808 14544 12860 14550
rect 12808 14486 12860 14492
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11900 12866 11928 12922
rect 11900 12838 12112 12866
rect 12912 12850 12940 13126
rect 13004 12986 13032 13126
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11900 12434 11928 12650
rect 11980 12436 12032 12442
rect 11900 12406 11980 12434
rect 11980 12378 12032 12384
rect 12084 12322 12112 12838
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 11900 12294 12112 12322
rect 11900 12238 11928 12294
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 12176 12102 12204 12378
rect 12820 12306 12848 12582
rect 13096 12442 13124 12582
rect 13084 12436 13136 12442
rect 13188 12434 13216 15558
rect 13188 12406 13308 12434
rect 13084 12378 13136 12384
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 13096 12170 13124 12378
rect 13280 12170 13308 12406
rect 13372 12374 13400 16390
rect 13450 16351 13506 16360
rect 13464 15570 13492 16351
rect 13556 15978 13584 17614
rect 13648 16998 13676 17614
rect 14016 17542 14044 18226
rect 14335 17980 14643 17989
rect 14335 17978 14341 17980
rect 14397 17978 14421 17980
rect 14477 17978 14501 17980
rect 14557 17978 14581 17980
rect 14637 17978 14643 17980
rect 14397 17926 14399 17978
rect 14579 17926 14581 17978
rect 14335 17924 14341 17926
rect 14397 17924 14421 17926
rect 14477 17924 14501 17926
rect 14557 17924 14581 17926
rect 14637 17924 14643 17926
rect 14335 17915 14643 17924
rect 14752 17762 14780 19994
rect 14844 18834 14872 20198
rect 14936 20058 14964 25230
rect 15016 23248 15068 23254
rect 15014 23216 15016 23225
rect 15068 23216 15070 23225
rect 15014 23151 15070 23160
rect 15028 21486 15056 23151
rect 15108 22976 15160 22982
rect 15212 22964 15240 26318
rect 15292 25696 15344 25702
rect 15292 25638 15344 25644
rect 15304 25498 15332 25638
rect 15292 25492 15344 25498
rect 15292 25434 15344 25440
rect 16132 24818 16160 26386
rect 16592 26042 16620 26386
rect 16580 26036 16632 26042
rect 16580 25978 16632 25984
rect 16684 25922 16712 26862
rect 16776 26246 16804 26998
rect 18156 26926 18184 27814
rect 19260 27674 19288 27950
rect 19892 27872 19944 27878
rect 19892 27814 19944 27820
rect 20076 27872 20128 27878
rect 20076 27814 20128 27820
rect 21640 27872 21692 27878
rect 21640 27814 21692 27820
rect 23848 27872 23900 27878
rect 23848 27814 23900 27820
rect 25872 27872 25924 27878
rect 25872 27814 25924 27820
rect 19248 27668 19300 27674
rect 19248 27610 19300 27616
rect 19904 27606 19932 27814
rect 19892 27600 19944 27606
rect 19892 27542 19944 27548
rect 18328 27532 18380 27538
rect 18328 27474 18380 27480
rect 18340 27130 18368 27474
rect 19432 27328 19484 27334
rect 19432 27270 19484 27276
rect 18328 27124 18380 27130
rect 18328 27066 18380 27072
rect 18144 26920 18196 26926
rect 18144 26862 18196 26868
rect 19444 26858 19472 27270
rect 20088 26858 20116 27814
rect 21304 27772 21612 27781
rect 21304 27770 21310 27772
rect 21366 27770 21390 27772
rect 21446 27770 21470 27772
rect 21526 27770 21550 27772
rect 21606 27770 21612 27772
rect 21366 27718 21368 27770
rect 21548 27718 21550 27770
rect 21304 27716 21310 27718
rect 21366 27716 21390 27718
rect 21446 27716 21470 27718
rect 21526 27716 21550 27718
rect 21606 27716 21612 27718
rect 21304 27707 21612 27716
rect 21652 27674 21680 27814
rect 21640 27668 21692 27674
rect 21640 27610 21692 27616
rect 22836 27532 22888 27538
rect 22836 27474 22888 27480
rect 23296 27532 23348 27538
rect 23296 27474 23348 27480
rect 20628 27396 20680 27402
rect 20628 27338 20680 27344
rect 20444 26920 20496 26926
rect 20444 26862 20496 26868
rect 19432 26852 19484 26858
rect 19432 26794 19484 26800
rect 20076 26852 20128 26858
rect 20076 26794 20128 26800
rect 16948 26784 17000 26790
rect 16948 26726 17000 26732
rect 18144 26784 18196 26790
rect 18144 26726 18196 26732
rect 20352 26784 20404 26790
rect 20352 26726 20404 26732
rect 16960 26586 16988 26726
rect 16948 26580 17000 26586
rect 16948 26522 17000 26528
rect 16764 26240 16816 26246
rect 16764 26182 16816 26188
rect 16856 26240 16908 26246
rect 16856 26182 16908 26188
rect 16592 25894 16712 25922
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 15568 24404 15620 24410
rect 15568 24346 15620 24352
rect 15580 23798 15608 24346
rect 16132 24274 16160 24754
rect 16120 24268 16172 24274
rect 16120 24210 16172 24216
rect 16132 23866 16160 24210
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 15568 23792 15620 23798
rect 15568 23734 15620 23740
rect 15580 23254 15608 23734
rect 15292 23248 15344 23254
rect 15292 23190 15344 23196
rect 15568 23248 15620 23254
rect 15568 23190 15620 23196
rect 15160 22936 15240 22964
rect 15108 22918 15160 22924
rect 15120 22030 15148 22918
rect 15304 22710 15332 23190
rect 15292 22704 15344 22710
rect 15292 22646 15344 22652
rect 15108 22024 15160 22030
rect 15108 21966 15160 21972
rect 15120 21894 15148 21966
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 15672 21690 15700 23802
rect 15844 22976 15896 22982
rect 15842 22944 15844 22953
rect 15896 22944 15898 22953
rect 15842 22879 15898 22888
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 15856 21690 15884 22578
rect 16120 22160 16172 22166
rect 16120 22102 16172 22108
rect 15660 21684 15712 21690
rect 15660 21626 15712 21632
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 15016 21480 15068 21486
rect 15016 21422 15068 21428
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 15856 21146 15884 21286
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 14924 20052 14976 20058
rect 14924 19994 14976 20000
rect 15028 19242 15056 20946
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15396 20058 15424 20402
rect 15384 20052 15436 20058
rect 15304 20012 15384 20040
rect 15016 19236 15068 19242
rect 15016 19178 15068 19184
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 14832 18080 14884 18086
rect 14832 18022 14884 18028
rect 14568 17734 14780 17762
rect 14844 17746 14872 18022
rect 14832 17740 14884 17746
rect 14568 17678 14596 17734
rect 15016 17740 15068 17746
rect 14832 17682 14884 17688
rect 14936 17700 15016 17728
rect 14556 17672 14608 17678
rect 14648 17672 14700 17678
rect 14556 17614 14608 17620
rect 14646 17640 14648 17649
rect 14700 17640 14702 17649
rect 14464 17604 14516 17610
rect 14464 17546 14516 17552
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 14476 17354 14504 17546
rect 14568 17542 14596 17614
rect 14646 17575 14702 17584
rect 14660 17542 14688 17575
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14936 17354 14964 17700
rect 15016 17682 15068 17688
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 15120 17354 15148 17682
rect 14004 17332 14056 17338
rect 14476 17326 14964 17354
rect 15028 17326 15148 17354
rect 15304 17338 15332 20012
rect 15384 19994 15436 20000
rect 16132 19990 16160 22102
rect 16304 21480 16356 21486
rect 16304 21422 16356 21428
rect 16316 20602 16344 21422
rect 16408 20602 16436 22714
rect 16488 22432 16540 22438
rect 16488 22374 16540 22380
rect 16500 22030 16528 22374
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16500 21146 16528 21966
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16304 20596 16356 20602
rect 16304 20538 16356 20544
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16408 20058 16436 20538
rect 16592 20398 16620 25894
rect 16776 25362 16804 26182
rect 16868 25430 16896 26182
rect 17820 26140 18128 26149
rect 17820 26138 17826 26140
rect 17882 26138 17906 26140
rect 17962 26138 17986 26140
rect 18042 26138 18066 26140
rect 18122 26138 18128 26140
rect 17882 26086 17884 26138
rect 18064 26086 18066 26138
rect 17820 26084 17826 26086
rect 17882 26084 17906 26086
rect 17962 26084 17986 26086
rect 18042 26084 18066 26086
rect 18122 26084 18128 26086
rect 17820 26075 18128 26084
rect 18156 25974 18184 26726
rect 19708 26308 19760 26314
rect 19708 26250 19760 26256
rect 18236 26240 18288 26246
rect 18236 26182 18288 26188
rect 18144 25968 18196 25974
rect 18144 25910 18196 25916
rect 16856 25424 16908 25430
rect 16856 25366 16908 25372
rect 16764 25356 16816 25362
rect 16764 25298 16816 25304
rect 18156 25158 18184 25910
rect 17132 25152 17184 25158
rect 17132 25094 17184 25100
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 17040 24064 17092 24070
rect 17040 24006 17092 24012
rect 16764 23792 16816 23798
rect 16764 23734 16816 23740
rect 16776 23186 16804 23734
rect 16856 23588 16908 23594
rect 16856 23530 16908 23536
rect 16868 23186 16896 23530
rect 16764 23180 16816 23186
rect 16764 23122 16816 23128
rect 16856 23180 16908 23186
rect 16856 23122 16908 23128
rect 16856 22976 16908 22982
rect 16856 22918 16908 22924
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16580 20392 16632 20398
rect 16580 20334 16632 20340
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 16120 19984 16172 19990
rect 16120 19926 16172 19932
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15396 18086 15424 19246
rect 16592 19174 16620 20334
rect 16580 19168 16632 19174
rect 16580 19110 16632 19116
rect 16488 18148 16540 18154
rect 16488 18090 16540 18096
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 16500 17678 16528 18090
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 15292 17332 15344 17338
rect 14004 17274 14056 17280
rect 14016 16998 14044 17274
rect 15028 17082 15056 17326
rect 15292 17274 15344 17280
rect 14936 17054 15056 17082
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 14016 16046 14044 16934
rect 14335 16892 14643 16901
rect 14335 16890 14341 16892
rect 14397 16890 14421 16892
rect 14477 16890 14501 16892
rect 14557 16890 14581 16892
rect 14637 16890 14643 16892
rect 14397 16838 14399 16890
rect 14579 16838 14581 16890
rect 14335 16836 14341 16838
rect 14397 16836 14421 16838
rect 14477 16836 14501 16838
rect 14557 16836 14581 16838
rect 14637 16836 14643 16838
rect 14335 16827 14643 16836
rect 14936 16726 14964 17054
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 15028 16726 15056 16934
rect 15212 16726 15240 17070
rect 15488 16794 15516 17070
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 14924 16720 14976 16726
rect 14924 16662 14976 16668
rect 15016 16720 15068 16726
rect 15016 16662 15068 16668
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 15568 16720 15620 16726
rect 15568 16662 15620 16668
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13648 15706 13676 15846
rect 14335 15804 14643 15813
rect 14335 15802 14341 15804
rect 14397 15802 14421 15804
rect 14477 15802 14501 15804
rect 14557 15802 14581 15804
rect 14637 15802 14643 15804
rect 14397 15750 14399 15802
rect 14579 15750 14581 15802
rect 14335 15748 14341 15750
rect 14397 15748 14421 15750
rect 14477 15748 14501 15750
rect 14557 15748 14581 15750
rect 14637 15748 14643 15750
rect 14335 15739 14643 15748
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 13912 15088 13964 15094
rect 13912 15030 13964 15036
rect 13820 14884 13872 14890
rect 13820 14826 13872 14832
rect 13832 14618 13860 14826
rect 13924 14822 13952 15030
rect 14096 14952 14148 14958
rect 14096 14894 14148 14900
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13452 13728 13504 13734
rect 13452 13670 13504 13676
rect 13464 12889 13492 13670
rect 13648 13462 13676 13806
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13636 13456 13688 13462
rect 13636 13398 13688 13404
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13556 12986 13584 13126
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13450 12880 13506 12889
rect 13450 12815 13506 12824
rect 13464 12714 13492 12815
rect 13740 12714 13768 13670
rect 13832 13462 13860 13806
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13924 13258 13952 14758
rect 14016 14618 14044 14758
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14108 14482 14136 14894
rect 14200 14822 14228 15438
rect 14844 14958 14872 16050
rect 15028 15910 15056 16662
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15304 16250 15332 16526
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15580 16046 15608 16662
rect 15568 16040 15620 16046
rect 15568 15982 15620 15988
rect 15016 15904 15068 15910
rect 15016 15846 15068 15852
rect 15028 14958 15056 15846
rect 14832 14952 14884 14958
rect 15016 14952 15068 14958
rect 14884 14912 14964 14940
rect 14832 14894 14884 14900
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 14016 13326 14044 14350
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 13912 13252 13964 13258
rect 13912 13194 13964 13200
rect 13924 12753 13952 13194
rect 13910 12744 13966 12753
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13728 12708 13780 12714
rect 14016 12714 14044 13262
rect 13910 12679 13966 12688
rect 14004 12708 14056 12714
rect 13728 12650 13780 12656
rect 14004 12650 14056 12656
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13360 12368 13412 12374
rect 13360 12310 13412 12316
rect 13556 12238 13584 12582
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13084 12164 13136 12170
rect 13084 12106 13136 12112
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 13096 11626 13124 12106
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 13280 11558 13308 12106
rect 13740 12102 13768 12650
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 14108 11830 14136 14418
rect 14200 13530 14228 14758
rect 14335 14716 14643 14725
rect 14335 14714 14341 14716
rect 14397 14714 14421 14716
rect 14477 14714 14501 14716
rect 14557 14714 14581 14716
rect 14637 14714 14643 14716
rect 14397 14662 14399 14714
rect 14579 14662 14581 14714
rect 14335 14660 14341 14662
rect 14397 14660 14421 14662
rect 14477 14660 14501 14662
rect 14557 14660 14581 14662
rect 14637 14660 14643 14662
rect 14335 14651 14643 14660
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14335 13628 14643 13637
rect 14335 13626 14341 13628
rect 14397 13626 14421 13628
rect 14477 13626 14501 13628
rect 14557 13626 14581 13628
rect 14637 13626 14643 13628
rect 14397 13574 14399 13626
rect 14579 13574 14581 13626
rect 14335 13572 14341 13574
rect 14397 13572 14421 13574
rect 14477 13572 14501 13574
rect 14557 13572 14581 13574
rect 14637 13572 14643 13574
rect 14335 13563 14643 13572
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14752 13462 14780 14418
rect 14936 14346 14964 14912
rect 15016 14894 15068 14900
rect 14924 14340 14976 14346
rect 14924 14282 14976 14288
rect 14740 13456 14792 13462
rect 14740 13398 14792 13404
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13464 11642 13492 11698
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13372 11354 13400 11630
rect 13464 11614 13584 11642
rect 13556 11558 13584 11614
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 14108 11286 14136 11766
rect 14200 11626 14228 13330
rect 14384 13240 14412 13330
rect 14556 13252 14608 13258
rect 14384 13212 14556 13240
rect 14384 12782 14412 13212
rect 14556 13194 14608 13200
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14335 12540 14643 12549
rect 14335 12538 14341 12540
rect 14397 12538 14421 12540
rect 14477 12538 14501 12540
rect 14557 12538 14581 12540
rect 14637 12538 14643 12540
rect 14397 12486 14399 12538
rect 14579 12486 14581 12538
rect 14335 12484 14341 12486
rect 14397 12484 14421 12486
rect 14477 12484 14501 12486
rect 14557 12484 14581 12486
rect 14637 12484 14643 12486
rect 14335 12475 14643 12484
rect 14752 11694 14780 12854
rect 14844 12714 14872 13126
rect 14832 12708 14884 12714
rect 14832 12650 14884 12656
rect 14936 12594 14964 14282
rect 15028 14278 15056 14894
rect 15580 14618 15608 15982
rect 15672 14958 15700 17614
rect 16684 17202 16712 21830
rect 16762 21448 16818 21457
rect 16762 21383 16818 21392
rect 16776 21350 16804 21383
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16776 20466 16804 20878
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16776 20058 16804 20402
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 16868 18834 16896 22918
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16960 19514 16988 20402
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 16856 18828 16908 18834
rect 16856 18770 16908 18776
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16776 17746 16804 18226
rect 17052 18222 17080 24006
rect 17144 23662 17172 25094
rect 17820 25052 18128 25061
rect 17820 25050 17826 25052
rect 17882 25050 17906 25052
rect 17962 25050 17986 25052
rect 18042 25050 18066 25052
rect 18122 25050 18128 25052
rect 17882 24998 17884 25050
rect 18064 24998 18066 25050
rect 17820 24996 17826 24998
rect 17882 24996 17906 24998
rect 17962 24996 17986 24998
rect 18042 24996 18066 24998
rect 18122 24996 18128 24998
rect 17820 24987 18128 24996
rect 18156 24682 18184 25094
rect 18144 24676 18196 24682
rect 18144 24618 18196 24624
rect 18052 24268 18104 24274
rect 18052 24210 18104 24216
rect 17684 24064 17736 24070
rect 18064 24052 18092 24210
rect 18064 24024 18184 24052
rect 17684 24006 17736 24012
rect 17696 23798 17724 24006
rect 17820 23964 18128 23973
rect 17820 23962 17826 23964
rect 17882 23962 17906 23964
rect 17962 23962 17986 23964
rect 18042 23962 18066 23964
rect 18122 23962 18128 23964
rect 17882 23910 17884 23962
rect 18064 23910 18066 23962
rect 17820 23908 17826 23910
rect 17882 23908 17906 23910
rect 17962 23908 17986 23910
rect 18042 23908 18066 23910
rect 18122 23908 18128 23910
rect 17820 23899 18128 23908
rect 17684 23792 17736 23798
rect 17684 23734 17736 23740
rect 17132 23656 17184 23662
rect 18156 23610 18184 24024
rect 17132 23598 17184 23604
rect 17408 23588 17460 23594
rect 17408 23530 17460 23536
rect 17868 23588 17920 23594
rect 17868 23530 17920 23536
rect 18064 23582 18184 23610
rect 17224 23180 17276 23186
rect 17224 23122 17276 23128
rect 17316 23180 17368 23186
rect 17316 23122 17368 23128
rect 17236 22166 17264 23122
rect 17328 23089 17356 23122
rect 17314 23080 17370 23089
rect 17314 23015 17370 23024
rect 17224 22160 17276 22166
rect 17224 22102 17276 22108
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 17236 21486 17264 21626
rect 17224 21480 17276 21486
rect 17224 21422 17276 21428
rect 17132 21004 17184 21010
rect 17132 20946 17184 20952
rect 17144 20466 17172 20946
rect 17224 20800 17276 20806
rect 17224 20742 17276 20748
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17236 20262 17264 20742
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17236 20058 17264 20198
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17420 19446 17448 23530
rect 17880 23322 17908 23530
rect 17868 23316 17920 23322
rect 17868 23258 17920 23264
rect 18064 23118 18092 23582
rect 18144 23520 18196 23526
rect 18144 23462 18196 23468
rect 18052 23112 18104 23118
rect 18052 23054 18104 23060
rect 18156 22982 18184 23462
rect 17592 22976 17644 22982
rect 17592 22918 17644 22924
rect 18144 22976 18196 22982
rect 18144 22918 18196 22924
rect 17604 21486 17632 22918
rect 17820 22876 18128 22885
rect 17820 22874 17826 22876
rect 17882 22874 17906 22876
rect 17962 22874 17986 22876
rect 18042 22874 18066 22876
rect 18122 22874 18128 22876
rect 17882 22822 17884 22874
rect 18064 22822 18066 22874
rect 17820 22820 17826 22822
rect 17882 22820 17906 22822
rect 17962 22820 17986 22822
rect 18042 22820 18066 22822
rect 18122 22820 18128 22822
rect 17820 22811 18128 22820
rect 18248 22642 18276 26182
rect 18420 25832 18472 25838
rect 18420 25774 18472 25780
rect 18432 25498 18460 25774
rect 18696 25696 18748 25702
rect 18696 25638 18748 25644
rect 18420 25492 18472 25498
rect 18420 25434 18472 25440
rect 18328 25424 18380 25430
rect 18604 25424 18656 25430
rect 18328 25366 18380 25372
rect 18602 25392 18604 25401
rect 18656 25392 18658 25401
rect 18340 24954 18368 25366
rect 18602 25327 18658 25336
rect 18708 25294 18736 25638
rect 19616 25356 19668 25362
rect 19616 25298 19668 25304
rect 18696 25288 18748 25294
rect 18696 25230 18748 25236
rect 19628 24954 19656 25298
rect 18328 24948 18380 24954
rect 18328 24890 18380 24896
rect 19248 24948 19300 24954
rect 19248 24890 19300 24896
rect 19616 24948 19668 24954
rect 19616 24890 19668 24896
rect 19260 24614 19288 24890
rect 19616 24676 19668 24682
rect 19616 24618 19668 24624
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18788 24608 18840 24614
rect 18788 24550 18840 24556
rect 19248 24608 19300 24614
rect 19248 24550 19300 24556
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 18524 24274 18552 24550
rect 18800 24410 18828 24550
rect 18788 24404 18840 24410
rect 18788 24346 18840 24352
rect 18616 24274 18920 24290
rect 18512 24268 18564 24274
rect 18512 24210 18564 24216
rect 18604 24268 18920 24274
rect 18656 24262 18920 24268
rect 18604 24210 18656 24216
rect 18328 24064 18380 24070
rect 18328 24006 18380 24012
rect 18420 24064 18472 24070
rect 18420 24006 18472 24012
rect 18340 23186 18368 24006
rect 18432 23186 18460 24006
rect 18328 23180 18380 23186
rect 18328 23122 18380 23128
rect 18420 23180 18472 23186
rect 18524 23168 18552 24210
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 18800 23730 18828 24142
rect 18788 23724 18840 23730
rect 18788 23666 18840 23672
rect 18800 23186 18828 23666
rect 18892 23186 18920 24262
rect 18972 23656 19024 23662
rect 18972 23598 19024 23604
rect 18696 23180 18748 23186
rect 18524 23140 18696 23168
rect 18420 23122 18472 23128
rect 18696 23122 18748 23128
rect 18788 23180 18840 23186
rect 18788 23122 18840 23128
rect 18880 23180 18932 23186
rect 18880 23122 18932 23128
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18144 22500 18196 22506
rect 18144 22442 18196 22448
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17696 21554 17724 21830
rect 17820 21788 18128 21797
rect 17820 21786 17826 21788
rect 17882 21786 17906 21788
rect 17962 21786 17986 21788
rect 18042 21786 18066 21788
rect 18122 21786 18128 21788
rect 17882 21734 17884 21786
rect 18064 21734 18066 21786
rect 17820 21732 17826 21734
rect 17882 21732 17906 21734
rect 17962 21732 17986 21734
rect 18042 21732 18066 21734
rect 18122 21732 18128 21734
rect 17820 21723 18128 21732
rect 18156 21604 18184 22442
rect 18064 21576 18184 21604
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17592 21480 17644 21486
rect 17592 21422 17644 21428
rect 17604 21010 17632 21422
rect 17696 21010 17724 21490
rect 18064 21486 18092 21576
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17684 21004 17736 21010
rect 17684 20946 17736 20952
rect 17820 20700 18128 20709
rect 17820 20698 17826 20700
rect 17882 20698 17906 20700
rect 17962 20698 17986 20700
rect 18042 20698 18066 20700
rect 18122 20698 18128 20700
rect 17882 20646 17884 20698
rect 18064 20646 18066 20698
rect 17820 20644 17826 20646
rect 17882 20644 17906 20646
rect 17962 20644 17986 20646
rect 18042 20644 18066 20646
rect 18122 20644 18128 20646
rect 17820 20635 18128 20644
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 17820 19612 18128 19621
rect 17820 19610 17826 19612
rect 17882 19610 17906 19612
rect 17962 19610 17986 19612
rect 18042 19610 18066 19612
rect 18122 19610 18128 19612
rect 17882 19558 17884 19610
rect 18064 19558 18066 19610
rect 17820 19556 17826 19558
rect 17882 19556 17906 19558
rect 17962 19556 17986 19558
rect 18042 19556 18066 19558
rect 18122 19556 18128 19558
rect 17820 19547 18128 19556
rect 17408 19440 17460 19446
rect 18156 19394 18184 20198
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 17408 19382 17460 19388
rect 17972 19366 18184 19394
rect 17972 19310 18000 19366
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17420 18902 17448 19246
rect 17408 18896 17460 18902
rect 17408 18838 17460 18844
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 16764 17740 16816 17746
rect 16764 17682 16816 17688
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 16948 17536 17000 17542
rect 16948 17478 17000 17484
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 15936 17128 15988 17134
rect 16868 17105 16896 17138
rect 15936 17070 15988 17076
rect 16854 17096 16910 17105
rect 15844 17060 15896 17066
rect 15844 17002 15896 17008
rect 15856 16658 15884 17002
rect 15948 16658 15976 17070
rect 16212 17060 16264 17066
rect 16212 17002 16264 17008
rect 16396 17060 16448 17066
rect 16854 17031 16910 17040
rect 16396 17002 16448 17008
rect 16224 16726 16252 17002
rect 16212 16720 16264 16726
rect 16212 16662 16264 16668
rect 16408 16658 16436 17002
rect 16580 16720 16632 16726
rect 16580 16662 16632 16668
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16592 16522 16620 16662
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15752 16176 15804 16182
rect 15750 16144 15752 16153
rect 15804 16144 15806 16153
rect 15750 16079 15806 16088
rect 15948 16017 15976 16390
rect 16592 16046 16620 16458
rect 16580 16040 16632 16046
rect 15934 16008 15990 16017
rect 16580 15982 16632 15988
rect 15934 15943 15990 15952
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 16120 14884 16172 14890
rect 16120 14826 16172 14832
rect 16132 14618 16160 14826
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16960 14482 16988 17478
rect 17052 17338 17080 17614
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 17420 17218 17448 18566
rect 17512 18358 17540 18770
rect 17604 18426 17632 18770
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 17696 17746 17724 19246
rect 17972 18970 18000 19246
rect 18064 18970 18092 19246
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 17820 18524 18128 18533
rect 17820 18522 17826 18524
rect 17882 18522 17906 18524
rect 17962 18522 17986 18524
rect 18042 18522 18066 18524
rect 18122 18522 18128 18524
rect 17882 18470 17884 18522
rect 18064 18470 18066 18522
rect 17820 18468 17826 18470
rect 17882 18468 17906 18470
rect 17962 18468 17986 18470
rect 18042 18468 18066 18470
rect 18122 18468 18128 18470
rect 17820 18459 18128 18468
rect 18156 18222 18184 19366
rect 18248 19310 18276 19654
rect 18512 19372 18564 19378
rect 18708 19334 18736 23122
rect 18786 23080 18842 23089
rect 18892 23066 18920 23122
rect 18842 23038 18920 23066
rect 18786 23015 18842 23024
rect 18984 22982 19012 23598
rect 19064 23180 19116 23186
rect 19064 23122 19116 23128
rect 18972 22976 19024 22982
rect 18972 22918 19024 22924
rect 18984 22710 19012 22918
rect 19076 22778 19104 23122
rect 19156 22976 19208 22982
rect 19156 22918 19208 22924
rect 19064 22772 19116 22778
rect 19064 22714 19116 22720
rect 18972 22704 19024 22710
rect 18972 22646 19024 22652
rect 19168 22642 19196 22918
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 18880 22160 18932 22166
rect 18880 22102 18932 22108
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18512 19314 18564 19320
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18340 18902 18368 19246
rect 18328 18896 18380 18902
rect 18328 18838 18380 18844
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18328 18148 18380 18154
rect 18328 18090 18380 18096
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 17820 17436 18128 17445
rect 17820 17434 17826 17436
rect 17882 17434 17906 17436
rect 17962 17434 17986 17436
rect 18042 17434 18066 17436
rect 18122 17434 18128 17436
rect 17882 17382 17884 17434
rect 18064 17382 18066 17434
rect 17820 17380 17826 17382
rect 17882 17380 17906 17382
rect 17962 17380 17986 17382
rect 18042 17380 18066 17382
rect 18122 17380 18128 17382
rect 17820 17371 18128 17380
rect 17420 17190 17632 17218
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 17132 16040 17184 16046
rect 17236 16028 17264 16526
rect 17316 16516 17368 16522
rect 17316 16458 17368 16464
rect 17184 16000 17264 16028
rect 17132 15982 17184 15988
rect 17052 15570 17080 15982
rect 17236 15570 17264 16000
rect 17328 15706 17356 16458
rect 17420 16250 17448 17070
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17512 16794 17540 16934
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17408 16244 17460 16250
rect 17408 16186 17460 16192
rect 17512 16046 17540 16526
rect 17604 16454 17632 17190
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17972 16794 18000 17070
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 17500 16040 17552 16046
rect 17500 15982 17552 15988
rect 17604 15910 17632 16390
rect 17820 16348 18128 16357
rect 17820 16346 17826 16348
rect 17882 16346 17906 16348
rect 17962 16346 17986 16348
rect 18042 16346 18066 16348
rect 18122 16346 18128 16348
rect 17882 16294 17884 16346
rect 18064 16294 18066 16346
rect 17820 16292 17826 16294
rect 17882 16292 17906 16294
rect 17962 16292 17986 16294
rect 18042 16292 18066 16294
rect 18122 16292 18128 16294
rect 17820 16283 18128 16292
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17774 16144 17830 16153
rect 17774 16079 17830 16088
rect 17788 15910 17816 16079
rect 17868 16040 17920 16046
rect 17866 16008 17868 16017
rect 17920 16008 17922 16017
rect 17866 15943 17922 15952
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17972 15706 18000 16186
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17052 14890 17080 15506
rect 17236 15094 17264 15506
rect 17328 15366 17356 15642
rect 18156 15502 18184 17138
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17040 14884 17092 14890
rect 17040 14826 17092 14832
rect 17328 14618 17356 15302
rect 17820 15260 18128 15269
rect 17820 15258 17826 15260
rect 17882 15258 17906 15260
rect 17962 15258 17986 15260
rect 18042 15258 18066 15260
rect 18122 15258 18128 15260
rect 17882 15206 17884 15258
rect 18064 15206 18066 15258
rect 17820 15204 17826 15206
rect 17882 15204 17906 15206
rect 17962 15204 17986 15206
rect 18042 15204 18066 15206
rect 18122 15204 18128 15206
rect 17820 15195 18128 15204
rect 18340 15026 18368 18090
rect 18524 16046 18552 19314
rect 18616 19306 18736 19334
rect 18616 17134 18644 19306
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 18708 17202 18736 17818
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18604 16992 18656 16998
rect 18604 16934 18656 16940
rect 18616 16454 18644 16934
rect 18708 16794 18736 17138
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18708 15502 18736 16594
rect 18800 16250 18828 21966
rect 18892 21690 18920 22102
rect 19076 22094 19104 22510
rect 19076 22066 19196 22094
rect 18880 21684 18932 21690
rect 18880 21626 18932 21632
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 18984 21146 19012 21422
rect 18972 21140 19024 21146
rect 18972 21082 19024 21088
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 18984 20330 19012 20878
rect 18972 20324 19024 20330
rect 18972 20266 19024 20272
rect 18880 19712 18932 19718
rect 18880 19654 18932 19660
rect 18892 18970 18920 19654
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 19168 18816 19196 22066
rect 19260 20806 19288 24550
rect 19340 22704 19392 22710
rect 19340 22646 19392 22652
rect 19352 21486 19380 22646
rect 19444 22098 19472 24550
rect 19628 24206 19656 24618
rect 19616 24200 19668 24206
rect 19616 24142 19668 24148
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19260 18834 19288 20742
rect 19352 20602 19380 21422
rect 19628 21400 19656 24142
rect 19720 22234 19748 26250
rect 20364 25838 20392 26726
rect 20456 26246 20484 26862
rect 20444 26240 20496 26246
rect 20444 26182 20496 26188
rect 20456 25906 20484 26182
rect 20444 25900 20496 25906
rect 20444 25842 20496 25848
rect 19984 25832 20036 25838
rect 19984 25774 20036 25780
rect 20352 25832 20404 25838
rect 20352 25774 20404 25780
rect 19996 25158 20024 25774
rect 19984 25152 20036 25158
rect 19984 25094 20036 25100
rect 19996 23866 20024 25094
rect 20640 24614 20668 27338
rect 20720 27328 20772 27334
rect 20720 27270 20772 27276
rect 20904 27328 20956 27334
rect 20904 27270 20956 27276
rect 20628 24608 20680 24614
rect 20628 24550 20680 24556
rect 20352 24268 20404 24274
rect 20352 24210 20404 24216
rect 19984 23860 20036 23866
rect 19984 23802 20036 23808
rect 20260 22704 20312 22710
rect 20260 22646 20312 22652
rect 20272 22506 20300 22646
rect 20364 22556 20392 24210
rect 20536 24200 20588 24206
rect 20536 24142 20588 24148
rect 20548 23866 20576 24142
rect 20536 23860 20588 23866
rect 20536 23802 20588 23808
rect 20732 22710 20760 27270
rect 20916 26926 20944 27270
rect 22848 27130 22876 27474
rect 22928 27328 22980 27334
rect 22928 27270 22980 27276
rect 22836 27124 22888 27130
rect 22836 27066 22888 27072
rect 20904 26920 20956 26926
rect 20904 26862 20956 26868
rect 21304 26684 21612 26693
rect 21304 26682 21310 26684
rect 21366 26682 21390 26684
rect 21446 26682 21470 26684
rect 21526 26682 21550 26684
rect 21606 26682 21612 26684
rect 21366 26630 21368 26682
rect 21548 26630 21550 26682
rect 21304 26628 21310 26630
rect 21366 26628 21390 26630
rect 21446 26628 21470 26630
rect 21526 26628 21550 26630
rect 21606 26628 21612 26630
rect 21304 26619 21612 26628
rect 20812 26444 20864 26450
rect 20812 26386 20864 26392
rect 20824 26042 20852 26386
rect 20812 26036 20864 26042
rect 20812 25978 20864 25984
rect 22940 25838 22968 27270
rect 23308 27130 23336 27474
rect 23296 27124 23348 27130
rect 23296 27066 23348 27072
rect 23860 26926 23888 27814
rect 24400 27328 24452 27334
rect 24400 27270 24452 27276
rect 24412 27130 24440 27270
rect 24789 27228 25097 27237
rect 24789 27226 24795 27228
rect 24851 27226 24875 27228
rect 24931 27226 24955 27228
rect 25011 27226 25035 27228
rect 25091 27226 25097 27228
rect 24851 27174 24853 27226
rect 25033 27174 25035 27226
rect 24789 27172 24795 27174
rect 24851 27172 24875 27174
rect 24931 27172 24955 27174
rect 25011 27172 25035 27174
rect 25091 27172 25097 27174
rect 24789 27163 25097 27172
rect 24400 27124 24452 27130
rect 24400 27066 24452 27072
rect 23848 26920 23900 26926
rect 23848 26862 23900 26868
rect 25884 26858 25912 27814
rect 23756 26852 23808 26858
rect 23756 26794 23808 26800
rect 25872 26852 25924 26858
rect 25872 26794 25924 26800
rect 22928 25832 22980 25838
rect 22928 25774 22980 25780
rect 21732 25764 21784 25770
rect 21732 25706 21784 25712
rect 21304 25596 21612 25605
rect 21304 25594 21310 25596
rect 21366 25594 21390 25596
rect 21446 25594 21470 25596
rect 21526 25594 21550 25596
rect 21606 25594 21612 25596
rect 21366 25542 21368 25594
rect 21548 25542 21550 25594
rect 21304 25540 21310 25542
rect 21366 25540 21390 25542
rect 21446 25540 21470 25542
rect 21526 25540 21550 25542
rect 21606 25540 21612 25542
rect 21304 25531 21612 25540
rect 21744 25498 21772 25706
rect 22652 25696 22704 25702
rect 22652 25638 22704 25644
rect 21732 25492 21784 25498
rect 21732 25434 21784 25440
rect 21456 25356 21508 25362
rect 21456 25298 21508 25304
rect 20996 25152 21048 25158
rect 20996 25094 21048 25100
rect 20812 24812 20864 24818
rect 20812 24754 20864 24760
rect 20824 23730 20852 24754
rect 21008 24138 21036 25094
rect 21468 24954 21496 25298
rect 22664 24954 22692 25638
rect 23204 25288 23256 25294
rect 23204 25230 23256 25236
rect 22928 25152 22980 25158
rect 22928 25094 22980 25100
rect 21456 24948 21508 24954
rect 21456 24890 21508 24896
rect 22652 24948 22704 24954
rect 22652 24890 22704 24896
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 21824 24744 21876 24750
rect 21824 24686 21876 24692
rect 21088 24608 21140 24614
rect 21088 24550 21140 24556
rect 20996 24132 21048 24138
rect 20996 24074 21048 24080
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 21008 23662 21036 24074
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 21008 23322 21036 23598
rect 20996 23316 21048 23322
rect 20996 23258 21048 23264
rect 20812 22772 20864 22778
rect 20812 22714 20864 22720
rect 20720 22704 20772 22710
rect 20720 22646 20772 22652
rect 20536 22568 20588 22574
rect 20364 22528 20536 22556
rect 20260 22500 20312 22506
rect 20260 22442 20312 22448
rect 19708 22228 19760 22234
rect 19708 22170 19760 22176
rect 20272 22098 20300 22442
rect 20260 22092 20312 22098
rect 20260 22034 20312 22040
rect 20272 21894 20300 22034
rect 20364 21962 20392 22528
rect 20536 22510 20588 22516
rect 20536 22432 20588 22438
rect 20536 22374 20588 22380
rect 20548 22098 20576 22374
rect 20536 22092 20588 22098
rect 20536 22034 20588 22040
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 20260 21888 20312 21894
rect 20260 21830 20312 21836
rect 19708 21412 19760 21418
rect 19628 21372 19708 21400
rect 19708 21354 19760 21360
rect 19984 21412 20036 21418
rect 19984 21354 20036 21360
rect 19524 21344 19576 21350
rect 19444 21304 19524 21332
rect 19444 20942 19472 21304
rect 19524 21286 19576 21292
rect 19524 21072 19576 21078
rect 19524 21014 19576 21020
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19536 20602 19564 21014
rect 19720 21010 19748 21354
rect 19996 21078 20024 21354
rect 20272 21350 20300 21830
rect 20352 21480 20404 21486
rect 20352 21422 20404 21428
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 19984 21072 20036 21078
rect 19984 21014 20036 21020
rect 20272 21010 20300 21286
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 20076 21004 20128 21010
rect 20076 20946 20128 20952
rect 20260 21004 20312 21010
rect 20260 20946 20312 20952
rect 20088 20806 20116 20946
rect 20076 20800 20128 20806
rect 20076 20742 20128 20748
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19352 19854 19380 20538
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 20088 19514 20116 19790
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 20168 19372 20220 19378
rect 20168 19314 20220 19320
rect 19076 18788 19196 18816
rect 19248 18828 19300 18834
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18788 15088 18840 15094
rect 18788 15030 18840 15036
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 15028 12782 15056 13126
rect 15212 12850 15240 13330
rect 15580 13190 15608 13398
rect 15856 13394 15884 14214
rect 17820 14172 18128 14181
rect 17820 14170 17826 14172
rect 17882 14170 17906 14172
rect 17962 14170 17986 14172
rect 18042 14170 18066 14172
rect 18122 14170 18128 14172
rect 17882 14118 17884 14170
rect 18064 14118 18066 14170
rect 17820 14116 17826 14118
rect 17882 14116 17906 14118
rect 17962 14116 17986 14118
rect 18042 14116 18066 14118
rect 18122 14116 18128 14118
rect 17820 14107 18128 14116
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16316 13394 16344 13466
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16132 12850 16160 13126
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 15016 12776 15068 12782
rect 15292 12776 15344 12782
rect 15016 12718 15068 12724
rect 15120 12724 15292 12730
rect 15120 12718 15344 12724
rect 15120 12702 15332 12718
rect 15120 12646 15148 12702
rect 15108 12640 15160 12646
rect 14844 12566 14964 12594
rect 15014 12608 15070 12617
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14200 11354 14228 11562
rect 14335 11452 14643 11461
rect 14335 11450 14341 11452
rect 14397 11450 14421 11452
rect 14477 11450 14501 11452
rect 14557 11450 14581 11452
rect 14637 11450 14643 11452
rect 14397 11398 14399 11450
rect 14579 11398 14581 11450
rect 14335 11396 14341 11398
rect 14397 11396 14421 11398
rect 14477 11396 14501 11398
rect 14557 11396 14581 11398
rect 14637 11396 14643 11398
rect 14335 11387 14643 11396
rect 14844 11354 14872 12566
rect 15108 12582 15160 12588
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15014 12543 15070 12552
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14936 11898 14964 12038
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14096 11280 14148 11286
rect 14096 11222 14148 11228
rect 14844 11218 14872 11290
rect 15028 11218 15056 12543
rect 15212 11830 15240 12582
rect 16224 12434 16252 13330
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16302 12880 16358 12889
rect 16302 12815 16358 12824
rect 16316 12782 16344 12815
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16776 12646 16804 13194
rect 17040 13184 17092 13190
rect 17040 13126 17092 13132
rect 17052 12782 17080 13126
rect 17236 12850 17264 13874
rect 18340 13870 18368 14758
rect 18800 14346 18828 15030
rect 18984 14550 19012 17138
rect 19076 15570 19104 18788
rect 19248 18770 19300 18776
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19904 18426 19932 18566
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19628 17882 19656 18022
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 19352 15570 19380 17206
rect 20180 16998 20208 19314
rect 20364 17134 20392 21422
rect 20548 20398 20576 22034
rect 20720 21548 20772 21554
rect 20720 21490 20772 21496
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20456 18766 20484 19110
rect 20548 18834 20576 20334
rect 20732 19446 20760 21490
rect 20824 21146 20852 22714
rect 20996 22568 21048 22574
rect 20996 22510 21048 22516
rect 21008 22234 21036 22510
rect 20996 22228 21048 22234
rect 20996 22170 21048 22176
rect 21100 22137 21128 24550
rect 21304 24508 21612 24517
rect 21304 24506 21310 24508
rect 21366 24506 21390 24508
rect 21446 24506 21470 24508
rect 21526 24506 21550 24508
rect 21606 24506 21612 24508
rect 21366 24454 21368 24506
rect 21548 24454 21550 24506
rect 21304 24452 21310 24454
rect 21366 24452 21390 24454
rect 21446 24452 21470 24454
rect 21526 24452 21550 24454
rect 21606 24452 21612 24454
rect 21304 24443 21612 24452
rect 21640 24268 21692 24274
rect 21640 24210 21692 24216
rect 21652 23730 21680 24210
rect 21836 24138 21864 24686
rect 22020 24188 22048 24754
rect 22664 24732 22692 24890
rect 22572 24704 22692 24732
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 22192 24200 22244 24206
rect 21928 24160 22192 24188
rect 21824 24132 21876 24138
rect 21824 24074 21876 24080
rect 21640 23724 21692 23730
rect 21640 23666 21692 23672
rect 21304 23420 21612 23429
rect 21304 23418 21310 23420
rect 21366 23418 21390 23420
rect 21446 23418 21470 23420
rect 21526 23418 21550 23420
rect 21606 23418 21612 23420
rect 21366 23366 21368 23418
rect 21548 23366 21550 23418
rect 21304 23364 21310 23366
rect 21366 23364 21390 23366
rect 21446 23364 21470 23366
rect 21526 23364 21550 23366
rect 21606 23364 21612 23366
rect 21304 23355 21612 23364
rect 21652 23322 21680 23666
rect 21928 23662 21956 24160
rect 22192 24142 22244 24148
rect 22480 24154 22508 24346
rect 22572 24274 22600 24704
rect 22652 24608 22704 24614
rect 22652 24550 22704 24556
rect 22664 24410 22692 24550
rect 22652 24404 22704 24410
rect 22652 24346 22704 24352
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22480 24126 22692 24154
rect 22468 24064 22520 24070
rect 22468 24006 22520 24012
rect 22480 23730 22508 24006
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 21916 23656 21968 23662
rect 21916 23598 21968 23604
rect 22376 23656 22428 23662
rect 22376 23598 22428 23604
rect 21640 23316 21692 23322
rect 21640 23258 21692 23264
rect 21928 23254 21956 23598
rect 21916 23248 21968 23254
rect 21916 23190 21968 23196
rect 21732 23044 21784 23050
rect 21732 22986 21784 22992
rect 21180 22704 21232 22710
rect 21180 22646 21232 22652
rect 21086 22128 21142 22137
rect 21086 22063 21142 22072
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 21008 21486 21036 21966
rect 21100 21690 21128 22063
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 21008 20890 21036 21422
rect 20824 20862 21036 20890
rect 20720 19440 20772 19446
rect 20720 19382 20772 19388
rect 20824 18902 20852 20862
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20916 20602 20944 20742
rect 21192 20602 21220 22646
rect 21640 22432 21692 22438
rect 21640 22374 21692 22380
rect 21304 22332 21612 22341
rect 21304 22330 21310 22332
rect 21366 22330 21390 22332
rect 21446 22330 21470 22332
rect 21526 22330 21550 22332
rect 21606 22330 21612 22332
rect 21366 22278 21368 22330
rect 21548 22278 21550 22330
rect 21304 22276 21310 22278
rect 21366 22276 21390 22278
rect 21446 22276 21470 22278
rect 21526 22276 21550 22278
rect 21606 22276 21612 22278
rect 21304 22267 21612 22276
rect 21652 21962 21680 22374
rect 21744 22166 21772 22986
rect 21824 22976 21876 22982
rect 21824 22918 21876 22924
rect 21732 22160 21784 22166
rect 21732 22102 21784 22108
rect 21640 21956 21692 21962
rect 21640 21898 21692 21904
rect 21652 21486 21680 21898
rect 21744 21894 21772 22102
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 21304 21244 21612 21253
rect 21304 21242 21310 21244
rect 21366 21242 21390 21244
rect 21446 21242 21470 21244
rect 21526 21242 21550 21244
rect 21606 21242 21612 21244
rect 21366 21190 21368 21242
rect 21548 21190 21550 21242
rect 21304 21188 21310 21190
rect 21366 21188 21390 21190
rect 21446 21188 21470 21190
rect 21526 21188 21550 21190
rect 21606 21188 21612 21190
rect 21304 21179 21612 21188
rect 21732 21072 21784 21078
rect 21732 21014 21784 21020
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 21008 20058 21036 20334
rect 20996 20052 21048 20058
rect 20996 19994 21048 20000
rect 21008 19310 21036 19994
rect 21192 19922 21220 20538
rect 21744 20398 21772 21014
rect 21836 21010 21864 22918
rect 22388 22778 22416 23598
rect 22664 23526 22692 24126
rect 22560 23520 22612 23526
rect 22560 23462 22612 23468
rect 22652 23520 22704 23526
rect 22652 23462 22704 23468
rect 22376 22772 22428 22778
rect 22376 22714 22428 22720
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 22112 22166 22140 22374
rect 22100 22160 22152 22166
rect 22100 22102 22152 22108
rect 22204 21486 22232 22578
rect 22572 22574 22600 23462
rect 22664 22794 22692 23462
rect 22940 23225 22968 25094
rect 23216 24274 23244 25230
rect 23204 24268 23256 24274
rect 23572 24268 23624 24274
rect 23256 24228 23336 24256
rect 23204 24210 23256 24216
rect 23112 24132 23164 24138
rect 23112 24074 23164 24080
rect 22926 23216 22982 23225
rect 22926 23151 22982 23160
rect 22664 22766 22784 22794
rect 22652 22636 22704 22642
rect 22652 22578 22704 22584
rect 22560 22568 22612 22574
rect 22560 22510 22612 22516
rect 22284 22432 22336 22438
rect 22284 22374 22336 22380
rect 22296 22166 22324 22374
rect 22572 22234 22600 22510
rect 22560 22228 22612 22234
rect 22560 22170 22612 22176
rect 22284 22160 22336 22166
rect 22284 22102 22336 22108
rect 22296 21622 22324 22102
rect 22664 22098 22692 22578
rect 22652 22092 22704 22098
rect 22652 22034 22704 22040
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 21916 21344 21968 21350
rect 21916 21286 21968 21292
rect 21824 21004 21876 21010
rect 21824 20946 21876 20952
rect 21836 20602 21864 20946
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21928 20482 21956 21286
rect 22480 20874 22508 21966
rect 22664 21554 22692 22034
rect 22756 21690 22784 22766
rect 23124 22506 23152 24074
rect 23204 24064 23256 24070
rect 23204 24006 23256 24012
rect 23216 23662 23244 24006
rect 23204 23656 23256 23662
rect 23204 23598 23256 23604
rect 23308 22642 23336 24228
rect 23572 24210 23624 24216
rect 23584 23866 23612 24210
rect 23572 23860 23624 23866
rect 23572 23802 23624 23808
rect 23388 23656 23440 23662
rect 23388 23598 23440 23604
rect 23296 22636 23348 22642
rect 23296 22578 23348 22584
rect 23112 22500 23164 22506
rect 23112 22442 23164 22448
rect 22928 22092 22980 22098
rect 22928 22034 22980 22040
rect 22940 21894 22968 22034
rect 22928 21888 22980 21894
rect 22928 21830 22980 21836
rect 22744 21684 22796 21690
rect 22744 21626 22796 21632
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 22756 21146 22784 21626
rect 22744 21140 22796 21146
rect 22744 21082 22796 21088
rect 22848 21078 22876 21626
rect 22940 21554 22968 21830
rect 22928 21548 22980 21554
rect 22928 21490 22980 21496
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 22836 21072 22888 21078
rect 22836 21014 22888 21020
rect 23032 21010 23060 21286
rect 23020 21004 23072 21010
rect 23020 20946 23072 20952
rect 22468 20868 22520 20874
rect 22468 20810 22520 20816
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22204 20602 22232 20742
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 21836 20454 21956 20482
rect 21732 20392 21784 20398
rect 21732 20334 21784 20340
rect 21640 20256 21692 20262
rect 21640 20198 21692 20204
rect 21304 20156 21612 20165
rect 21304 20154 21310 20156
rect 21366 20154 21390 20156
rect 21446 20154 21470 20156
rect 21526 20154 21550 20156
rect 21606 20154 21612 20156
rect 21366 20102 21368 20154
rect 21548 20102 21550 20154
rect 21304 20100 21310 20102
rect 21366 20100 21390 20102
rect 21446 20100 21470 20102
rect 21526 20100 21550 20102
rect 21606 20100 21612 20102
rect 21304 20091 21612 20100
rect 21652 19922 21680 20198
rect 21180 19916 21232 19922
rect 21180 19858 21232 19864
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 20996 19304 21048 19310
rect 20996 19246 21048 19252
rect 21192 19174 21220 19858
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21284 19514 21312 19654
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21548 19304 21600 19310
rect 21546 19272 21548 19281
rect 21600 19272 21602 19281
rect 21546 19207 21602 19216
rect 21836 19224 21864 20454
rect 22480 20398 22508 20810
rect 22100 20392 22152 20398
rect 22100 20334 22152 20340
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22112 20058 22140 20334
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 21916 19984 21968 19990
rect 21916 19926 21968 19932
rect 21928 19334 21956 19926
rect 22112 19514 22140 19994
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 21928 19310 22140 19334
rect 22296 19310 22324 19858
rect 21928 19306 22152 19310
rect 22100 19304 22152 19306
rect 22100 19246 22152 19252
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 21916 19236 21968 19242
rect 21836 19196 21916 19224
rect 21916 19178 21968 19184
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21640 19168 21692 19174
rect 21640 19110 21692 19116
rect 21304 19068 21612 19077
rect 21304 19066 21310 19068
rect 21366 19066 21390 19068
rect 21446 19066 21470 19068
rect 21526 19066 21550 19068
rect 21606 19066 21612 19068
rect 21366 19014 21368 19066
rect 21548 19014 21550 19066
rect 21304 19012 21310 19014
rect 21366 19012 21390 19014
rect 21446 19012 21470 19014
rect 21526 19012 21550 19014
rect 21606 19012 21612 19014
rect 21304 19003 21612 19012
rect 21652 18970 21680 19110
rect 21640 18964 21692 18970
rect 21640 18906 21692 18912
rect 20812 18896 20864 18902
rect 20812 18838 20864 18844
rect 20536 18828 20588 18834
rect 20536 18770 20588 18776
rect 21928 18766 21956 19178
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 21916 18760 21968 18766
rect 21916 18702 21968 18708
rect 20536 18692 20588 18698
rect 20536 18634 20588 18640
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20180 16658 20208 16934
rect 19892 16652 19944 16658
rect 19892 16594 19944 16600
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19064 15360 19116 15366
rect 19064 15302 19116 15308
rect 18972 14544 19024 14550
rect 18972 14486 19024 14492
rect 18788 14340 18840 14346
rect 18788 14282 18840 14288
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18800 13462 18828 14282
rect 18984 13938 19012 14486
rect 19076 14482 19104 15302
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 18880 13728 18932 13734
rect 18880 13670 18932 13676
rect 17684 13456 17736 13462
rect 17684 13398 17736 13404
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 17696 12986 17724 13398
rect 18052 13320 18104 13326
rect 18604 13320 18656 13326
rect 18104 13268 18184 13274
rect 18052 13262 18184 13268
rect 18604 13262 18656 13268
rect 18064 13246 18184 13262
rect 17820 13084 18128 13093
rect 17820 13082 17826 13084
rect 17882 13082 17906 13084
rect 17962 13082 17986 13084
rect 18042 13082 18066 13084
rect 18122 13082 18128 13084
rect 17882 13030 17884 13082
rect 18064 13030 18066 13082
rect 17820 13028 17826 13030
rect 17882 13028 17906 13030
rect 17962 13028 17986 13030
rect 18042 13028 18066 13030
rect 18122 13028 18128 13030
rect 17820 13019 18128 13028
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 17236 12646 17264 12786
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 16132 12406 16252 12434
rect 16132 12374 16160 12406
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15304 11354 15332 11562
rect 15396 11558 15424 11630
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15396 11286 15424 11494
rect 15580 11354 15608 11494
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15384 11280 15436 11286
rect 15384 11222 15436 11228
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 11808 10810 11836 11154
rect 14844 11082 14872 11154
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 16132 11014 16160 12310
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 11354 16252 11494
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16408 11286 16436 12038
rect 16396 11280 16448 11286
rect 16396 11222 16448 11228
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 16592 10674 16620 10950
rect 16868 10810 16896 11086
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 17604 10606 17632 12854
rect 17820 11996 18128 12005
rect 17820 11994 17826 11996
rect 17882 11994 17906 11996
rect 17962 11994 17986 11996
rect 18042 11994 18066 11996
rect 18122 11994 18128 11996
rect 17882 11942 17884 11994
rect 18064 11942 18066 11994
rect 17820 11940 17826 11942
rect 17882 11940 17906 11942
rect 17962 11940 17986 11942
rect 18042 11940 18066 11942
rect 18122 11940 18128 11942
rect 17820 11931 18128 11940
rect 18156 11898 18184 13246
rect 18616 12306 18644 13262
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18156 11218 18184 11834
rect 18800 11694 18828 13398
rect 18892 13326 18920 13670
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18984 13258 19012 13874
rect 19076 13870 19104 14418
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19352 14074 19380 14214
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19444 13954 19472 16526
rect 19904 15570 19932 16594
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 20088 15706 20116 16390
rect 20548 16182 20576 18634
rect 20732 17882 20760 18702
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 21304 17980 21612 17989
rect 21304 17978 21310 17980
rect 21366 17978 21390 17980
rect 21446 17978 21470 17980
rect 21526 17978 21550 17980
rect 21606 17978 21612 17980
rect 21366 17926 21368 17978
rect 21548 17926 21550 17978
rect 21304 17924 21310 17926
rect 21366 17924 21390 17926
rect 21446 17924 21470 17926
rect 21526 17924 21550 17926
rect 21606 17924 21612 17926
rect 21304 17915 21612 17924
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 21304 16892 21612 16901
rect 21304 16890 21310 16892
rect 21366 16890 21390 16892
rect 21446 16890 21470 16892
rect 21526 16890 21550 16892
rect 21606 16890 21612 16892
rect 21366 16838 21368 16890
rect 21548 16838 21550 16890
rect 21304 16836 21310 16838
rect 21366 16836 21390 16838
rect 21446 16836 21470 16838
rect 21526 16836 21550 16838
rect 21606 16836 21612 16838
rect 21304 16827 21612 16836
rect 20536 16176 20588 16182
rect 20536 16118 20588 16124
rect 20168 15972 20220 15978
rect 20168 15914 20220 15920
rect 20180 15706 20208 15914
rect 20548 15706 20576 16118
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 21304 15804 21612 15813
rect 21304 15802 21310 15804
rect 21366 15802 21390 15804
rect 21446 15802 21470 15804
rect 21526 15802 21550 15804
rect 21606 15802 21612 15804
rect 21366 15750 21368 15802
rect 21548 15750 21550 15802
rect 21304 15748 21310 15750
rect 21366 15748 21390 15750
rect 21446 15748 21470 15750
rect 21526 15748 21550 15750
rect 21606 15748 21612 15750
rect 21304 15739 21612 15748
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 20168 15700 20220 15706
rect 20168 15642 20220 15648
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 19892 15564 19944 15570
rect 19892 15506 19944 15512
rect 19984 15564 20036 15570
rect 19984 15506 20036 15512
rect 19996 15162 20024 15506
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 20272 15094 20300 15302
rect 20260 15088 20312 15094
rect 20260 15030 20312 15036
rect 19352 13926 19472 13954
rect 19064 13864 19116 13870
rect 19116 13812 19196 13818
rect 19064 13806 19196 13812
rect 19076 13790 19196 13806
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 19168 12306 19196 13790
rect 19352 13530 19380 13926
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19444 13734 19472 13806
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19444 13394 19472 13670
rect 19536 13530 19564 13806
rect 19904 13530 19932 13806
rect 20272 13734 20300 15030
rect 20364 13870 20392 15302
rect 20444 14952 20496 14958
rect 20548 14940 20576 15642
rect 20996 15632 21048 15638
rect 20996 15574 21048 15580
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20640 15026 20668 15506
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 21008 14958 21036 15574
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21284 15162 21312 15506
rect 21640 15360 21692 15366
rect 21640 15302 21692 15308
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 20496 14912 20576 14940
rect 20996 14952 21048 14958
rect 20444 14894 20496 14900
rect 20996 14894 21048 14900
rect 21652 14890 21680 15302
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 20628 14884 20680 14890
rect 20628 14826 20680 14832
rect 21640 14884 21692 14890
rect 21640 14826 21692 14832
rect 20640 13870 20668 14826
rect 21304 14716 21612 14725
rect 21304 14714 21310 14716
rect 21366 14714 21390 14716
rect 21446 14714 21470 14716
rect 21526 14714 21550 14716
rect 21606 14714 21612 14716
rect 21366 14662 21368 14714
rect 21548 14662 21550 14714
rect 21304 14660 21310 14662
rect 21366 14660 21390 14662
rect 21446 14660 21470 14662
rect 21526 14660 21550 14662
rect 21606 14660 21612 14662
rect 21304 14651 21612 14660
rect 21640 14476 21692 14482
rect 21640 14418 21692 14424
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19892 13524 19944 13530
rect 19892 13466 19944 13472
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19616 13184 19668 13190
rect 19616 13126 19668 13132
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19168 11762 19196 12242
rect 19260 11830 19288 12242
rect 19628 12170 19656 13126
rect 19996 12918 20024 13670
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 19708 12708 19760 12714
rect 19708 12650 19760 12656
rect 19720 12306 19748 12650
rect 19996 12306 20024 12854
rect 20364 12646 20392 13262
rect 20640 12714 20668 13806
rect 21088 13728 21140 13734
rect 21088 13670 21140 13676
rect 21100 13530 21128 13670
rect 21304 13628 21612 13637
rect 21304 13626 21310 13628
rect 21366 13626 21390 13628
rect 21446 13626 21470 13628
rect 21526 13626 21550 13628
rect 21606 13626 21612 13628
rect 21366 13574 21368 13626
rect 21548 13574 21550 13626
rect 21304 13572 21310 13574
rect 21366 13572 21390 13574
rect 21446 13572 21470 13574
rect 21526 13572 21550 13574
rect 21606 13572 21612 13574
rect 21304 13563 21612 13572
rect 21652 13530 21680 14418
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21928 13326 21956 14894
rect 22112 13818 22140 16050
rect 22204 14958 22232 18566
rect 22480 15638 22508 20334
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22848 19310 22876 20198
rect 23032 20058 23060 20946
rect 23020 20052 23072 20058
rect 23020 19994 23072 20000
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 22928 19848 22980 19854
rect 22928 19790 22980 19796
rect 22560 19304 22612 19310
rect 22560 19246 22612 19252
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 22572 18630 22600 19246
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 22940 16114 22968 19790
rect 23216 19514 23244 19858
rect 23204 19508 23256 19514
rect 23204 19450 23256 19456
rect 23308 18902 23336 22578
rect 23400 22114 23428 23598
rect 23480 22568 23532 22574
rect 23480 22510 23532 22516
rect 23492 22386 23520 22510
rect 23664 22432 23716 22438
rect 23492 22358 23612 22386
rect 23664 22374 23716 22380
rect 23478 22128 23534 22137
rect 23400 22086 23478 22114
rect 23478 22063 23480 22072
rect 23532 22063 23534 22072
rect 23480 22034 23532 22040
rect 23388 20800 23440 20806
rect 23388 20742 23440 20748
rect 23400 20602 23428 20742
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23492 20398 23520 22034
rect 23584 21962 23612 22358
rect 23676 22234 23704 22374
rect 23664 22228 23716 22234
rect 23664 22170 23716 22176
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23296 18896 23348 18902
rect 23296 18838 23348 18844
rect 23308 17270 23336 18838
rect 23768 18834 23796 26794
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 23848 25832 23900 25838
rect 23848 25774 23900 25780
rect 23860 25430 23888 25774
rect 23848 25424 23900 25430
rect 23848 25366 23900 25372
rect 23860 24206 23888 25366
rect 24228 25362 24256 26726
rect 24789 26140 25097 26149
rect 24789 26138 24795 26140
rect 24851 26138 24875 26140
rect 24931 26138 24955 26140
rect 25011 26138 25035 26140
rect 25091 26138 25097 26140
rect 24851 26086 24853 26138
rect 25033 26086 25035 26138
rect 24789 26084 24795 26086
rect 24851 26084 24875 26086
rect 24931 26084 24955 26086
rect 25011 26084 25035 26086
rect 25091 26084 25097 26086
rect 24789 26075 25097 26084
rect 24216 25356 24268 25362
rect 24216 25298 24268 25304
rect 24789 25052 25097 25061
rect 24789 25050 24795 25052
rect 24851 25050 24875 25052
rect 24931 25050 24955 25052
rect 25011 25050 25035 25052
rect 25091 25050 25097 25052
rect 24851 24998 24853 25050
rect 25033 24998 25035 25050
rect 24789 24996 24795 24998
rect 24851 24996 24875 24998
rect 24931 24996 24955 24998
rect 25011 24996 25035 24998
rect 25091 24996 25097 24998
rect 24789 24987 25097 24996
rect 24492 24268 24544 24274
rect 24492 24210 24544 24216
rect 23848 24200 23900 24206
rect 23848 24142 23900 24148
rect 23860 22642 23888 24142
rect 24216 24064 24268 24070
rect 24216 24006 24268 24012
rect 24228 23866 24256 24006
rect 24504 23866 24532 24210
rect 24584 24064 24636 24070
rect 24584 24006 24636 24012
rect 24216 23860 24268 23866
rect 24216 23802 24268 23808
rect 24492 23860 24544 23866
rect 24492 23802 24544 23808
rect 24596 23662 24624 24006
rect 24789 23964 25097 23973
rect 24789 23962 24795 23964
rect 24851 23962 24875 23964
rect 24931 23962 24955 23964
rect 25011 23962 25035 23964
rect 25091 23962 25097 23964
rect 24851 23910 24853 23962
rect 25033 23910 25035 23962
rect 24789 23908 24795 23910
rect 24851 23908 24875 23910
rect 24931 23908 24955 23910
rect 25011 23908 25035 23910
rect 25091 23908 25097 23910
rect 24789 23899 25097 23908
rect 24400 23656 24452 23662
rect 24400 23598 24452 23604
rect 24584 23656 24636 23662
rect 24584 23598 24636 23604
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 24308 22500 24360 22506
rect 24308 22442 24360 22448
rect 24320 22234 24348 22442
rect 24308 22228 24360 22234
rect 24308 22170 24360 22176
rect 24308 21548 24360 21554
rect 24308 21490 24360 21496
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 23860 21146 23888 21286
rect 23848 21140 23900 21146
rect 23848 21082 23900 21088
rect 24320 20058 24348 21490
rect 24412 20874 24440 23598
rect 24789 22876 25097 22885
rect 24789 22874 24795 22876
rect 24851 22874 24875 22876
rect 24931 22874 24955 22876
rect 25011 22874 25035 22876
rect 25091 22874 25097 22876
rect 24851 22822 24853 22874
rect 25033 22822 25035 22874
rect 24789 22820 24795 22822
rect 24851 22820 24875 22822
rect 24931 22820 24955 22822
rect 25011 22820 25035 22822
rect 25091 22820 25097 22822
rect 24789 22811 25097 22820
rect 25228 22432 25280 22438
rect 25228 22374 25280 22380
rect 24789 21788 25097 21797
rect 24789 21786 24795 21788
rect 24851 21786 24875 21788
rect 24931 21786 24955 21788
rect 25011 21786 25035 21788
rect 25091 21786 25097 21788
rect 24851 21734 24853 21786
rect 25033 21734 25035 21786
rect 24789 21732 24795 21734
rect 24851 21732 24875 21734
rect 24931 21732 24955 21734
rect 25011 21732 25035 21734
rect 25091 21732 25097 21734
rect 24789 21723 25097 21732
rect 25240 21486 25268 22374
rect 25228 21480 25280 21486
rect 25228 21422 25280 21428
rect 24400 20868 24452 20874
rect 24400 20810 24452 20816
rect 24789 20700 25097 20709
rect 24789 20698 24795 20700
rect 24851 20698 24875 20700
rect 24931 20698 24955 20700
rect 25011 20698 25035 20700
rect 25091 20698 25097 20700
rect 24851 20646 24853 20698
rect 25033 20646 25035 20698
rect 24789 20644 24795 20646
rect 24851 20644 24875 20646
rect 24931 20644 24955 20646
rect 25011 20644 25035 20646
rect 25091 20644 25097 20646
rect 24789 20635 25097 20644
rect 24308 20052 24360 20058
rect 24308 19994 24360 20000
rect 24789 19612 25097 19621
rect 24789 19610 24795 19612
rect 24851 19610 24875 19612
rect 24931 19610 24955 19612
rect 25011 19610 25035 19612
rect 25091 19610 25097 19612
rect 24851 19558 24853 19610
rect 25033 19558 25035 19610
rect 24789 19556 24795 19558
rect 24851 19556 24875 19558
rect 24931 19556 24955 19558
rect 25011 19556 25035 19558
rect 25091 19556 25097 19558
rect 24789 19547 25097 19556
rect 27632 19281 27660 28600
rect 28273 27772 28581 27781
rect 28273 27770 28279 27772
rect 28335 27770 28359 27772
rect 28415 27770 28439 27772
rect 28495 27770 28519 27772
rect 28575 27770 28581 27772
rect 28335 27718 28337 27770
rect 28517 27718 28519 27770
rect 28273 27716 28279 27718
rect 28335 27716 28359 27718
rect 28415 27716 28439 27718
rect 28495 27716 28519 27718
rect 28575 27716 28581 27718
rect 28273 27707 28581 27716
rect 28273 26684 28581 26693
rect 28273 26682 28279 26684
rect 28335 26682 28359 26684
rect 28415 26682 28439 26684
rect 28495 26682 28519 26684
rect 28575 26682 28581 26684
rect 28335 26630 28337 26682
rect 28517 26630 28519 26682
rect 28273 26628 28279 26630
rect 28335 26628 28359 26630
rect 28415 26628 28439 26630
rect 28495 26628 28519 26630
rect 28575 26628 28581 26630
rect 28273 26619 28581 26628
rect 28273 25596 28581 25605
rect 28273 25594 28279 25596
rect 28335 25594 28359 25596
rect 28415 25594 28439 25596
rect 28495 25594 28519 25596
rect 28575 25594 28581 25596
rect 28335 25542 28337 25594
rect 28517 25542 28519 25594
rect 28273 25540 28279 25542
rect 28335 25540 28359 25542
rect 28415 25540 28439 25542
rect 28495 25540 28519 25542
rect 28575 25540 28581 25542
rect 28273 25531 28581 25540
rect 28273 24508 28581 24517
rect 28273 24506 28279 24508
rect 28335 24506 28359 24508
rect 28415 24506 28439 24508
rect 28495 24506 28519 24508
rect 28575 24506 28581 24508
rect 28335 24454 28337 24506
rect 28517 24454 28519 24506
rect 28273 24452 28279 24454
rect 28335 24452 28359 24454
rect 28415 24452 28439 24454
rect 28495 24452 28519 24454
rect 28575 24452 28581 24454
rect 28273 24443 28581 24452
rect 28273 23420 28581 23429
rect 28273 23418 28279 23420
rect 28335 23418 28359 23420
rect 28415 23418 28439 23420
rect 28495 23418 28519 23420
rect 28575 23418 28581 23420
rect 28335 23366 28337 23418
rect 28517 23366 28519 23418
rect 28273 23364 28279 23366
rect 28335 23364 28359 23366
rect 28415 23364 28439 23366
rect 28495 23364 28519 23366
rect 28575 23364 28581 23366
rect 28273 23355 28581 23364
rect 28273 22332 28581 22341
rect 28273 22330 28279 22332
rect 28335 22330 28359 22332
rect 28415 22330 28439 22332
rect 28495 22330 28519 22332
rect 28575 22330 28581 22332
rect 28335 22278 28337 22330
rect 28517 22278 28519 22330
rect 28273 22276 28279 22278
rect 28335 22276 28359 22278
rect 28415 22276 28439 22278
rect 28495 22276 28519 22278
rect 28575 22276 28581 22278
rect 28273 22267 28581 22276
rect 28273 21244 28581 21253
rect 28273 21242 28279 21244
rect 28335 21242 28359 21244
rect 28415 21242 28439 21244
rect 28495 21242 28519 21244
rect 28575 21242 28581 21244
rect 28335 21190 28337 21242
rect 28517 21190 28519 21242
rect 28273 21188 28279 21190
rect 28335 21188 28359 21190
rect 28415 21188 28439 21190
rect 28495 21188 28519 21190
rect 28575 21188 28581 21190
rect 28273 21179 28581 21188
rect 28273 20156 28581 20165
rect 28273 20154 28279 20156
rect 28335 20154 28359 20156
rect 28415 20154 28439 20156
rect 28495 20154 28519 20156
rect 28575 20154 28581 20156
rect 28335 20102 28337 20154
rect 28517 20102 28519 20154
rect 28273 20100 28279 20102
rect 28335 20100 28359 20102
rect 28415 20100 28439 20102
rect 28495 20100 28519 20102
rect 28575 20100 28581 20102
rect 28273 20091 28581 20100
rect 27618 19272 27674 19281
rect 27618 19207 27674 19216
rect 28273 19068 28581 19077
rect 28273 19066 28279 19068
rect 28335 19066 28359 19068
rect 28415 19066 28439 19068
rect 28495 19066 28519 19068
rect 28575 19066 28581 19068
rect 28335 19014 28337 19066
rect 28517 19014 28519 19066
rect 28273 19012 28279 19014
rect 28335 19012 28359 19014
rect 28415 19012 28439 19014
rect 28495 19012 28519 19014
rect 28575 19012 28581 19014
rect 28273 19003 28581 19012
rect 23756 18828 23808 18834
rect 23756 18770 23808 18776
rect 24789 18524 25097 18533
rect 24789 18522 24795 18524
rect 24851 18522 24875 18524
rect 24931 18522 24955 18524
rect 25011 18522 25035 18524
rect 25091 18522 25097 18524
rect 24851 18470 24853 18522
rect 25033 18470 25035 18522
rect 24789 18468 24795 18470
rect 24851 18468 24875 18470
rect 24931 18468 24955 18470
rect 25011 18468 25035 18470
rect 25091 18468 25097 18470
rect 24789 18459 25097 18468
rect 28273 17980 28581 17989
rect 28273 17978 28279 17980
rect 28335 17978 28359 17980
rect 28415 17978 28439 17980
rect 28495 17978 28519 17980
rect 28575 17978 28581 17980
rect 28335 17926 28337 17978
rect 28517 17926 28519 17978
rect 28273 17924 28279 17926
rect 28335 17924 28359 17926
rect 28415 17924 28439 17926
rect 28495 17924 28519 17926
rect 28575 17924 28581 17926
rect 28273 17915 28581 17924
rect 24789 17436 25097 17445
rect 24789 17434 24795 17436
rect 24851 17434 24875 17436
rect 24931 17434 24955 17436
rect 25011 17434 25035 17436
rect 25091 17434 25097 17436
rect 24851 17382 24853 17434
rect 25033 17382 25035 17434
rect 24789 17380 24795 17382
rect 24851 17380 24875 17382
rect 24931 17380 24955 17382
rect 25011 17380 25035 17382
rect 25091 17380 25097 17382
rect 24789 17371 25097 17380
rect 23296 17264 23348 17270
rect 23296 17206 23348 17212
rect 28273 16892 28581 16901
rect 28273 16890 28279 16892
rect 28335 16890 28359 16892
rect 28415 16890 28439 16892
rect 28495 16890 28519 16892
rect 28575 16890 28581 16892
rect 28335 16838 28337 16890
rect 28517 16838 28519 16890
rect 28273 16836 28279 16838
rect 28335 16836 28359 16838
rect 28415 16836 28439 16838
rect 28495 16836 28519 16838
rect 28575 16836 28581 16838
rect 28273 16827 28581 16836
rect 24789 16348 25097 16357
rect 24789 16346 24795 16348
rect 24851 16346 24875 16348
rect 24931 16346 24955 16348
rect 25011 16346 25035 16348
rect 25091 16346 25097 16348
rect 24851 16294 24853 16346
rect 25033 16294 25035 16346
rect 24789 16292 24795 16294
rect 24851 16292 24875 16294
rect 24931 16292 24955 16294
rect 25011 16292 25035 16294
rect 25091 16292 25097 16294
rect 24789 16283 25097 16292
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 22468 15632 22520 15638
rect 22468 15574 22520 15580
rect 22940 15570 22968 16050
rect 28273 15804 28581 15813
rect 28273 15802 28279 15804
rect 28335 15802 28359 15804
rect 28415 15802 28439 15804
rect 28495 15802 28519 15804
rect 28575 15802 28581 15804
rect 28335 15750 28337 15802
rect 28517 15750 28519 15802
rect 28273 15748 28279 15750
rect 28335 15748 28359 15750
rect 28415 15748 28439 15750
rect 28495 15748 28519 15750
rect 28575 15748 28581 15750
rect 28273 15739 28581 15748
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 24789 15260 25097 15269
rect 24789 15258 24795 15260
rect 24851 15258 24875 15260
rect 24931 15258 24955 15260
rect 25011 15258 25035 15260
rect 25091 15258 25097 15260
rect 24851 15206 24853 15258
rect 25033 15206 25035 15258
rect 24789 15204 24795 15206
rect 24851 15204 24875 15206
rect 24931 15204 24955 15206
rect 25011 15204 25035 15206
rect 25091 15204 25097 15206
rect 24789 15195 25097 15204
rect 22192 14952 22244 14958
rect 22192 14894 22244 14900
rect 28273 14716 28581 14725
rect 28273 14714 28279 14716
rect 28335 14714 28359 14716
rect 28415 14714 28439 14716
rect 28495 14714 28519 14716
rect 28575 14714 28581 14716
rect 28335 14662 28337 14714
rect 28517 14662 28519 14714
rect 28273 14660 28279 14662
rect 28335 14660 28359 14662
rect 28415 14660 28439 14662
rect 28495 14660 28519 14662
rect 28575 14660 28581 14662
rect 28273 14651 28581 14660
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22020 13802 22140 13818
rect 22296 13802 22324 14214
rect 24789 14172 25097 14181
rect 24789 14170 24795 14172
rect 24851 14170 24875 14172
rect 24931 14170 24955 14172
rect 25011 14170 25035 14172
rect 25091 14170 25097 14172
rect 24851 14118 24853 14170
rect 25033 14118 25035 14170
rect 24789 14116 24795 14118
rect 24851 14116 24875 14118
rect 24931 14116 24955 14118
rect 25011 14116 25035 14118
rect 25091 14116 25097 14118
rect 24789 14107 25097 14116
rect 22008 13796 22140 13802
rect 22060 13790 22140 13796
rect 22284 13796 22336 13802
rect 22008 13738 22060 13744
rect 22284 13738 22336 13744
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 20628 12708 20680 12714
rect 20628 12650 20680 12656
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20364 12306 20392 12582
rect 21304 12540 21612 12549
rect 21304 12538 21310 12540
rect 21366 12538 21390 12540
rect 21446 12538 21470 12540
rect 21526 12538 21550 12540
rect 21606 12538 21612 12540
rect 21366 12486 21368 12538
rect 21548 12486 21550 12538
rect 21304 12484 21310 12486
rect 21366 12484 21390 12486
rect 21446 12484 21470 12486
rect 21526 12484 21550 12486
rect 21606 12484 21612 12486
rect 21304 12475 21612 12484
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 20352 12300 20404 12306
rect 20352 12242 20404 12248
rect 19616 12164 19668 12170
rect 19616 12106 19668 12112
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 19248 11824 19300 11830
rect 19248 11766 19300 11772
rect 19156 11756 19208 11762
rect 19156 11698 19208 11704
rect 20916 11694 20944 12038
rect 22020 11898 22048 13738
rect 28273 13628 28581 13637
rect 28273 13626 28279 13628
rect 28335 13626 28359 13628
rect 28415 13626 28439 13628
rect 28495 13626 28519 13628
rect 28575 13626 28581 13628
rect 28335 13574 28337 13626
rect 28517 13574 28519 13626
rect 28273 13572 28279 13574
rect 28335 13572 28359 13574
rect 28415 13572 28439 13574
rect 28495 13572 28519 13574
rect 28575 13572 28581 13574
rect 28273 13563 28581 13572
rect 24789 13084 25097 13093
rect 24789 13082 24795 13084
rect 24851 13082 24875 13084
rect 24931 13082 24955 13084
rect 25011 13082 25035 13084
rect 25091 13082 25097 13084
rect 24851 13030 24853 13082
rect 25033 13030 25035 13082
rect 24789 13028 24795 13030
rect 24851 13028 24875 13030
rect 24931 13028 24955 13030
rect 25011 13028 25035 13030
rect 25091 13028 25097 13030
rect 24789 13019 25097 13028
rect 28273 12540 28581 12549
rect 28273 12538 28279 12540
rect 28335 12538 28359 12540
rect 28415 12538 28439 12540
rect 28495 12538 28519 12540
rect 28575 12538 28581 12540
rect 28335 12486 28337 12538
rect 28517 12486 28519 12538
rect 28273 12484 28279 12486
rect 28335 12484 28359 12486
rect 28415 12484 28439 12486
rect 28495 12484 28519 12486
rect 28575 12484 28581 12486
rect 28273 12475 28581 12484
rect 24789 11996 25097 12005
rect 24789 11994 24795 11996
rect 24851 11994 24875 11996
rect 24931 11994 24955 11996
rect 25011 11994 25035 11996
rect 25091 11994 25097 11996
rect 24851 11942 24853 11994
rect 25033 11942 25035 11994
rect 24789 11940 24795 11942
rect 24851 11940 24875 11942
rect 24931 11940 24955 11942
rect 25011 11940 25035 11942
rect 25091 11940 25097 11942
rect 24789 11931 25097 11940
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 21304 11452 21612 11461
rect 21304 11450 21310 11452
rect 21366 11450 21390 11452
rect 21446 11450 21470 11452
rect 21526 11450 21550 11452
rect 21606 11450 21612 11452
rect 21366 11398 21368 11450
rect 21548 11398 21550 11450
rect 21304 11396 21310 11398
rect 21366 11396 21390 11398
rect 21446 11396 21470 11398
rect 21526 11396 21550 11398
rect 21606 11396 21612 11398
rect 21304 11387 21612 11396
rect 28273 11452 28581 11461
rect 28273 11450 28279 11452
rect 28335 11450 28359 11452
rect 28415 11450 28439 11452
rect 28495 11450 28519 11452
rect 28575 11450 28581 11452
rect 28335 11398 28337 11450
rect 28517 11398 28519 11450
rect 28273 11396 28279 11398
rect 28335 11396 28359 11398
rect 28415 11396 28439 11398
rect 28495 11396 28519 11398
rect 28575 11396 28581 11398
rect 28273 11387 28581 11396
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 17820 10908 18128 10917
rect 17820 10906 17826 10908
rect 17882 10906 17906 10908
rect 17962 10906 17986 10908
rect 18042 10906 18066 10908
rect 18122 10906 18128 10908
rect 17882 10854 17884 10906
rect 18064 10854 18066 10906
rect 17820 10852 17826 10854
rect 17882 10852 17906 10854
rect 17962 10852 17986 10854
rect 18042 10852 18066 10854
rect 18122 10852 18128 10854
rect 17820 10843 18128 10852
rect 24789 10908 25097 10917
rect 24789 10906 24795 10908
rect 24851 10906 24875 10908
rect 24931 10906 24955 10908
rect 25011 10906 25035 10908
rect 25091 10906 25097 10908
rect 24851 10854 24853 10906
rect 25033 10854 25035 10906
rect 24789 10852 24795 10854
rect 24851 10852 24875 10854
rect 24931 10852 24955 10854
rect 25011 10852 25035 10854
rect 25091 10852 25097 10854
rect 24789 10843 25097 10852
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 17592 10600 17644 10606
rect 17592 10542 17644 10548
rect 10140 10532 10192 10538
rect 10140 10474 10192 10480
rect 14335 10364 14643 10373
rect 14335 10362 14341 10364
rect 14397 10362 14421 10364
rect 14477 10362 14501 10364
rect 14557 10362 14581 10364
rect 14637 10362 14643 10364
rect 14397 10310 14399 10362
rect 14579 10310 14581 10362
rect 14335 10308 14341 10310
rect 14397 10308 14421 10310
rect 14477 10308 14501 10310
rect 14557 10308 14581 10310
rect 14637 10308 14643 10310
rect 14335 10299 14643 10308
rect 21304 10364 21612 10373
rect 21304 10362 21310 10364
rect 21366 10362 21390 10364
rect 21446 10362 21470 10364
rect 21526 10362 21550 10364
rect 21606 10362 21612 10364
rect 21366 10310 21368 10362
rect 21548 10310 21550 10362
rect 21304 10308 21310 10310
rect 21366 10308 21390 10310
rect 21446 10308 21470 10310
rect 21526 10308 21550 10310
rect 21606 10308 21612 10310
rect 21304 10299 21612 10308
rect 28273 10364 28581 10373
rect 28273 10362 28279 10364
rect 28335 10362 28359 10364
rect 28415 10362 28439 10364
rect 28495 10362 28519 10364
rect 28575 10362 28581 10364
rect 28335 10310 28337 10362
rect 28517 10310 28519 10362
rect 28273 10308 28279 10310
rect 28335 10308 28359 10310
rect 28415 10308 28439 10310
rect 28495 10308 28519 10310
rect 28575 10308 28581 10310
rect 28273 10299 28581 10308
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 3882 9820 4190 9829
rect 3882 9818 3888 9820
rect 3944 9818 3968 9820
rect 4024 9818 4048 9820
rect 4104 9818 4128 9820
rect 4184 9818 4190 9820
rect 3944 9766 3946 9818
rect 4126 9766 4128 9818
rect 3882 9764 3888 9766
rect 3944 9764 3968 9766
rect 4024 9764 4048 9766
rect 4104 9764 4128 9766
rect 4184 9764 4190 9766
rect 3882 9755 4190 9764
rect 10851 9820 11159 9829
rect 10851 9818 10857 9820
rect 10913 9818 10937 9820
rect 10993 9818 11017 9820
rect 11073 9818 11097 9820
rect 11153 9818 11159 9820
rect 10913 9766 10915 9818
rect 11095 9766 11097 9818
rect 10851 9764 10857 9766
rect 10913 9764 10937 9766
rect 10993 9764 11017 9766
rect 11073 9764 11097 9766
rect 11153 9764 11159 9766
rect 10851 9755 11159 9764
rect 17820 9820 18128 9829
rect 17820 9818 17826 9820
rect 17882 9818 17906 9820
rect 17962 9818 17986 9820
rect 18042 9818 18066 9820
rect 18122 9818 18128 9820
rect 17882 9766 17884 9818
rect 18064 9766 18066 9818
rect 17820 9764 17826 9766
rect 17882 9764 17906 9766
rect 17962 9764 17986 9766
rect 18042 9764 18066 9766
rect 18122 9764 18128 9766
rect 17820 9755 18128 9764
rect 24789 9820 25097 9829
rect 24789 9818 24795 9820
rect 24851 9818 24875 9820
rect 24931 9818 24955 9820
rect 25011 9818 25035 9820
rect 25091 9818 25097 9820
rect 24851 9766 24853 9818
rect 25033 9766 25035 9818
rect 24789 9764 24795 9766
rect 24851 9764 24875 9766
rect 24931 9764 24955 9766
rect 25011 9764 25035 9766
rect 25091 9764 25097 9766
rect 24789 9755 25097 9764
rect 7366 9276 7674 9285
rect 7366 9274 7372 9276
rect 7428 9274 7452 9276
rect 7508 9274 7532 9276
rect 7588 9274 7612 9276
rect 7668 9274 7674 9276
rect 7428 9222 7430 9274
rect 7610 9222 7612 9274
rect 7366 9220 7372 9222
rect 7428 9220 7452 9222
rect 7508 9220 7532 9222
rect 7588 9220 7612 9222
rect 7668 9220 7674 9222
rect 7366 9211 7674 9220
rect 14335 9276 14643 9285
rect 14335 9274 14341 9276
rect 14397 9274 14421 9276
rect 14477 9274 14501 9276
rect 14557 9274 14581 9276
rect 14637 9274 14643 9276
rect 14397 9222 14399 9274
rect 14579 9222 14581 9274
rect 14335 9220 14341 9222
rect 14397 9220 14421 9222
rect 14477 9220 14501 9222
rect 14557 9220 14581 9222
rect 14637 9220 14643 9222
rect 14335 9211 14643 9220
rect 21304 9276 21612 9285
rect 21304 9274 21310 9276
rect 21366 9274 21390 9276
rect 21446 9274 21470 9276
rect 21526 9274 21550 9276
rect 21606 9274 21612 9276
rect 21366 9222 21368 9274
rect 21548 9222 21550 9274
rect 21304 9220 21310 9222
rect 21366 9220 21390 9222
rect 21446 9220 21470 9222
rect 21526 9220 21550 9222
rect 21606 9220 21612 9222
rect 21304 9211 21612 9220
rect 28273 9276 28581 9285
rect 28273 9274 28279 9276
rect 28335 9274 28359 9276
rect 28415 9274 28439 9276
rect 28495 9274 28519 9276
rect 28575 9274 28581 9276
rect 28335 9222 28337 9274
rect 28517 9222 28519 9274
rect 28273 9220 28279 9222
rect 28335 9220 28359 9222
rect 28415 9220 28439 9222
rect 28495 9220 28519 9222
rect 28575 9220 28581 9222
rect 28273 9211 28581 9220
rect 3882 8732 4190 8741
rect 3882 8730 3888 8732
rect 3944 8730 3968 8732
rect 4024 8730 4048 8732
rect 4104 8730 4128 8732
rect 4184 8730 4190 8732
rect 3944 8678 3946 8730
rect 4126 8678 4128 8730
rect 3882 8676 3888 8678
rect 3944 8676 3968 8678
rect 4024 8676 4048 8678
rect 4104 8676 4128 8678
rect 4184 8676 4190 8678
rect 3882 8667 4190 8676
rect 10851 8732 11159 8741
rect 10851 8730 10857 8732
rect 10913 8730 10937 8732
rect 10993 8730 11017 8732
rect 11073 8730 11097 8732
rect 11153 8730 11159 8732
rect 10913 8678 10915 8730
rect 11095 8678 11097 8730
rect 10851 8676 10857 8678
rect 10913 8676 10937 8678
rect 10993 8676 11017 8678
rect 11073 8676 11097 8678
rect 11153 8676 11159 8678
rect 10851 8667 11159 8676
rect 17820 8732 18128 8741
rect 17820 8730 17826 8732
rect 17882 8730 17906 8732
rect 17962 8730 17986 8732
rect 18042 8730 18066 8732
rect 18122 8730 18128 8732
rect 17882 8678 17884 8730
rect 18064 8678 18066 8730
rect 17820 8676 17826 8678
rect 17882 8676 17906 8678
rect 17962 8676 17986 8678
rect 18042 8676 18066 8678
rect 18122 8676 18128 8678
rect 17820 8667 18128 8676
rect 24789 8732 25097 8741
rect 24789 8730 24795 8732
rect 24851 8730 24875 8732
rect 24931 8730 24955 8732
rect 25011 8730 25035 8732
rect 25091 8730 25097 8732
rect 24851 8678 24853 8730
rect 25033 8678 25035 8730
rect 24789 8676 24795 8678
rect 24851 8676 24875 8678
rect 24931 8676 24955 8678
rect 25011 8676 25035 8678
rect 25091 8676 25097 8678
rect 24789 8667 25097 8676
rect 7366 8188 7674 8197
rect 7366 8186 7372 8188
rect 7428 8186 7452 8188
rect 7508 8186 7532 8188
rect 7588 8186 7612 8188
rect 7668 8186 7674 8188
rect 7428 8134 7430 8186
rect 7610 8134 7612 8186
rect 7366 8132 7372 8134
rect 7428 8132 7452 8134
rect 7508 8132 7532 8134
rect 7588 8132 7612 8134
rect 7668 8132 7674 8134
rect 7366 8123 7674 8132
rect 14335 8188 14643 8197
rect 14335 8186 14341 8188
rect 14397 8186 14421 8188
rect 14477 8186 14501 8188
rect 14557 8186 14581 8188
rect 14637 8186 14643 8188
rect 14397 8134 14399 8186
rect 14579 8134 14581 8186
rect 14335 8132 14341 8134
rect 14397 8132 14421 8134
rect 14477 8132 14501 8134
rect 14557 8132 14581 8134
rect 14637 8132 14643 8134
rect 14335 8123 14643 8132
rect 21304 8188 21612 8197
rect 21304 8186 21310 8188
rect 21366 8186 21390 8188
rect 21446 8186 21470 8188
rect 21526 8186 21550 8188
rect 21606 8186 21612 8188
rect 21366 8134 21368 8186
rect 21548 8134 21550 8186
rect 21304 8132 21310 8134
rect 21366 8132 21390 8134
rect 21446 8132 21470 8134
rect 21526 8132 21550 8134
rect 21606 8132 21612 8134
rect 21304 8123 21612 8132
rect 28273 8188 28581 8197
rect 28273 8186 28279 8188
rect 28335 8186 28359 8188
rect 28415 8186 28439 8188
rect 28495 8186 28519 8188
rect 28575 8186 28581 8188
rect 28335 8134 28337 8186
rect 28517 8134 28519 8186
rect 28273 8132 28279 8134
rect 28335 8132 28359 8134
rect 28415 8132 28439 8134
rect 28495 8132 28519 8134
rect 28575 8132 28581 8134
rect 28273 8123 28581 8132
rect 3882 7644 4190 7653
rect 3882 7642 3888 7644
rect 3944 7642 3968 7644
rect 4024 7642 4048 7644
rect 4104 7642 4128 7644
rect 4184 7642 4190 7644
rect 3944 7590 3946 7642
rect 4126 7590 4128 7642
rect 3882 7588 3888 7590
rect 3944 7588 3968 7590
rect 4024 7588 4048 7590
rect 4104 7588 4128 7590
rect 4184 7588 4190 7590
rect 3882 7579 4190 7588
rect 10851 7644 11159 7653
rect 10851 7642 10857 7644
rect 10913 7642 10937 7644
rect 10993 7642 11017 7644
rect 11073 7642 11097 7644
rect 11153 7642 11159 7644
rect 10913 7590 10915 7642
rect 11095 7590 11097 7642
rect 10851 7588 10857 7590
rect 10913 7588 10937 7590
rect 10993 7588 11017 7590
rect 11073 7588 11097 7590
rect 11153 7588 11159 7590
rect 10851 7579 11159 7588
rect 17820 7644 18128 7653
rect 17820 7642 17826 7644
rect 17882 7642 17906 7644
rect 17962 7642 17986 7644
rect 18042 7642 18066 7644
rect 18122 7642 18128 7644
rect 17882 7590 17884 7642
rect 18064 7590 18066 7642
rect 17820 7588 17826 7590
rect 17882 7588 17906 7590
rect 17962 7588 17986 7590
rect 18042 7588 18066 7590
rect 18122 7588 18128 7590
rect 17820 7579 18128 7588
rect 24789 7644 25097 7653
rect 24789 7642 24795 7644
rect 24851 7642 24875 7644
rect 24931 7642 24955 7644
rect 25011 7642 25035 7644
rect 25091 7642 25097 7644
rect 24851 7590 24853 7642
rect 25033 7590 25035 7642
rect 24789 7588 24795 7590
rect 24851 7588 24875 7590
rect 24931 7588 24955 7590
rect 25011 7588 25035 7590
rect 25091 7588 25097 7590
rect 24789 7579 25097 7588
rect 7366 7100 7674 7109
rect 7366 7098 7372 7100
rect 7428 7098 7452 7100
rect 7508 7098 7532 7100
rect 7588 7098 7612 7100
rect 7668 7098 7674 7100
rect 7428 7046 7430 7098
rect 7610 7046 7612 7098
rect 7366 7044 7372 7046
rect 7428 7044 7452 7046
rect 7508 7044 7532 7046
rect 7588 7044 7612 7046
rect 7668 7044 7674 7046
rect 7366 7035 7674 7044
rect 14335 7100 14643 7109
rect 14335 7098 14341 7100
rect 14397 7098 14421 7100
rect 14477 7098 14501 7100
rect 14557 7098 14581 7100
rect 14637 7098 14643 7100
rect 14397 7046 14399 7098
rect 14579 7046 14581 7098
rect 14335 7044 14341 7046
rect 14397 7044 14421 7046
rect 14477 7044 14501 7046
rect 14557 7044 14581 7046
rect 14637 7044 14643 7046
rect 14335 7035 14643 7044
rect 21304 7100 21612 7109
rect 21304 7098 21310 7100
rect 21366 7098 21390 7100
rect 21446 7098 21470 7100
rect 21526 7098 21550 7100
rect 21606 7098 21612 7100
rect 21366 7046 21368 7098
rect 21548 7046 21550 7098
rect 21304 7044 21310 7046
rect 21366 7044 21390 7046
rect 21446 7044 21470 7046
rect 21526 7044 21550 7046
rect 21606 7044 21612 7046
rect 21304 7035 21612 7044
rect 28273 7100 28581 7109
rect 28273 7098 28279 7100
rect 28335 7098 28359 7100
rect 28415 7098 28439 7100
rect 28495 7098 28519 7100
rect 28575 7098 28581 7100
rect 28335 7046 28337 7098
rect 28517 7046 28519 7098
rect 28273 7044 28279 7046
rect 28335 7044 28359 7046
rect 28415 7044 28439 7046
rect 28495 7044 28519 7046
rect 28575 7044 28581 7046
rect 28273 7035 28581 7044
rect 3882 6556 4190 6565
rect 3882 6554 3888 6556
rect 3944 6554 3968 6556
rect 4024 6554 4048 6556
rect 4104 6554 4128 6556
rect 4184 6554 4190 6556
rect 3944 6502 3946 6554
rect 4126 6502 4128 6554
rect 3882 6500 3888 6502
rect 3944 6500 3968 6502
rect 4024 6500 4048 6502
rect 4104 6500 4128 6502
rect 4184 6500 4190 6502
rect 3882 6491 4190 6500
rect 10851 6556 11159 6565
rect 10851 6554 10857 6556
rect 10913 6554 10937 6556
rect 10993 6554 11017 6556
rect 11073 6554 11097 6556
rect 11153 6554 11159 6556
rect 10913 6502 10915 6554
rect 11095 6502 11097 6554
rect 10851 6500 10857 6502
rect 10913 6500 10937 6502
rect 10993 6500 11017 6502
rect 11073 6500 11097 6502
rect 11153 6500 11159 6502
rect 10851 6491 11159 6500
rect 17820 6556 18128 6565
rect 17820 6554 17826 6556
rect 17882 6554 17906 6556
rect 17962 6554 17986 6556
rect 18042 6554 18066 6556
rect 18122 6554 18128 6556
rect 17882 6502 17884 6554
rect 18064 6502 18066 6554
rect 17820 6500 17826 6502
rect 17882 6500 17906 6502
rect 17962 6500 17986 6502
rect 18042 6500 18066 6502
rect 18122 6500 18128 6502
rect 17820 6491 18128 6500
rect 24789 6556 25097 6565
rect 24789 6554 24795 6556
rect 24851 6554 24875 6556
rect 24931 6554 24955 6556
rect 25011 6554 25035 6556
rect 25091 6554 25097 6556
rect 24851 6502 24853 6554
rect 25033 6502 25035 6554
rect 24789 6500 24795 6502
rect 24851 6500 24875 6502
rect 24931 6500 24955 6502
rect 25011 6500 25035 6502
rect 25091 6500 25097 6502
rect 24789 6491 25097 6500
rect 7366 6012 7674 6021
rect 7366 6010 7372 6012
rect 7428 6010 7452 6012
rect 7508 6010 7532 6012
rect 7588 6010 7612 6012
rect 7668 6010 7674 6012
rect 7428 5958 7430 6010
rect 7610 5958 7612 6010
rect 7366 5956 7372 5958
rect 7428 5956 7452 5958
rect 7508 5956 7532 5958
rect 7588 5956 7612 5958
rect 7668 5956 7674 5958
rect 7366 5947 7674 5956
rect 14335 6012 14643 6021
rect 14335 6010 14341 6012
rect 14397 6010 14421 6012
rect 14477 6010 14501 6012
rect 14557 6010 14581 6012
rect 14637 6010 14643 6012
rect 14397 5958 14399 6010
rect 14579 5958 14581 6010
rect 14335 5956 14341 5958
rect 14397 5956 14421 5958
rect 14477 5956 14501 5958
rect 14557 5956 14581 5958
rect 14637 5956 14643 5958
rect 14335 5947 14643 5956
rect 21304 6012 21612 6021
rect 21304 6010 21310 6012
rect 21366 6010 21390 6012
rect 21446 6010 21470 6012
rect 21526 6010 21550 6012
rect 21606 6010 21612 6012
rect 21366 5958 21368 6010
rect 21548 5958 21550 6010
rect 21304 5956 21310 5958
rect 21366 5956 21390 5958
rect 21446 5956 21470 5958
rect 21526 5956 21550 5958
rect 21606 5956 21612 5958
rect 21304 5947 21612 5956
rect 28273 6012 28581 6021
rect 28273 6010 28279 6012
rect 28335 6010 28359 6012
rect 28415 6010 28439 6012
rect 28495 6010 28519 6012
rect 28575 6010 28581 6012
rect 28335 5958 28337 6010
rect 28517 5958 28519 6010
rect 28273 5956 28279 5958
rect 28335 5956 28359 5958
rect 28415 5956 28439 5958
rect 28495 5956 28519 5958
rect 28575 5956 28581 5958
rect 28273 5947 28581 5956
rect 3882 5468 4190 5477
rect 3882 5466 3888 5468
rect 3944 5466 3968 5468
rect 4024 5466 4048 5468
rect 4104 5466 4128 5468
rect 4184 5466 4190 5468
rect 3944 5414 3946 5466
rect 4126 5414 4128 5466
rect 3882 5412 3888 5414
rect 3944 5412 3968 5414
rect 4024 5412 4048 5414
rect 4104 5412 4128 5414
rect 4184 5412 4190 5414
rect 3882 5403 4190 5412
rect 10851 5468 11159 5477
rect 10851 5466 10857 5468
rect 10913 5466 10937 5468
rect 10993 5466 11017 5468
rect 11073 5466 11097 5468
rect 11153 5466 11159 5468
rect 10913 5414 10915 5466
rect 11095 5414 11097 5466
rect 10851 5412 10857 5414
rect 10913 5412 10937 5414
rect 10993 5412 11017 5414
rect 11073 5412 11097 5414
rect 11153 5412 11159 5414
rect 10851 5403 11159 5412
rect 17820 5468 18128 5477
rect 17820 5466 17826 5468
rect 17882 5466 17906 5468
rect 17962 5466 17986 5468
rect 18042 5466 18066 5468
rect 18122 5466 18128 5468
rect 17882 5414 17884 5466
rect 18064 5414 18066 5466
rect 17820 5412 17826 5414
rect 17882 5412 17906 5414
rect 17962 5412 17986 5414
rect 18042 5412 18066 5414
rect 18122 5412 18128 5414
rect 17820 5403 18128 5412
rect 24789 5468 25097 5477
rect 24789 5466 24795 5468
rect 24851 5466 24875 5468
rect 24931 5466 24955 5468
rect 25011 5466 25035 5468
rect 25091 5466 25097 5468
rect 24851 5414 24853 5466
rect 25033 5414 25035 5466
rect 24789 5412 24795 5414
rect 24851 5412 24875 5414
rect 24931 5412 24955 5414
rect 25011 5412 25035 5414
rect 25091 5412 25097 5414
rect 24789 5403 25097 5412
rect 7366 4924 7674 4933
rect 7366 4922 7372 4924
rect 7428 4922 7452 4924
rect 7508 4922 7532 4924
rect 7588 4922 7612 4924
rect 7668 4922 7674 4924
rect 7428 4870 7430 4922
rect 7610 4870 7612 4922
rect 7366 4868 7372 4870
rect 7428 4868 7452 4870
rect 7508 4868 7532 4870
rect 7588 4868 7612 4870
rect 7668 4868 7674 4870
rect 7366 4859 7674 4868
rect 14335 4924 14643 4933
rect 14335 4922 14341 4924
rect 14397 4922 14421 4924
rect 14477 4922 14501 4924
rect 14557 4922 14581 4924
rect 14637 4922 14643 4924
rect 14397 4870 14399 4922
rect 14579 4870 14581 4922
rect 14335 4868 14341 4870
rect 14397 4868 14421 4870
rect 14477 4868 14501 4870
rect 14557 4868 14581 4870
rect 14637 4868 14643 4870
rect 14335 4859 14643 4868
rect 21304 4924 21612 4933
rect 21304 4922 21310 4924
rect 21366 4922 21390 4924
rect 21446 4922 21470 4924
rect 21526 4922 21550 4924
rect 21606 4922 21612 4924
rect 21366 4870 21368 4922
rect 21548 4870 21550 4922
rect 21304 4868 21310 4870
rect 21366 4868 21390 4870
rect 21446 4868 21470 4870
rect 21526 4868 21550 4870
rect 21606 4868 21612 4870
rect 21304 4859 21612 4868
rect 28273 4924 28581 4933
rect 28273 4922 28279 4924
rect 28335 4922 28359 4924
rect 28415 4922 28439 4924
rect 28495 4922 28519 4924
rect 28575 4922 28581 4924
rect 28335 4870 28337 4922
rect 28517 4870 28519 4922
rect 28273 4868 28279 4870
rect 28335 4868 28359 4870
rect 28415 4868 28439 4870
rect 28495 4868 28519 4870
rect 28575 4868 28581 4870
rect 28273 4859 28581 4868
rect 3882 4380 4190 4389
rect 3882 4378 3888 4380
rect 3944 4378 3968 4380
rect 4024 4378 4048 4380
rect 4104 4378 4128 4380
rect 4184 4378 4190 4380
rect 3944 4326 3946 4378
rect 4126 4326 4128 4378
rect 3882 4324 3888 4326
rect 3944 4324 3968 4326
rect 4024 4324 4048 4326
rect 4104 4324 4128 4326
rect 4184 4324 4190 4326
rect 3882 4315 4190 4324
rect 10851 4380 11159 4389
rect 10851 4378 10857 4380
rect 10913 4378 10937 4380
rect 10993 4378 11017 4380
rect 11073 4378 11097 4380
rect 11153 4378 11159 4380
rect 10913 4326 10915 4378
rect 11095 4326 11097 4378
rect 10851 4324 10857 4326
rect 10913 4324 10937 4326
rect 10993 4324 11017 4326
rect 11073 4324 11097 4326
rect 11153 4324 11159 4326
rect 10851 4315 11159 4324
rect 17820 4380 18128 4389
rect 17820 4378 17826 4380
rect 17882 4378 17906 4380
rect 17962 4378 17986 4380
rect 18042 4378 18066 4380
rect 18122 4378 18128 4380
rect 17882 4326 17884 4378
rect 18064 4326 18066 4378
rect 17820 4324 17826 4326
rect 17882 4324 17906 4326
rect 17962 4324 17986 4326
rect 18042 4324 18066 4326
rect 18122 4324 18128 4326
rect 17820 4315 18128 4324
rect 24789 4380 25097 4389
rect 24789 4378 24795 4380
rect 24851 4378 24875 4380
rect 24931 4378 24955 4380
rect 25011 4378 25035 4380
rect 25091 4378 25097 4380
rect 24851 4326 24853 4378
rect 25033 4326 25035 4378
rect 24789 4324 24795 4326
rect 24851 4324 24875 4326
rect 24931 4324 24955 4326
rect 25011 4324 25035 4326
rect 25091 4324 25097 4326
rect 24789 4315 25097 4324
rect 7366 3836 7674 3845
rect 7366 3834 7372 3836
rect 7428 3834 7452 3836
rect 7508 3834 7532 3836
rect 7588 3834 7612 3836
rect 7668 3834 7674 3836
rect 7428 3782 7430 3834
rect 7610 3782 7612 3834
rect 7366 3780 7372 3782
rect 7428 3780 7452 3782
rect 7508 3780 7532 3782
rect 7588 3780 7612 3782
rect 7668 3780 7674 3782
rect 7366 3771 7674 3780
rect 14335 3836 14643 3845
rect 14335 3834 14341 3836
rect 14397 3834 14421 3836
rect 14477 3834 14501 3836
rect 14557 3834 14581 3836
rect 14637 3834 14643 3836
rect 14397 3782 14399 3834
rect 14579 3782 14581 3834
rect 14335 3780 14341 3782
rect 14397 3780 14421 3782
rect 14477 3780 14501 3782
rect 14557 3780 14581 3782
rect 14637 3780 14643 3782
rect 14335 3771 14643 3780
rect 21304 3836 21612 3845
rect 21304 3834 21310 3836
rect 21366 3834 21390 3836
rect 21446 3834 21470 3836
rect 21526 3834 21550 3836
rect 21606 3834 21612 3836
rect 21366 3782 21368 3834
rect 21548 3782 21550 3834
rect 21304 3780 21310 3782
rect 21366 3780 21390 3782
rect 21446 3780 21470 3782
rect 21526 3780 21550 3782
rect 21606 3780 21612 3782
rect 21304 3771 21612 3780
rect 28273 3836 28581 3845
rect 28273 3834 28279 3836
rect 28335 3834 28359 3836
rect 28415 3834 28439 3836
rect 28495 3834 28519 3836
rect 28575 3834 28581 3836
rect 28335 3782 28337 3834
rect 28517 3782 28519 3834
rect 28273 3780 28279 3782
rect 28335 3780 28359 3782
rect 28415 3780 28439 3782
rect 28495 3780 28519 3782
rect 28575 3780 28581 3782
rect 28273 3771 28581 3780
rect 3882 3292 4190 3301
rect 3882 3290 3888 3292
rect 3944 3290 3968 3292
rect 4024 3290 4048 3292
rect 4104 3290 4128 3292
rect 4184 3290 4190 3292
rect 3944 3238 3946 3290
rect 4126 3238 4128 3290
rect 3882 3236 3888 3238
rect 3944 3236 3968 3238
rect 4024 3236 4048 3238
rect 4104 3236 4128 3238
rect 4184 3236 4190 3238
rect 3882 3227 4190 3236
rect 10851 3292 11159 3301
rect 10851 3290 10857 3292
rect 10913 3290 10937 3292
rect 10993 3290 11017 3292
rect 11073 3290 11097 3292
rect 11153 3290 11159 3292
rect 10913 3238 10915 3290
rect 11095 3238 11097 3290
rect 10851 3236 10857 3238
rect 10913 3236 10937 3238
rect 10993 3236 11017 3238
rect 11073 3236 11097 3238
rect 11153 3236 11159 3238
rect 10851 3227 11159 3236
rect 17820 3292 18128 3301
rect 17820 3290 17826 3292
rect 17882 3290 17906 3292
rect 17962 3290 17986 3292
rect 18042 3290 18066 3292
rect 18122 3290 18128 3292
rect 17882 3238 17884 3290
rect 18064 3238 18066 3290
rect 17820 3236 17826 3238
rect 17882 3236 17906 3238
rect 17962 3236 17986 3238
rect 18042 3236 18066 3238
rect 18122 3236 18128 3238
rect 17820 3227 18128 3236
rect 24789 3292 25097 3301
rect 24789 3290 24795 3292
rect 24851 3290 24875 3292
rect 24931 3290 24955 3292
rect 25011 3290 25035 3292
rect 25091 3290 25097 3292
rect 24851 3238 24853 3290
rect 25033 3238 25035 3290
rect 24789 3236 24795 3238
rect 24851 3236 24875 3238
rect 24931 3236 24955 3238
rect 25011 3236 25035 3238
rect 25091 3236 25097 3238
rect 24789 3227 25097 3236
rect 7366 2748 7674 2757
rect 7366 2746 7372 2748
rect 7428 2746 7452 2748
rect 7508 2746 7532 2748
rect 7588 2746 7612 2748
rect 7668 2746 7674 2748
rect 7428 2694 7430 2746
rect 7610 2694 7612 2746
rect 7366 2692 7372 2694
rect 7428 2692 7452 2694
rect 7508 2692 7532 2694
rect 7588 2692 7612 2694
rect 7668 2692 7674 2694
rect 7366 2683 7674 2692
rect 14335 2748 14643 2757
rect 14335 2746 14341 2748
rect 14397 2746 14421 2748
rect 14477 2746 14501 2748
rect 14557 2746 14581 2748
rect 14637 2746 14643 2748
rect 14397 2694 14399 2746
rect 14579 2694 14581 2746
rect 14335 2692 14341 2694
rect 14397 2692 14421 2694
rect 14477 2692 14501 2694
rect 14557 2692 14581 2694
rect 14637 2692 14643 2694
rect 14335 2683 14643 2692
rect 21304 2748 21612 2757
rect 21304 2746 21310 2748
rect 21366 2746 21390 2748
rect 21446 2746 21470 2748
rect 21526 2746 21550 2748
rect 21606 2746 21612 2748
rect 21366 2694 21368 2746
rect 21548 2694 21550 2746
rect 21304 2692 21310 2694
rect 21366 2692 21390 2694
rect 21446 2692 21470 2694
rect 21526 2692 21550 2694
rect 21606 2692 21612 2694
rect 21304 2683 21612 2692
rect 28273 2748 28581 2757
rect 28273 2746 28279 2748
rect 28335 2746 28359 2748
rect 28415 2746 28439 2748
rect 28495 2746 28519 2748
rect 28575 2746 28581 2748
rect 28335 2694 28337 2746
rect 28517 2694 28519 2746
rect 28273 2692 28279 2694
rect 28335 2692 28359 2694
rect 28415 2692 28439 2694
rect 28495 2692 28519 2694
rect 28575 2692 28581 2694
rect 28273 2683 28581 2692
rect 3882 2204 4190 2213
rect 3882 2202 3888 2204
rect 3944 2202 3968 2204
rect 4024 2202 4048 2204
rect 4104 2202 4128 2204
rect 4184 2202 4190 2204
rect 3944 2150 3946 2202
rect 4126 2150 4128 2202
rect 3882 2148 3888 2150
rect 3944 2148 3968 2150
rect 4024 2148 4048 2150
rect 4104 2148 4128 2150
rect 4184 2148 4190 2150
rect 3882 2139 4190 2148
rect 10851 2204 11159 2213
rect 10851 2202 10857 2204
rect 10913 2202 10937 2204
rect 10993 2202 11017 2204
rect 11073 2202 11097 2204
rect 11153 2202 11159 2204
rect 10913 2150 10915 2202
rect 11095 2150 11097 2202
rect 10851 2148 10857 2150
rect 10913 2148 10937 2150
rect 10993 2148 11017 2150
rect 11073 2148 11097 2150
rect 11153 2148 11159 2150
rect 10851 2139 11159 2148
rect 17820 2204 18128 2213
rect 17820 2202 17826 2204
rect 17882 2202 17906 2204
rect 17962 2202 17986 2204
rect 18042 2202 18066 2204
rect 18122 2202 18128 2204
rect 17882 2150 17884 2202
rect 18064 2150 18066 2202
rect 17820 2148 17826 2150
rect 17882 2148 17906 2150
rect 17962 2148 17986 2150
rect 18042 2148 18066 2150
rect 18122 2148 18128 2150
rect 17820 2139 18128 2148
rect 24789 2204 25097 2213
rect 24789 2202 24795 2204
rect 24851 2202 24875 2204
rect 24931 2202 24955 2204
rect 25011 2202 25035 2204
rect 25091 2202 25097 2204
rect 24851 2150 24853 2202
rect 25033 2150 25035 2202
rect 24789 2148 24795 2150
rect 24851 2148 24875 2150
rect 24931 2148 24955 2150
rect 25011 2148 25035 2150
rect 25091 2148 25097 2150
rect 24789 2139 25097 2148
rect 7366 1660 7674 1669
rect 7366 1658 7372 1660
rect 7428 1658 7452 1660
rect 7508 1658 7532 1660
rect 7588 1658 7612 1660
rect 7668 1658 7674 1660
rect 7428 1606 7430 1658
rect 7610 1606 7612 1658
rect 7366 1604 7372 1606
rect 7428 1604 7452 1606
rect 7508 1604 7532 1606
rect 7588 1604 7612 1606
rect 7668 1604 7674 1606
rect 7366 1595 7674 1604
rect 14335 1660 14643 1669
rect 14335 1658 14341 1660
rect 14397 1658 14421 1660
rect 14477 1658 14501 1660
rect 14557 1658 14581 1660
rect 14637 1658 14643 1660
rect 14397 1606 14399 1658
rect 14579 1606 14581 1658
rect 14335 1604 14341 1606
rect 14397 1604 14421 1606
rect 14477 1604 14501 1606
rect 14557 1604 14581 1606
rect 14637 1604 14643 1606
rect 14335 1595 14643 1604
rect 21304 1660 21612 1669
rect 21304 1658 21310 1660
rect 21366 1658 21390 1660
rect 21446 1658 21470 1660
rect 21526 1658 21550 1660
rect 21606 1658 21612 1660
rect 21366 1606 21368 1658
rect 21548 1606 21550 1658
rect 21304 1604 21310 1606
rect 21366 1604 21390 1606
rect 21446 1604 21470 1606
rect 21526 1604 21550 1606
rect 21606 1604 21612 1606
rect 21304 1595 21612 1604
rect 28273 1660 28581 1669
rect 28273 1658 28279 1660
rect 28335 1658 28359 1660
rect 28415 1658 28439 1660
rect 28495 1658 28519 1660
rect 28575 1658 28581 1660
rect 28335 1606 28337 1658
rect 28517 1606 28519 1658
rect 28273 1604 28279 1606
rect 28335 1604 28359 1606
rect 28415 1604 28439 1606
rect 28495 1604 28519 1606
rect 28575 1604 28581 1606
rect 28273 1595 28581 1604
rect 3882 1116 4190 1125
rect 3882 1114 3888 1116
rect 3944 1114 3968 1116
rect 4024 1114 4048 1116
rect 4104 1114 4128 1116
rect 4184 1114 4190 1116
rect 3944 1062 3946 1114
rect 4126 1062 4128 1114
rect 3882 1060 3888 1062
rect 3944 1060 3968 1062
rect 4024 1060 4048 1062
rect 4104 1060 4128 1062
rect 4184 1060 4190 1062
rect 3882 1051 4190 1060
rect 10851 1116 11159 1125
rect 10851 1114 10857 1116
rect 10913 1114 10937 1116
rect 10993 1114 11017 1116
rect 11073 1114 11097 1116
rect 11153 1114 11159 1116
rect 10913 1062 10915 1114
rect 11095 1062 11097 1114
rect 10851 1060 10857 1062
rect 10913 1060 10937 1062
rect 10993 1060 11017 1062
rect 11073 1060 11097 1062
rect 11153 1060 11159 1062
rect 10851 1051 11159 1060
rect 17820 1116 18128 1125
rect 17820 1114 17826 1116
rect 17882 1114 17906 1116
rect 17962 1114 17986 1116
rect 18042 1114 18066 1116
rect 18122 1114 18128 1116
rect 17882 1062 17884 1114
rect 18064 1062 18066 1114
rect 17820 1060 17826 1062
rect 17882 1060 17906 1062
rect 17962 1060 17986 1062
rect 18042 1060 18066 1062
rect 18122 1060 18128 1062
rect 17820 1051 18128 1060
rect 24789 1116 25097 1125
rect 24789 1114 24795 1116
rect 24851 1114 24875 1116
rect 24931 1114 24955 1116
rect 25011 1114 25035 1116
rect 25091 1114 25097 1116
rect 24851 1062 24853 1114
rect 25033 1062 25035 1114
rect 24789 1060 24795 1062
rect 24851 1060 24875 1062
rect 24931 1060 24955 1062
rect 25011 1060 25035 1062
rect 25091 1060 25097 1062
rect 24789 1051 25097 1060
rect 7366 572 7674 581
rect 7366 570 7372 572
rect 7428 570 7452 572
rect 7508 570 7532 572
rect 7588 570 7612 572
rect 7668 570 7674 572
rect 7428 518 7430 570
rect 7610 518 7612 570
rect 7366 516 7372 518
rect 7428 516 7452 518
rect 7508 516 7532 518
rect 7588 516 7612 518
rect 7668 516 7674 518
rect 7366 507 7674 516
rect 14335 572 14643 581
rect 14335 570 14341 572
rect 14397 570 14421 572
rect 14477 570 14501 572
rect 14557 570 14581 572
rect 14637 570 14643 572
rect 14397 518 14399 570
rect 14579 518 14581 570
rect 14335 516 14341 518
rect 14397 516 14421 518
rect 14477 516 14501 518
rect 14557 516 14581 518
rect 14637 516 14643 518
rect 14335 507 14643 516
rect 21304 572 21612 581
rect 21304 570 21310 572
rect 21366 570 21390 572
rect 21446 570 21470 572
rect 21526 570 21550 572
rect 21606 570 21612 572
rect 21366 518 21368 570
rect 21548 518 21550 570
rect 21304 516 21310 518
rect 21366 516 21390 518
rect 21446 516 21470 518
rect 21526 516 21550 518
rect 21606 516 21612 518
rect 21304 507 21612 516
rect 28273 572 28581 581
rect 28273 570 28279 572
rect 28335 570 28359 572
rect 28415 570 28439 572
rect 28495 570 28519 572
rect 28575 570 28581 572
rect 28335 518 28337 570
rect 28517 518 28519 570
rect 28273 516 28279 518
rect 28335 516 28359 518
rect 28415 516 28439 518
rect 28495 516 28519 518
rect 28575 516 28581 518
rect 28273 507 28581 516
<< via2 >>
rect 3888 28314 3944 28316
rect 3968 28314 4024 28316
rect 4048 28314 4104 28316
rect 4128 28314 4184 28316
rect 3888 28262 3934 28314
rect 3934 28262 3944 28314
rect 3968 28262 3998 28314
rect 3998 28262 4010 28314
rect 4010 28262 4024 28314
rect 4048 28262 4062 28314
rect 4062 28262 4074 28314
rect 4074 28262 4104 28314
rect 4128 28262 4138 28314
rect 4138 28262 4184 28314
rect 3888 28260 3944 28262
rect 3968 28260 4024 28262
rect 4048 28260 4104 28262
rect 4128 28260 4184 28262
rect 3888 27226 3944 27228
rect 3968 27226 4024 27228
rect 4048 27226 4104 27228
rect 4128 27226 4184 27228
rect 3888 27174 3934 27226
rect 3934 27174 3944 27226
rect 3968 27174 3998 27226
rect 3998 27174 4010 27226
rect 4010 27174 4024 27226
rect 4048 27174 4062 27226
rect 4062 27174 4074 27226
rect 4074 27174 4104 27226
rect 4128 27174 4138 27226
rect 4138 27174 4184 27226
rect 3888 27172 3944 27174
rect 3968 27172 4024 27174
rect 4048 27172 4104 27174
rect 4128 27172 4184 27174
rect 3888 26138 3944 26140
rect 3968 26138 4024 26140
rect 4048 26138 4104 26140
rect 4128 26138 4184 26140
rect 3888 26086 3934 26138
rect 3934 26086 3944 26138
rect 3968 26086 3998 26138
rect 3998 26086 4010 26138
rect 4010 26086 4024 26138
rect 4048 26086 4062 26138
rect 4062 26086 4074 26138
rect 4074 26086 4104 26138
rect 4128 26086 4138 26138
rect 4138 26086 4184 26138
rect 3888 26084 3944 26086
rect 3968 26084 4024 26086
rect 4048 26084 4104 26086
rect 4128 26084 4184 26086
rect 3888 25050 3944 25052
rect 3968 25050 4024 25052
rect 4048 25050 4104 25052
rect 4128 25050 4184 25052
rect 3888 24998 3934 25050
rect 3934 24998 3944 25050
rect 3968 24998 3998 25050
rect 3998 24998 4010 25050
rect 4010 24998 4024 25050
rect 4048 24998 4062 25050
rect 4062 24998 4074 25050
rect 4074 24998 4104 25050
rect 4128 24998 4138 25050
rect 4138 24998 4184 25050
rect 3888 24996 3944 24998
rect 3968 24996 4024 24998
rect 4048 24996 4104 24998
rect 4128 24996 4184 24998
rect 2226 23024 2282 23080
rect 3888 23962 3944 23964
rect 3968 23962 4024 23964
rect 4048 23962 4104 23964
rect 4128 23962 4184 23964
rect 3888 23910 3934 23962
rect 3934 23910 3944 23962
rect 3968 23910 3998 23962
rect 3998 23910 4010 23962
rect 4010 23910 4024 23962
rect 4048 23910 4062 23962
rect 4062 23910 4074 23962
rect 4074 23910 4104 23962
rect 4128 23910 4138 23962
rect 4138 23910 4184 23962
rect 3888 23908 3944 23910
rect 3968 23908 4024 23910
rect 4048 23908 4104 23910
rect 4128 23908 4184 23910
rect 3888 22874 3944 22876
rect 3968 22874 4024 22876
rect 4048 22874 4104 22876
rect 4128 22874 4184 22876
rect 3888 22822 3934 22874
rect 3934 22822 3944 22874
rect 3968 22822 3998 22874
rect 3998 22822 4010 22874
rect 4010 22822 4024 22874
rect 4048 22822 4062 22874
rect 4062 22822 4074 22874
rect 4074 22822 4104 22874
rect 4128 22822 4138 22874
rect 4138 22822 4184 22874
rect 3888 22820 3944 22822
rect 3968 22820 4024 22822
rect 4048 22820 4104 22822
rect 4128 22820 4184 22822
rect 4342 22500 4398 22536
rect 4342 22480 4344 22500
rect 4344 22480 4396 22500
rect 4396 22480 4398 22500
rect 3888 21786 3944 21788
rect 3968 21786 4024 21788
rect 4048 21786 4104 21788
rect 4128 21786 4184 21788
rect 3888 21734 3934 21786
rect 3934 21734 3944 21786
rect 3968 21734 3998 21786
rect 3998 21734 4010 21786
rect 4010 21734 4024 21786
rect 4048 21734 4062 21786
rect 4062 21734 4074 21786
rect 4074 21734 4104 21786
rect 4128 21734 4138 21786
rect 4138 21734 4184 21786
rect 3888 21732 3944 21734
rect 3968 21732 4024 21734
rect 4048 21732 4104 21734
rect 4128 21732 4184 21734
rect 3888 20698 3944 20700
rect 3968 20698 4024 20700
rect 4048 20698 4104 20700
rect 4128 20698 4184 20700
rect 3888 20646 3934 20698
rect 3934 20646 3944 20698
rect 3968 20646 3998 20698
rect 3998 20646 4010 20698
rect 4010 20646 4024 20698
rect 4048 20646 4062 20698
rect 4062 20646 4074 20698
rect 4074 20646 4104 20698
rect 4128 20646 4138 20698
rect 4138 20646 4184 20698
rect 3888 20644 3944 20646
rect 3968 20644 4024 20646
rect 4048 20644 4104 20646
rect 4128 20644 4184 20646
rect 3606 19372 3662 19408
rect 3606 19352 3608 19372
rect 3608 19352 3660 19372
rect 3660 19352 3662 19372
rect 3888 19610 3944 19612
rect 3968 19610 4024 19612
rect 4048 19610 4104 19612
rect 4128 19610 4184 19612
rect 3888 19558 3934 19610
rect 3934 19558 3944 19610
rect 3968 19558 3998 19610
rect 3998 19558 4010 19610
rect 4010 19558 4024 19610
rect 4048 19558 4062 19610
rect 4062 19558 4074 19610
rect 4074 19558 4104 19610
rect 4128 19558 4138 19610
rect 4138 19558 4184 19610
rect 3888 19556 3944 19558
rect 3968 19556 4024 19558
rect 4048 19556 4104 19558
rect 4128 19556 4184 19558
rect 3888 18522 3944 18524
rect 3968 18522 4024 18524
rect 4048 18522 4104 18524
rect 4128 18522 4184 18524
rect 3888 18470 3934 18522
rect 3934 18470 3944 18522
rect 3968 18470 3998 18522
rect 3998 18470 4010 18522
rect 4010 18470 4024 18522
rect 4048 18470 4062 18522
rect 4062 18470 4074 18522
rect 4074 18470 4104 18522
rect 4128 18470 4138 18522
rect 4138 18470 4184 18522
rect 3888 18468 3944 18470
rect 3968 18468 4024 18470
rect 4048 18468 4104 18470
rect 4128 18468 4184 18470
rect 3888 17434 3944 17436
rect 3968 17434 4024 17436
rect 4048 17434 4104 17436
rect 4128 17434 4184 17436
rect 3888 17382 3934 17434
rect 3934 17382 3944 17434
rect 3968 17382 3998 17434
rect 3998 17382 4010 17434
rect 4010 17382 4024 17434
rect 4048 17382 4062 17434
rect 4062 17382 4074 17434
rect 4074 17382 4104 17434
rect 4128 17382 4138 17434
rect 4138 17382 4184 17434
rect 3888 17380 3944 17382
rect 3968 17380 4024 17382
rect 4048 17380 4104 17382
rect 4128 17380 4184 17382
rect 3888 16346 3944 16348
rect 3968 16346 4024 16348
rect 4048 16346 4104 16348
rect 4128 16346 4184 16348
rect 3888 16294 3934 16346
rect 3934 16294 3944 16346
rect 3968 16294 3998 16346
rect 3998 16294 4010 16346
rect 4010 16294 4024 16346
rect 4048 16294 4062 16346
rect 4062 16294 4074 16346
rect 4074 16294 4104 16346
rect 4128 16294 4138 16346
rect 4138 16294 4184 16346
rect 3888 16292 3944 16294
rect 3968 16292 4024 16294
rect 4048 16292 4104 16294
rect 4128 16292 4184 16294
rect 3888 15258 3944 15260
rect 3968 15258 4024 15260
rect 4048 15258 4104 15260
rect 4128 15258 4184 15260
rect 3888 15206 3934 15258
rect 3934 15206 3944 15258
rect 3968 15206 3998 15258
rect 3998 15206 4010 15258
rect 4010 15206 4024 15258
rect 4048 15206 4062 15258
rect 4062 15206 4074 15258
rect 4074 15206 4104 15258
rect 4128 15206 4138 15258
rect 4138 15206 4184 15258
rect 3888 15204 3944 15206
rect 3968 15204 4024 15206
rect 4048 15204 4104 15206
rect 4128 15204 4184 15206
rect 3888 14170 3944 14172
rect 3968 14170 4024 14172
rect 4048 14170 4104 14172
rect 4128 14170 4184 14172
rect 3888 14118 3934 14170
rect 3934 14118 3944 14170
rect 3968 14118 3998 14170
rect 3998 14118 4010 14170
rect 4010 14118 4024 14170
rect 4048 14118 4062 14170
rect 4062 14118 4074 14170
rect 4074 14118 4104 14170
rect 4128 14118 4138 14170
rect 4138 14118 4184 14170
rect 3888 14116 3944 14118
rect 3968 14116 4024 14118
rect 4048 14116 4104 14118
rect 4128 14116 4184 14118
rect 3888 13082 3944 13084
rect 3968 13082 4024 13084
rect 4048 13082 4104 13084
rect 4128 13082 4184 13084
rect 3888 13030 3934 13082
rect 3934 13030 3944 13082
rect 3968 13030 3998 13082
rect 3998 13030 4010 13082
rect 4010 13030 4024 13082
rect 4048 13030 4062 13082
rect 4062 13030 4074 13082
rect 4074 13030 4104 13082
rect 4128 13030 4138 13082
rect 4138 13030 4184 13082
rect 3888 13028 3944 13030
rect 3968 13028 4024 13030
rect 4048 13028 4104 13030
rect 4128 13028 4184 13030
rect 5354 22516 5356 22536
rect 5356 22516 5408 22536
rect 5408 22516 5410 22536
rect 5354 22480 5410 22516
rect 5722 20440 5778 20496
rect 6182 19372 6238 19408
rect 6182 19352 6184 19372
rect 6184 19352 6236 19372
rect 6236 19352 6238 19372
rect 7372 27770 7428 27772
rect 7452 27770 7508 27772
rect 7532 27770 7588 27772
rect 7612 27770 7668 27772
rect 7372 27718 7418 27770
rect 7418 27718 7428 27770
rect 7452 27718 7482 27770
rect 7482 27718 7494 27770
rect 7494 27718 7508 27770
rect 7532 27718 7546 27770
rect 7546 27718 7558 27770
rect 7558 27718 7588 27770
rect 7612 27718 7622 27770
rect 7622 27718 7668 27770
rect 7372 27716 7428 27718
rect 7452 27716 7508 27718
rect 7532 27716 7588 27718
rect 7612 27716 7668 27718
rect 7372 26682 7428 26684
rect 7452 26682 7508 26684
rect 7532 26682 7588 26684
rect 7612 26682 7668 26684
rect 7372 26630 7418 26682
rect 7418 26630 7428 26682
rect 7452 26630 7482 26682
rect 7482 26630 7494 26682
rect 7494 26630 7508 26682
rect 7532 26630 7546 26682
rect 7546 26630 7558 26682
rect 7558 26630 7588 26682
rect 7612 26630 7622 26682
rect 7622 26630 7668 26682
rect 7372 26628 7428 26630
rect 7452 26628 7508 26630
rect 7532 26628 7588 26630
rect 7612 26628 7668 26630
rect 7372 25594 7428 25596
rect 7452 25594 7508 25596
rect 7532 25594 7588 25596
rect 7612 25594 7668 25596
rect 7372 25542 7418 25594
rect 7418 25542 7428 25594
rect 7452 25542 7482 25594
rect 7482 25542 7494 25594
rect 7494 25542 7508 25594
rect 7532 25542 7546 25594
rect 7546 25542 7558 25594
rect 7558 25542 7588 25594
rect 7612 25542 7622 25594
rect 7622 25542 7668 25594
rect 7372 25540 7428 25542
rect 7452 25540 7508 25542
rect 7532 25540 7588 25542
rect 7612 25540 7668 25542
rect 7372 24506 7428 24508
rect 7452 24506 7508 24508
rect 7532 24506 7588 24508
rect 7612 24506 7668 24508
rect 7372 24454 7418 24506
rect 7418 24454 7428 24506
rect 7452 24454 7482 24506
rect 7482 24454 7494 24506
rect 7494 24454 7508 24506
rect 7532 24454 7546 24506
rect 7546 24454 7558 24506
rect 7558 24454 7588 24506
rect 7612 24454 7622 24506
rect 7622 24454 7668 24506
rect 7372 24452 7428 24454
rect 7452 24452 7508 24454
rect 7532 24452 7588 24454
rect 7612 24452 7668 24454
rect 7372 23418 7428 23420
rect 7452 23418 7508 23420
rect 7532 23418 7588 23420
rect 7612 23418 7668 23420
rect 7372 23366 7418 23418
rect 7418 23366 7428 23418
rect 7452 23366 7482 23418
rect 7482 23366 7494 23418
rect 7494 23366 7508 23418
rect 7532 23366 7546 23418
rect 7546 23366 7558 23418
rect 7558 23366 7588 23418
rect 7612 23366 7622 23418
rect 7622 23366 7668 23418
rect 7372 23364 7428 23366
rect 7452 23364 7508 23366
rect 7532 23364 7588 23366
rect 7612 23364 7668 23366
rect 7372 22330 7428 22332
rect 7452 22330 7508 22332
rect 7532 22330 7588 22332
rect 7612 22330 7668 22332
rect 7372 22278 7418 22330
rect 7418 22278 7428 22330
rect 7452 22278 7482 22330
rect 7482 22278 7494 22330
rect 7494 22278 7508 22330
rect 7532 22278 7546 22330
rect 7546 22278 7558 22330
rect 7558 22278 7588 22330
rect 7612 22278 7622 22330
rect 7622 22278 7668 22330
rect 7372 22276 7428 22278
rect 7452 22276 7508 22278
rect 7532 22276 7588 22278
rect 7612 22276 7668 22278
rect 7746 21936 7802 21992
rect 7372 21242 7428 21244
rect 7452 21242 7508 21244
rect 7532 21242 7588 21244
rect 7612 21242 7668 21244
rect 7372 21190 7418 21242
rect 7418 21190 7428 21242
rect 7452 21190 7482 21242
rect 7482 21190 7494 21242
rect 7494 21190 7508 21242
rect 7532 21190 7546 21242
rect 7546 21190 7558 21242
rect 7558 21190 7588 21242
rect 7612 21190 7622 21242
rect 7622 21190 7668 21242
rect 7372 21188 7428 21190
rect 7452 21188 7508 21190
rect 7532 21188 7588 21190
rect 7612 21188 7668 21190
rect 7372 20154 7428 20156
rect 7452 20154 7508 20156
rect 7532 20154 7588 20156
rect 7612 20154 7668 20156
rect 7372 20102 7418 20154
rect 7418 20102 7428 20154
rect 7452 20102 7482 20154
rect 7482 20102 7494 20154
rect 7494 20102 7508 20154
rect 7532 20102 7546 20154
rect 7546 20102 7558 20154
rect 7558 20102 7588 20154
rect 7612 20102 7622 20154
rect 7622 20102 7668 20154
rect 7372 20100 7428 20102
rect 7452 20100 7508 20102
rect 7532 20100 7588 20102
rect 7612 20100 7668 20102
rect 10857 28314 10913 28316
rect 10937 28314 10993 28316
rect 11017 28314 11073 28316
rect 11097 28314 11153 28316
rect 10857 28262 10903 28314
rect 10903 28262 10913 28314
rect 10937 28262 10967 28314
rect 10967 28262 10979 28314
rect 10979 28262 10993 28314
rect 11017 28262 11031 28314
rect 11031 28262 11043 28314
rect 11043 28262 11073 28314
rect 11097 28262 11107 28314
rect 11107 28262 11153 28314
rect 10857 28260 10913 28262
rect 10937 28260 10993 28262
rect 11017 28260 11073 28262
rect 11097 28260 11153 28262
rect 7372 19066 7428 19068
rect 7452 19066 7508 19068
rect 7532 19066 7588 19068
rect 7612 19066 7668 19068
rect 7372 19014 7418 19066
rect 7418 19014 7428 19066
rect 7452 19014 7482 19066
rect 7482 19014 7494 19066
rect 7494 19014 7508 19066
rect 7532 19014 7546 19066
rect 7546 19014 7558 19066
rect 7558 19014 7588 19066
rect 7612 19014 7622 19066
rect 7622 19014 7668 19066
rect 7372 19012 7428 19014
rect 7452 19012 7508 19014
rect 7532 19012 7588 19014
rect 7612 19012 7668 19014
rect 7372 17978 7428 17980
rect 7452 17978 7508 17980
rect 7532 17978 7588 17980
rect 7612 17978 7668 17980
rect 7372 17926 7418 17978
rect 7418 17926 7428 17978
rect 7452 17926 7482 17978
rect 7482 17926 7494 17978
rect 7494 17926 7508 17978
rect 7532 17926 7546 17978
rect 7546 17926 7558 17978
rect 7558 17926 7588 17978
rect 7612 17926 7622 17978
rect 7622 17926 7668 17978
rect 7372 17924 7428 17926
rect 7452 17924 7508 17926
rect 7532 17924 7588 17926
rect 7612 17924 7668 17926
rect 7372 16890 7428 16892
rect 7452 16890 7508 16892
rect 7532 16890 7588 16892
rect 7612 16890 7668 16892
rect 7372 16838 7418 16890
rect 7418 16838 7428 16890
rect 7452 16838 7482 16890
rect 7482 16838 7494 16890
rect 7494 16838 7508 16890
rect 7532 16838 7546 16890
rect 7546 16838 7558 16890
rect 7558 16838 7588 16890
rect 7612 16838 7622 16890
rect 7622 16838 7668 16890
rect 7372 16836 7428 16838
rect 7452 16836 7508 16838
rect 7532 16836 7588 16838
rect 7612 16836 7668 16838
rect 7372 15802 7428 15804
rect 7452 15802 7508 15804
rect 7532 15802 7588 15804
rect 7612 15802 7668 15804
rect 7372 15750 7418 15802
rect 7418 15750 7428 15802
rect 7452 15750 7482 15802
rect 7482 15750 7494 15802
rect 7494 15750 7508 15802
rect 7532 15750 7546 15802
rect 7546 15750 7558 15802
rect 7558 15750 7588 15802
rect 7612 15750 7622 15802
rect 7622 15750 7668 15802
rect 7372 15748 7428 15750
rect 7452 15748 7508 15750
rect 7532 15748 7588 15750
rect 7612 15748 7668 15750
rect 3888 11994 3944 11996
rect 3968 11994 4024 11996
rect 4048 11994 4104 11996
rect 4128 11994 4184 11996
rect 3888 11942 3934 11994
rect 3934 11942 3944 11994
rect 3968 11942 3998 11994
rect 3998 11942 4010 11994
rect 4010 11942 4024 11994
rect 4048 11942 4062 11994
rect 4062 11942 4074 11994
rect 4074 11942 4104 11994
rect 4128 11942 4138 11994
rect 4138 11942 4184 11994
rect 3888 11940 3944 11942
rect 3968 11940 4024 11942
rect 4048 11940 4104 11942
rect 4128 11940 4184 11942
rect 7372 14714 7428 14716
rect 7452 14714 7508 14716
rect 7532 14714 7588 14716
rect 7612 14714 7668 14716
rect 7372 14662 7418 14714
rect 7418 14662 7428 14714
rect 7452 14662 7482 14714
rect 7482 14662 7494 14714
rect 7494 14662 7508 14714
rect 7532 14662 7546 14714
rect 7546 14662 7558 14714
rect 7558 14662 7588 14714
rect 7612 14662 7622 14714
rect 7622 14662 7668 14714
rect 7372 14660 7428 14662
rect 7452 14660 7508 14662
rect 7532 14660 7588 14662
rect 7612 14660 7668 14662
rect 7372 13626 7428 13628
rect 7452 13626 7508 13628
rect 7532 13626 7588 13628
rect 7612 13626 7668 13628
rect 7372 13574 7418 13626
rect 7418 13574 7428 13626
rect 7452 13574 7482 13626
rect 7482 13574 7494 13626
rect 7494 13574 7508 13626
rect 7532 13574 7546 13626
rect 7546 13574 7558 13626
rect 7558 13574 7588 13626
rect 7612 13574 7622 13626
rect 7622 13574 7668 13626
rect 7372 13572 7428 13574
rect 7452 13572 7508 13574
rect 7532 13572 7588 13574
rect 7612 13572 7668 13574
rect 7372 12538 7428 12540
rect 7452 12538 7508 12540
rect 7532 12538 7588 12540
rect 7612 12538 7668 12540
rect 7372 12486 7418 12538
rect 7418 12486 7428 12538
rect 7452 12486 7482 12538
rect 7482 12486 7494 12538
rect 7494 12486 7508 12538
rect 7532 12486 7546 12538
rect 7546 12486 7558 12538
rect 7558 12486 7588 12538
rect 7612 12486 7622 12538
rect 7622 12486 7668 12538
rect 7372 12484 7428 12486
rect 7452 12484 7508 12486
rect 7532 12484 7588 12486
rect 7612 12484 7668 12486
rect 3888 10906 3944 10908
rect 3968 10906 4024 10908
rect 4048 10906 4104 10908
rect 4128 10906 4184 10908
rect 3888 10854 3934 10906
rect 3934 10854 3944 10906
rect 3968 10854 3998 10906
rect 3998 10854 4010 10906
rect 4010 10854 4024 10906
rect 4048 10854 4062 10906
rect 4062 10854 4074 10906
rect 4074 10854 4104 10906
rect 4128 10854 4138 10906
rect 4138 10854 4184 10906
rect 3888 10852 3944 10854
rect 3968 10852 4024 10854
rect 4048 10852 4104 10854
rect 4128 10852 4184 10854
rect 10857 27226 10913 27228
rect 10937 27226 10993 27228
rect 11017 27226 11073 27228
rect 11097 27226 11153 27228
rect 10857 27174 10903 27226
rect 10903 27174 10913 27226
rect 10937 27174 10967 27226
rect 10967 27174 10979 27226
rect 10979 27174 10993 27226
rect 11017 27174 11031 27226
rect 11031 27174 11043 27226
rect 11043 27174 11073 27226
rect 11097 27174 11107 27226
rect 11107 27174 11153 27226
rect 10857 27172 10913 27174
rect 10937 27172 10993 27174
rect 11017 27172 11073 27174
rect 11097 27172 11153 27174
rect 10857 26138 10913 26140
rect 10937 26138 10993 26140
rect 11017 26138 11073 26140
rect 11097 26138 11153 26140
rect 10857 26086 10903 26138
rect 10903 26086 10913 26138
rect 10937 26086 10967 26138
rect 10967 26086 10979 26138
rect 10979 26086 10993 26138
rect 11017 26086 11031 26138
rect 11031 26086 11043 26138
rect 11043 26086 11073 26138
rect 11097 26086 11107 26138
rect 11107 26086 11153 26138
rect 10857 26084 10913 26086
rect 10937 26084 10993 26086
rect 11017 26084 11073 26086
rect 11097 26084 11153 26086
rect 10857 25050 10913 25052
rect 10937 25050 10993 25052
rect 11017 25050 11073 25052
rect 11097 25050 11153 25052
rect 10857 24998 10903 25050
rect 10903 24998 10913 25050
rect 10937 24998 10967 25050
rect 10967 24998 10979 25050
rect 10979 24998 10993 25050
rect 11017 24998 11031 25050
rect 11031 24998 11043 25050
rect 11043 24998 11073 25050
rect 11097 24998 11107 25050
rect 11107 24998 11153 25050
rect 10857 24996 10913 24998
rect 10937 24996 10993 24998
rect 11017 24996 11073 24998
rect 11097 24996 11153 24998
rect 10857 23962 10913 23964
rect 10937 23962 10993 23964
rect 11017 23962 11073 23964
rect 11097 23962 11153 23964
rect 10857 23910 10903 23962
rect 10903 23910 10913 23962
rect 10937 23910 10967 23962
rect 10967 23910 10979 23962
rect 10979 23910 10993 23962
rect 11017 23910 11031 23962
rect 11031 23910 11043 23962
rect 11043 23910 11073 23962
rect 11097 23910 11107 23962
rect 11107 23910 11153 23962
rect 10857 23908 10913 23910
rect 10937 23908 10993 23910
rect 11017 23908 11073 23910
rect 11097 23908 11153 23910
rect 9862 20884 9864 20904
rect 9864 20884 9916 20904
rect 9916 20884 9918 20904
rect 9862 20848 9918 20884
rect 7372 11450 7428 11452
rect 7452 11450 7508 11452
rect 7532 11450 7588 11452
rect 7612 11450 7668 11452
rect 7372 11398 7418 11450
rect 7418 11398 7428 11450
rect 7452 11398 7482 11450
rect 7482 11398 7494 11450
rect 7494 11398 7508 11450
rect 7532 11398 7546 11450
rect 7546 11398 7558 11450
rect 7558 11398 7588 11450
rect 7612 11398 7622 11450
rect 7622 11398 7668 11450
rect 7372 11396 7428 11398
rect 7452 11396 7508 11398
rect 7532 11396 7588 11398
rect 7612 11396 7668 11398
rect 10857 22874 10913 22876
rect 10937 22874 10993 22876
rect 11017 22874 11073 22876
rect 11097 22874 11153 22876
rect 10857 22822 10903 22874
rect 10903 22822 10913 22874
rect 10937 22822 10967 22874
rect 10967 22822 10979 22874
rect 10979 22822 10993 22874
rect 11017 22822 11031 22874
rect 11031 22822 11043 22874
rect 11043 22822 11073 22874
rect 11097 22822 11107 22874
rect 11107 22822 11153 22874
rect 10857 22820 10913 22822
rect 10937 22820 10993 22822
rect 11017 22820 11073 22822
rect 11097 22820 11153 22822
rect 14341 27770 14397 27772
rect 14421 27770 14477 27772
rect 14501 27770 14557 27772
rect 14581 27770 14637 27772
rect 14341 27718 14387 27770
rect 14387 27718 14397 27770
rect 14421 27718 14451 27770
rect 14451 27718 14463 27770
rect 14463 27718 14477 27770
rect 14501 27718 14515 27770
rect 14515 27718 14527 27770
rect 14527 27718 14557 27770
rect 14581 27718 14591 27770
rect 14591 27718 14637 27770
rect 14341 27716 14397 27718
rect 14421 27716 14477 27718
rect 14501 27716 14557 27718
rect 14581 27716 14637 27718
rect 17826 28314 17882 28316
rect 17906 28314 17962 28316
rect 17986 28314 18042 28316
rect 18066 28314 18122 28316
rect 17826 28262 17872 28314
rect 17872 28262 17882 28314
rect 17906 28262 17936 28314
rect 17936 28262 17948 28314
rect 17948 28262 17962 28314
rect 17986 28262 18000 28314
rect 18000 28262 18012 28314
rect 18012 28262 18042 28314
rect 18066 28262 18076 28314
rect 18076 28262 18122 28314
rect 17826 28260 17882 28262
rect 17906 28260 17962 28262
rect 17986 28260 18042 28262
rect 18066 28260 18122 28262
rect 24795 28314 24851 28316
rect 24875 28314 24931 28316
rect 24955 28314 25011 28316
rect 25035 28314 25091 28316
rect 24795 28262 24841 28314
rect 24841 28262 24851 28314
rect 24875 28262 24905 28314
rect 24905 28262 24917 28314
rect 24917 28262 24931 28314
rect 24955 28262 24969 28314
rect 24969 28262 24981 28314
rect 24981 28262 25011 28314
rect 25035 28262 25045 28314
rect 25045 28262 25091 28314
rect 24795 28260 24851 28262
rect 24875 28260 24931 28262
rect 24955 28260 25011 28262
rect 25035 28260 25091 28262
rect 10857 21786 10913 21788
rect 10937 21786 10993 21788
rect 11017 21786 11073 21788
rect 11097 21786 11153 21788
rect 10857 21734 10903 21786
rect 10903 21734 10913 21786
rect 10937 21734 10967 21786
rect 10967 21734 10979 21786
rect 10979 21734 10993 21786
rect 11017 21734 11031 21786
rect 11031 21734 11043 21786
rect 11043 21734 11073 21786
rect 11097 21734 11107 21786
rect 11107 21734 11153 21786
rect 10857 21732 10913 21734
rect 10937 21732 10993 21734
rect 11017 21732 11073 21734
rect 11097 21732 11153 21734
rect 10857 20698 10913 20700
rect 10937 20698 10993 20700
rect 11017 20698 11073 20700
rect 11097 20698 11153 20700
rect 10857 20646 10903 20698
rect 10903 20646 10913 20698
rect 10937 20646 10967 20698
rect 10967 20646 10979 20698
rect 10979 20646 10993 20698
rect 11017 20646 11031 20698
rect 11031 20646 11043 20698
rect 11043 20646 11073 20698
rect 11097 20646 11107 20698
rect 11107 20646 11153 20698
rect 10857 20644 10913 20646
rect 10937 20644 10993 20646
rect 11017 20644 11073 20646
rect 11097 20644 11153 20646
rect 11058 20440 11114 20496
rect 11610 21392 11666 21448
rect 10857 19610 10913 19612
rect 10937 19610 10993 19612
rect 11017 19610 11073 19612
rect 11097 19610 11153 19612
rect 10857 19558 10903 19610
rect 10903 19558 10913 19610
rect 10937 19558 10967 19610
rect 10967 19558 10979 19610
rect 10979 19558 10993 19610
rect 11017 19558 11031 19610
rect 11031 19558 11043 19610
rect 11043 19558 11073 19610
rect 11097 19558 11107 19610
rect 11107 19558 11153 19610
rect 10857 19556 10913 19558
rect 10937 19556 10993 19558
rect 11017 19556 11073 19558
rect 11097 19556 11153 19558
rect 10857 18522 10913 18524
rect 10937 18522 10993 18524
rect 11017 18522 11073 18524
rect 11097 18522 11153 18524
rect 10857 18470 10903 18522
rect 10903 18470 10913 18522
rect 10937 18470 10967 18522
rect 10967 18470 10979 18522
rect 10979 18470 10993 18522
rect 11017 18470 11031 18522
rect 11031 18470 11043 18522
rect 11043 18470 11073 18522
rect 11097 18470 11107 18522
rect 11107 18470 11153 18522
rect 10857 18468 10913 18470
rect 10937 18468 10993 18470
rect 11017 18468 11073 18470
rect 11097 18468 11153 18470
rect 10857 17434 10913 17436
rect 10937 17434 10993 17436
rect 11017 17434 11073 17436
rect 11097 17434 11153 17436
rect 10857 17382 10903 17434
rect 10903 17382 10913 17434
rect 10937 17382 10967 17434
rect 10967 17382 10979 17434
rect 10979 17382 10993 17434
rect 11017 17382 11031 17434
rect 11031 17382 11043 17434
rect 11043 17382 11073 17434
rect 11097 17382 11107 17434
rect 11107 17382 11153 17434
rect 10857 17380 10913 17382
rect 10937 17380 10993 17382
rect 11017 17380 11073 17382
rect 11097 17380 11153 17382
rect 10857 16346 10913 16348
rect 10937 16346 10993 16348
rect 11017 16346 11073 16348
rect 11097 16346 11153 16348
rect 10857 16294 10903 16346
rect 10903 16294 10913 16346
rect 10937 16294 10967 16346
rect 10967 16294 10979 16346
rect 10979 16294 10993 16346
rect 11017 16294 11031 16346
rect 11031 16294 11043 16346
rect 11043 16294 11073 16346
rect 11097 16294 11107 16346
rect 11107 16294 11153 16346
rect 10857 16292 10913 16294
rect 10937 16292 10993 16294
rect 11017 16292 11073 16294
rect 11097 16292 11153 16294
rect 11886 21392 11942 21448
rect 12346 22888 12402 22944
rect 14341 26682 14397 26684
rect 14421 26682 14477 26684
rect 14501 26682 14557 26684
rect 14581 26682 14637 26684
rect 14341 26630 14387 26682
rect 14387 26630 14397 26682
rect 14421 26630 14451 26682
rect 14451 26630 14463 26682
rect 14463 26630 14477 26682
rect 14501 26630 14515 26682
rect 14515 26630 14527 26682
rect 14527 26630 14557 26682
rect 14581 26630 14591 26682
rect 14591 26630 14637 26682
rect 14341 26628 14397 26630
rect 14421 26628 14477 26630
rect 14501 26628 14557 26630
rect 14581 26628 14637 26630
rect 14341 25594 14397 25596
rect 14421 25594 14477 25596
rect 14501 25594 14557 25596
rect 14581 25594 14637 25596
rect 14341 25542 14387 25594
rect 14387 25542 14397 25594
rect 14421 25542 14451 25594
rect 14451 25542 14463 25594
rect 14463 25542 14477 25594
rect 14501 25542 14515 25594
rect 14515 25542 14527 25594
rect 14527 25542 14557 25594
rect 14581 25542 14591 25594
rect 14591 25542 14637 25594
rect 14341 25540 14397 25542
rect 14421 25540 14477 25542
rect 14501 25540 14557 25542
rect 14581 25540 14637 25542
rect 13726 25356 13782 25392
rect 13726 25336 13728 25356
rect 13728 25336 13780 25356
rect 13780 25336 13782 25356
rect 17826 27226 17882 27228
rect 17906 27226 17962 27228
rect 17986 27226 18042 27228
rect 18066 27226 18122 27228
rect 17826 27174 17872 27226
rect 17872 27174 17882 27226
rect 17906 27174 17936 27226
rect 17936 27174 17948 27226
rect 17948 27174 17962 27226
rect 17986 27174 18000 27226
rect 18000 27174 18012 27226
rect 18012 27174 18042 27226
rect 18066 27174 18076 27226
rect 18076 27174 18122 27226
rect 17826 27172 17882 27174
rect 17906 27172 17962 27174
rect 17986 27172 18042 27174
rect 18066 27172 18122 27174
rect 14341 24506 14397 24508
rect 14421 24506 14477 24508
rect 14501 24506 14557 24508
rect 14581 24506 14637 24508
rect 14341 24454 14387 24506
rect 14387 24454 14397 24506
rect 14421 24454 14451 24506
rect 14451 24454 14463 24506
rect 14463 24454 14477 24506
rect 14501 24454 14515 24506
rect 14515 24454 14527 24506
rect 14527 24454 14557 24506
rect 14581 24454 14591 24506
rect 14591 24454 14637 24506
rect 14341 24452 14397 24454
rect 14421 24452 14477 24454
rect 14501 24452 14557 24454
rect 14581 24452 14637 24454
rect 13174 23044 13230 23080
rect 13174 23024 13176 23044
rect 13176 23024 13228 23044
rect 13228 23024 13230 23044
rect 13726 23024 13782 23080
rect 14341 23418 14397 23420
rect 14421 23418 14477 23420
rect 14501 23418 14557 23420
rect 14581 23418 14637 23420
rect 14341 23366 14387 23418
rect 14387 23366 14397 23418
rect 14421 23366 14451 23418
rect 14451 23366 14463 23418
rect 14463 23366 14477 23418
rect 14501 23366 14515 23418
rect 14515 23366 14527 23418
rect 14527 23366 14557 23418
rect 14581 23366 14591 23418
rect 14591 23366 14637 23418
rect 14341 23364 14397 23366
rect 14421 23364 14477 23366
rect 14501 23364 14557 23366
rect 14581 23364 14637 23366
rect 13726 21936 13782 21992
rect 10857 15258 10913 15260
rect 10937 15258 10993 15260
rect 11017 15258 11073 15260
rect 11097 15258 11153 15260
rect 10857 15206 10903 15258
rect 10903 15206 10913 15258
rect 10937 15206 10967 15258
rect 10967 15206 10979 15258
rect 10979 15206 10993 15258
rect 11017 15206 11031 15258
rect 11031 15206 11043 15258
rect 11043 15206 11073 15258
rect 11097 15206 11107 15258
rect 11107 15206 11153 15258
rect 10857 15204 10913 15206
rect 10937 15204 10993 15206
rect 11017 15204 11073 15206
rect 11097 15204 11153 15206
rect 10322 14864 10378 14920
rect 10857 14170 10913 14172
rect 10937 14170 10993 14172
rect 11017 14170 11073 14172
rect 11097 14170 11153 14172
rect 10857 14118 10903 14170
rect 10903 14118 10913 14170
rect 10937 14118 10967 14170
rect 10967 14118 10979 14170
rect 10979 14118 10993 14170
rect 11017 14118 11031 14170
rect 11031 14118 11043 14170
rect 11043 14118 11073 14170
rect 11097 14118 11107 14170
rect 11107 14118 11153 14170
rect 10857 14116 10913 14118
rect 10937 14116 10993 14118
rect 11017 14116 11073 14118
rect 11097 14116 11153 14118
rect 11702 14900 11704 14920
rect 11704 14900 11756 14920
rect 11756 14900 11758 14920
rect 11702 14864 11758 14900
rect 10857 13082 10913 13084
rect 10937 13082 10993 13084
rect 11017 13082 11073 13084
rect 11097 13082 11153 13084
rect 10857 13030 10903 13082
rect 10903 13030 10913 13082
rect 10937 13030 10967 13082
rect 10967 13030 10979 13082
rect 10979 13030 10993 13082
rect 11017 13030 11031 13082
rect 11031 13030 11043 13082
rect 11043 13030 11073 13082
rect 11097 13030 11107 13082
rect 11107 13030 11153 13082
rect 10857 13028 10913 13030
rect 10937 13028 10993 13030
rect 11017 13028 11073 13030
rect 11097 13028 11153 13030
rect 7372 10362 7428 10364
rect 7452 10362 7508 10364
rect 7532 10362 7588 10364
rect 7612 10362 7668 10364
rect 7372 10310 7418 10362
rect 7418 10310 7428 10362
rect 7452 10310 7482 10362
rect 7482 10310 7494 10362
rect 7494 10310 7508 10362
rect 7532 10310 7546 10362
rect 7546 10310 7558 10362
rect 7558 10310 7588 10362
rect 7612 10310 7622 10362
rect 7622 10310 7668 10362
rect 7372 10308 7428 10310
rect 7452 10308 7508 10310
rect 7532 10308 7588 10310
rect 7612 10308 7668 10310
rect 10857 11994 10913 11996
rect 10937 11994 10993 11996
rect 11017 11994 11073 11996
rect 11097 11994 11153 11996
rect 10857 11942 10903 11994
rect 10903 11942 10913 11994
rect 10937 11942 10967 11994
rect 10967 11942 10979 11994
rect 10979 11942 10993 11994
rect 11017 11942 11031 11994
rect 11031 11942 11043 11994
rect 11043 11942 11073 11994
rect 11097 11942 11107 11994
rect 11107 11942 11153 11994
rect 10857 11940 10913 11942
rect 10937 11940 10993 11942
rect 11017 11940 11073 11942
rect 11097 11940 11153 11942
rect 10857 10906 10913 10908
rect 10937 10906 10993 10908
rect 11017 10906 11073 10908
rect 11097 10906 11153 10908
rect 10857 10854 10903 10906
rect 10903 10854 10913 10906
rect 10937 10854 10967 10906
rect 10967 10854 10979 10906
rect 10979 10854 10993 10906
rect 11017 10854 11031 10906
rect 11031 10854 11043 10906
rect 11043 10854 11073 10906
rect 11097 10854 11107 10906
rect 11107 10854 11153 10906
rect 10857 10852 10913 10854
rect 10937 10852 10993 10854
rect 11017 10852 11073 10854
rect 11097 10852 11153 10854
rect 12990 17040 13046 17096
rect 14341 22330 14397 22332
rect 14421 22330 14477 22332
rect 14501 22330 14557 22332
rect 14581 22330 14637 22332
rect 14341 22278 14387 22330
rect 14387 22278 14397 22330
rect 14421 22278 14451 22330
rect 14451 22278 14463 22330
rect 14463 22278 14477 22330
rect 14501 22278 14515 22330
rect 14515 22278 14527 22330
rect 14527 22278 14557 22330
rect 14581 22278 14591 22330
rect 14591 22278 14637 22330
rect 14341 22276 14397 22278
rect 14421 22276 14477 22278
rect 14501 22276 14557 22278
rect 14581 22276 14637 22278
rect 14341 21242 14397 21244
rect 14421 21242 14477 21244
rect 14501 21242 14557 21244
rect 14581 21242 14637 21244
rect 14341 21190 14387 21242
rect 14387 21190 14397 21242
rect 14421 21190 14451 21242
rect 14451 21190 14463 21242
rect 14463 21190 14477 21242
rect 14501 21190 14515 21242
rect 14515 21190 14527 21242
rect 14527 21190 14557 21242
rect 14581 21190 14591 21242
rect 14591 21190 14637 21242
rect 14341 21188 14397 21190
rect 14421 21188 14477 21190
rect 14501 21188 14557 21190
rect 14581 21188 14637 21190
rect 14094 20748 14096 20768
rect 14096 20748 14148 20768
rect 14148 20748 14150 20768
rect 14094 20712 14150 20748
rect 14341 20154 14397 20156
rect 14421 20154 14477 20156
rect 14501 20154 14557 20156
rect 14581 20154 14637 20156
rect 14341 20102 14387 20154
rect 14387 20102 14397 20154
rect 14421 20102 14451 20154
rect 14451 20102 14463 20154
rect 14463 20102 14477 20154
rect 14501 20102 14515 20154
rect 14515 20102 14527 20154
rect 14527 20102 14557 20154
rect 14581 20102 14591 20154
rect 14591 20102 14637 20154
rect 14341 20100 14397 20102
rect 14421 20100 14477 20102
rect 14501 20100 14557 20102
rect 14581 20100 14637 20102
rect 13358 17584 13414 17640
rect 14341 19066 14397 19068
rect 14421 19066 14477 19068
rect 14501 19066 14557 19068
rect 14581 19066 14637 19068
rect 14341 19014 14387 19066
rect 14387 19014 14397 19066
rect 14421 19014 14451 19066
rect 14451 19014 14463 19066
rect 14463 19014 14477 19066
rect 14501 19014 14515 19066
rect 14515 19014 14527 19066
rect 14527 19014 14557 19066
rect 14581 19014 14591 19066
rect 14591 19014 14637 19066
rect 14341 19012 14397 19014
rect 14421 19012 14477 19014
rect 14501 19012 14557 19014
rect 14581 19012 14637 19014
rect 13450 16360 13506 16416
rect 14341 17978 14397 17980
rect 14421 17978 14477 17980
rect 14501 17978 14557 17980
rect 14581 17978 14637 17980
rect 14341 17926 14387 17978
rect 14387 17926 14397 17978
rect 14421 17926 14451 17978
rect 14451 17926 14463 17978
rect 14463 17926 14477 17978
rect 14501 17926 14515 17978
rect 14515 17926 14527 17978
rect 14527 17926 14557 17978
rect 14581 17926 14591 17978
rect 14591 17926 14637 17978
rect 14341 17924 14397 17926
rect 14421 17924 14477 17926
rect 14501 17924 14557 17926
rect 14581 17924 14637 17926
rect 15014 23196 15016 23216
rect 15016 23196 15068 23216
rect 15068 23196 15070 23216
rect 15014 23160 15070 23196
rect 21310 27770 21366 27772
rect 21390 27770 21446 27772
rect 21470 27770 21526 27772
rect 21550 27770 21606 27772
rect 21310 27718 21356 27770
rect 21356 27718 21366 27770
rect 21390 27718 21420 27770
rect 21420 27718 21432 27770
rect 21432 27718 21446 27770
rect 21470 27718 21484 27770
rect 21484 27718 21496 27770
rect 21496 27718 21526 27770
rect 21550 27718 21560 27770
rect 21560 27718 21606 27770
rect 21310 27716 21366 27718
rect 21390 27716 21446 27718
rect 21470 27716 21526 27718
rect 21550 27716 21606 27718
rect 15842 22924 15844 22944
rect 15844 22924 15896 22944
rect 15896 22924 15898 22944
rect 15842 22888 15898 22924
rect 14646 17620 14648 17640
rect 14648 17620 14700 17640
rect 14700 17620 14702 17640
rect 14646 17584 14702 17620
rect 17826 26138 17882 26140
rect 17906 26138 17962 26140
rect 17986 26138 18042 26140
rect 18066 26138 18122 26140
rect 17826 26086 17872 26138
rect 17872 26086 17882 26138
rect 17906 26086 17936 26138
rect 17936 26086 17948 26138
rect 17948 26086 17962 26138
rect 17986 26086 18000 26138
rect 18000 26086 18012 26138
rect 18012 26086 18042 26138
rect 18066 26086 18076 26138
rect 18076 26086 18122 26138
rect 17826 26084 17882 26086
rect 17906 26084 17962 26086
rect 17986 26084 18042 26086
rect 18066 26084 18122 26086
rect 14341 16890 14397 16892
rect 14421 16890 14477 16892
rect 14501 16890 14557 16892
rect 14581 16890 14637 16892
rect 14341 16838 14387 16890
rect 14387 16838 14397 16890
rect 14421 16838 14451 16890
rect 14451 16838 14463 16890
rect 14463 16838 14477 16890
rect 14501 16838 14515 16890
rect 14515 16838 14527 16890
rect 14527 16838 14557 16890
rect 14581 16838 14591 16890
rect 14591 16838 14637 16890
rect 14341 16836 14397 16838
rect 14421 16836 14477 16838
rect 14501 16836 14557 16838
rect 14581 16836 14637 16838
rect 14341 15802 14397 15804
rect 14421 15802 14477 15804
rect 14501 15802 14557 15804
rect 14581 15802 14637 15804
rect 14341 15750 14387 15802
rect 14387 15750 14397 15802
rect 14421 15750 14451 15802
rect 14451 15750 14463 15802
rect 14463 15750 14477 15802
rect 14501 15750 14515 15802
rect 14515 15750 14527 15802
rect 14527 15750 14557 15802
rect 14581 15750 14591 15802
rect 14591 15750 14637 15802
rect 14341 15748 14397 15750
rect 14421 15748 14477 15750
rect 14501 15748 14557 15750
rect 14581 15748 14637 15750
rect 13450 12824 13506 12880
rect 13910 12688 13966 12744
rect 14341 14714 14397 14716
rect 14421 14714 14477 14716
rect 14501 14714 14557 14716
rect 14581 14714 14637 14716
rect 14341 14662 14387 14714
rect 14387 14662 14397 14714
rect 14421 14662 14451 14714
rect 14451 14662 14463 14714
rect 14463 14662 14477 14714
rect 14501 14662 14515 14714
rect 14515 14662 14527 14714
rect 14527 14662 14557 14714
rect 14581 14662 14591 14714
rect 14591 14662 14637 14714
rect 14341 14660 14397 14662
rect 14421 14660 14477 14662
rect 14501 14660 14557 14662
rect 14581 14660 14637 14662
rect 14341 13626 14397 13628
rect 14421 13626 14477 13628
rect 14501 13626 14557 13628
rect 14581 13626 14637 13628
rect 14341 13574 14387 13626
rect 14387 13574 14397 13626
rect 14421 13574 14451 13626
rect 14451 13574 14463 13626
rect 14463 13574 14477 13626
rect 14501 13574 14515 13626
rect 14515 13574 14527 13626
rect 14527 13574 14557 13626
rect 14581 13574 14591 13626
rect 14591 13574 14637 13626
rect 14341 13572 14397 13574
rect 14421 13572 14477 13574
rect 14501 13572 14557 13574
rect 14581 13572 14637 13574
rect 14341 12538 14397 12540
rect 14421 12538 14477 12540
rect 14501 12538 14557 12540
rect 14581 12538 14637 12540
rect 14341 12486 14387 12538
rect 14387 12486 14397 12538
rect 14421 12486 14451 12538
rect 14451 12486 14463 12538
rect 14463 12486 14477 12538
rect 14501 12486 14515 12538
rect 14515 12486 14527 12538
rect 14527 12486 14557 12538
rect 14581 12486 14591 12538
rect 14591 12486 14637 12538
rect 14341 12484 14397 12486
rect 14421 12484 14477 12486
rect 14501 12484 14557 12486
rect 14581 12484 14637 12486
rect 16762 21392 16818 21448
rect 17826 25050 17882 25052
rect 17906 25050 17962 25052
rect 17986 25050 18042 25052
rect 18066 25050 18122 25052
rect 17826 24998 17872 25050
rect 17872 24998 17882 25050
rect 17906 24998 17936 25050
rect 17936 24998 17948 25050
rect 17948 24998 17962 25050
rect 17986 24998 18000 25050
rect 18000 24998 18012 25050
rect 18012 24998 18042 25050
rect 18066 24998 18076 25050
rect 18076 24998 18122 25050
rect 17826 24996 17882 24998
rect 17906 24996 17962 24998
rect 17986 24996 18042 24998
rect 18066 24996 18122 24998
rect 17826 23962 17882 23964
rect 17906 23962 17962 23964
rect 17986 23962 18042 23964
rect 18066 23962 18122 23964
rect 17826 23910 17872 23962
rect 17872 23910 17882 23962
rect 17906 23910 17936 23962
rect 17936 23910 17948 23962
rect 17948 23910 17962 23962
rect 17986 23910 18000 23962
rect 18000 23910 18012 23962
rect 18012 23910 18042 23962
rect 18066 23910 18076 23962
rect 18076 23910 18122 23962
rect 17826 23908 17882 23910
rect 17906 23908 17962 23910
rect 17986 23908 18042 23910
rect 18066 23908 18122 23910
rect 17314 23024 17370 23080
rect 17826 22874 17882 22876
rect 17906 22874 17962 22876
rect 17986 22874 18042 22876
rect 18066 22874 18122 22876
rect 17826 22822 17872 22874
rect 17872 22822 17882 22874
rect 17906 22822 17936 22874
rect 17936 22822 17948 22874
rect 17948 22822 17962 22874
rect 17986 22822 18000 22874
rect 18000 22822 18012 22874
rect 18012 22822 18042 22874
rect 18066 22822 18076 22874
rect 18076 22822 18122 22874
rect 17826 22820 17882 22822
rect 17906 22820 17962 22822
rect 17986 22820 18042 22822
rect 18066 22820 18122 22822
rect 18602 25372 18604 25392
rect 18604 25372 18656 25392
rect 18656 25372 18658 25392
rect 18602 25336 18658 25372
rect 17826 21786 17882 21788
rect 17906 21786 17962 21788
rect 17986 21786 18042 21788
rect 18066 21786 18122 21788
rect 17826 21734 17872 21786
rect 17872 21734 17882 21786
rect 17906 21734 17936 21786
rect 17936 21734 17948 21786
rect 17948 21734 17962 21786
rect 17986 21734 18000 21786
rect 18000 21734 18012 21786
rect 18012 21734 18042 21786
rect 18066 21734 18076 21786
rect 18076 21734 18122 21786
rect 17826 21732 17882 21734
rect 17906 21732 17962 21734
rect 17986 21732 18042 21734
rect 18066 21732 18122 21734
rect 17826 20698 17882 20700
rect 17906 20698 17962 20700
rect 17986 20698 18042 20700
rect 18066 20698 18122 20700
rect 17826 20646 17872 20698
rect 17872 20646 17882 20698
rect 17906 20646 17936 20698
rect 17936 20646 17948 20698
rect 17948 20646 17962 20698
rect 17986 20646 18000 20698
rect 18000 20646 18012 20698
rect 18012 20646 18042 20698
rect 18066 20646 18076 20698
rect 18076 20646 18122 20698
rect 17826 20644 17882 20646
rect 17906 20644 17962 20646
rect 17986 20644 18042 20646
rect 18066 20644 18122 20646
rect 17826 19610 17882 19612
rect 17906 19610 17962 19612
rect 17986 19610 18042 19612
rect 18066 19610 18122 19612
rect 17826 19558 17872 19610
rect 17872 19558 17882 19610
rect 17906 19558 17936 19610
rect 17936 19558 17948 19610
rect 17948 19558 17962 19610
rect 17986 19558 18000 19610
rect 18000 19558 18012 19610
rect 18012 19558 18042 19610
rect 18066 19558 18076 19610
rect 18076 19558 18122 19610
rect 17826 19556 17882 19558
rect 17906 19556 17962 19558
rect 17986 19556 18042 19558
rect 18066 19556 18122 19558
rect 16854 17040 16910 17096
rect 15750 16124 15752 16144
rect 15752 16124 15804 16144
rect 15804 16124 15806 16144
rect 15750 16088 15806 16124
rect 15934 15952 15990 16008
rect 17826 18522 17882 18524
rect 17906 18522 17962 18524
rect 17986 18522 18042 18524
rect 18066 18522 18122 18524
rect 17826 18470 17872 18522
rect 17872 18470 17882 18522
rect 17906 18470 17936 18522
rect 17936 18470 17948 18522
rect 17948 18470 17962 18522
rect 17986 18470 18000 18522
rect 18000 18470 18012 18522
rect 18012 18470 18042 18522
rect 18066 18470 18076 18522
rect 18076 18470 18122 18522
rect 17826 18468 17882 18470
rect 17906 18468 17962 18470
rect 17986 18468 18042 18470
rect 18066 18468 18122 18470
rect 18786 23024 18842 23080
rect 17826 17434 17882 17436
rect 17906 17434 17962 17436
rect 17986 17434 18042 17436
rect 18066 17434 18122 17436
rect 17826 17382 17872 17434
rect 17872 17382 17882 17434
rect 17906 17382 17936 17434
rect 17936 17382 17948 17434
rect 17948 17382 17962 17434
rect 17986 17382 18000 17434
rect 18000 17382 18012 17434
rect 18012 17382 18042 17434
rect 18066 17382 18076 17434
rect 18076 17382 18122 17434
rect 17826 17380 17882 17382
rect 17906 17380 17962 17382
rect 17986 17380 18042 17382
rect 18066 17380 18122 17382
rect 17826 16346 17882 16348
rect 17906 16346 17962 16348
rect 17986 16346 18042 16348
rect 18066 16346 18122 16348
rect 17826 16294 17872 16346
rect 17872 16294 17882 16346
rect 17906 16294 17936 16346
rect 17936 16294 17948 16346
rect 17948 16294 17962 16346
rect 17986 16294 18000 16346
rect 18000 16294 18012 16346
rect 18012 16294 18042 16346
rect 18066 16294 18076 16346
rect 18076 16294 18122 16346
rect 17826 16292 17882 16294
rect 17906 16292 17962 16294
rect 17986 16292 18042 16294
rect 18066 16292 18122 16294
rect 17774 16088 17830 16144
rect 17866 15988 17868 16008
rect 17868 15988 17920 16008
rect 17920 15988 17922 16008
rect 17866 15952 17922 15988
rect 17826 15258 17882 15260
rect 17906 15258 17962 15260
rect 17986 15258 18042 15260
rect 18066 15258 18122 15260
rect 17826 15206 17872 15258
rect 17872 15206 17882 15258
rect 17906 15206 17936 15258
rect 17936 15206 17948 15258
rect 17948 15206 17962 15258
rect 17986 15206 18000 15258
rect 18000 15206 18012 15258
rect 18012 15206 18042 15258
rect 18066 15206 18076 15258
rect 18076 15206 18122 15258
rect 17826 15204 17882 15206
rect 17906 15204 17962 15206
rect 17986 15204 18042 15206
rect 18066 15204 18122 15206
rect 21310 26682 21366 26684
rect 21390 26682 21446 26684
rect 21470 26682 21526 26684
rect 21550 26682 21606 26684
rect 21310 26630 21356 26682
rect 21356 26630 21366 26682
rect 21390 26630 21420 26682
rect 21420 26630 21432 26682
rect 21432 26630 21446 26682
rect 21470 26630 21484 26682
rect 21484 26630 21496 26682
rect 21496 26630 21526 26682
rect 21550 26630 21560 26682
rect 21560 26630 21606 26682
rect 21310 26628 21366 26630
rect 21390 26628 21446 26630
rect 21470 26628 21526 26630
rect 21550 26628 21606 26630
rect 24795 27226 24851 27228
rect 24875 27226 24931 27228
rect 24955 27226 25011 27228
rect 25035 27226 25091 27228
rect 24795 27174 24841 27226
rect 24841 27174 24851 27226
rect 24875 27174 24905 27226
rect 24905 27174 24917 27226
rect 24917 27174 24931 27226
rect 24955 27174 24969 27226
rect 24969 27174 24981 27226
rect 24981 27174 25011 27226
rect 25035 27174 25045 27226
rect 25045 27174 25091 27226
rect 24795 27172 24851 27174
rect 24875 27172 24931 27174
rect 24955 27172 25011 27174
rect 25035 27172 25091 27174
rect 21310 25594 21366 25596
rect 21390 25594 21446 25596
rect 21470 25594 21526 25596
rect 21550 25594 21606 25596
rect 21310 25542 21356 25594
rect 21356 25542 21366 25594
rect 21390 25542 21420 25594
rect 21420 25542 21432 25594
rect 21432 25542 21446 25594
rect 21470 25542 21484 25594
rect 21484 25542 21496 25594
rect 21496 25542 21526 25594
rect 21550 25542 21560 25594
rect 21560 25542 21606 25594
rect 21310 25540 21366 25542
rect 21390 25540 21446 25542
rect 21470 25540 21526 25542
rect 21550 25540 21606 25542
rect 17826 14170 17882 14172
rect 17906 14170 17962 14172
rect 17986 14170 18042 14172
rect 18066 14170 18122 14172
rect 17826 14118 17872 14170
rect 17872 14118 17882 14170
rect 17906 14118 17936 14170
rect 17936 14118 17948 14170
rect 17948 14118 17962 14170
rect 17986 14118 18000 14170
rect 18000 14118 18012 14170
rect 18012 14118 18042 14170
rect 18066 14118 18076 14170
rect 18076 14118 18122 14170
rect 17826 14116 17882 14118
rect 17906 14116 17962 14118
rect 17986 14116 18042 14118
rect 18066 14116 18122 14118
rect 14341 11450 14397 11452
rect 14421 11450 14477 11452
rect 14501 11450 14557 11452
rect 14581 11450 14637 11452
rect 14341 11398 14387 11450
rect 14387 11398 14397 11450
rect 14421 11398 14451 11450
rect 14451 11398 14463 11450
rect 14463 11398 14477 11450
rect 14501 11398 14515 11450
rect 14515 11398 14527 11450
rect 14527 11398 14557 11450
rect 14581 11398 14591 11450
rect 14591 11398 14637 11450
rect 14341 11396 14397 11398
rect 14421 11396 14477 11398
rect 14501 11396 14557 11398
rect 14581 11396 14637 11398
rect 15014 12552 15070 12608
rect 16302 12824 16358 12880
rect 21310 24506 21366 24508
rect 21390 24506 21446 24508
rect 21470 24506 21526 24508
rect 21550 24506 21606 24508
rect 21310 24454 21356 24506
rect 21356 24454 21366 24506
rect 21390 24454 21420 24506
rect 21420 24454 21432 24506
rect 21432 24454 21446 24506
rect 21470 24454 21484 24506
rect 21484 24454 21496 24506
rect 21496 24454 21526 24506
rect 21550 24454 21560 24506
rect 21560 24454 21606 24506
rect 21310 24452 21366 24454
rect 21390 24452 21446 24454
rect 21470 24452 21526 24454
rect 21550 24452 21606 24454
rect 21310 23418 21366 23420
rect 21390 23418 21446 23420
rect 21470 23418 21526 23420
rect 21550 23418 21606 23420
rect 21310 23366 21356 23418
rect 21356 23366 21366 23418
rect 21390 23366 21420 23418
rect 21420 23366 21432 23418
rect 21432 23366 21446 23418
rect 21470 23366 21484 23418
rect 21484 23366 21496 23418
rect 21496 23366 21526 23418
rect 21550 23366 21560 23418
rect 21560 23366 21606 23418
rect 21310 23364 21366 23366
rect 21390 23364 21446 23366
rect 21470 23364 21526 23366
rect 21550 23364 21606 23366
rect 21086 22072 21142 22128
rect 21310 22330 21366 22332
rect 21390 22330 21446 22332
rect 21470 22330 21526 22332
rect 21550 22330 21606 22332
rect 21310 22278 21356 22330
rect 21356 22278 21366 22330
rect 21390 22278 21420 22330
rect 21420 22278 21432 22330
rect 21432 22278 21446 22330
rect 21470 22278 21484 22330
rect 21484 22278 21496 22330
rect 21496 22278 21526 22330
rect 21550 22278 21560 22330
rect 21560 22278 21606 22330
rect 21310 22276 21366 22278
rect 21390 22276 21446 22278
rect 21470 22276 21526 22278
rect 21550 22276 21606 22278
rect 21310 21242 21366 21244
rect 21390 21242 21446 21244
rect 21470 21242 21526 21244
rect 21550 21242 21606 21244
rect 21310 21190 21356 21242
rect 21356 21190 21366 21242
rect 21390 21190 21420 21242
rect 21420 21190 21432 21242
rect 21432 21190 21446 21242
rect 21470 21190 21484 21242
rect 21484 21190 21496 21242
rect 21496 21190 21526 21242
rect 21550 21190 21560 21242
rect 21560 21190 21606 21242
rect 21310 21188 21366 21190
rect 21390 21188 21446 21190
rect 21470 21188 21526 21190
rect 21550 21188 21606 21190
rect 22926 23160 22982 23216
rect 21310 20154 21366 20156
rect 21390 20154 21446 20156
rect 21470 20154 21526 20156
rect 21550 20154 21606 20156
rect 21310 20102 21356 20154
rect 21356 20102 21366 20154
rect 21390 20102 21420 20154
rect 21420 20102 21432 20154
rect 21432 20102 21446 20154
rect 21470 20102 21484 20154
rect 21484 20102 21496 20154
rect 21496 20102 21526 20154
rect 21550 20102 21560 20154
rect 21560 20102 21606 20154
rect 21310 20100 21366 20102
rect 21390 20100 21446 20102
rect 21470 20100 21526 20102
rect 21550 20100 21606 20102
rect 21546 19252 21548 19272
rect 21548 19252 21600 19272
rect 21600 19252 21602 19272
rect 21546 19216 21602 19252
rect 21310 19066 21366 19068
rect 21390 19066 21446 19068
rect 21470 19066 21526 19068
rect 21550 19066 21606 19068
rect 21310 19014 21356 19066
rect 21356 19014 21366 19066
rect 21390 19014 21420 19066
rect 21420 19014 21432 19066
rect 21432 19014 21446 19066
rect 21470 19014 21484 19066
rect 21484 19014 21496 19066
rect 21496 19014 21526 19066
rect 21550 19014 21560 19066
rect 21560 19014 21606 19066
rect 21310 19012 21366 19014
rect 21390 19012 21446 19014
rect 21470 19012 21526 19014
rect 21550 19012 21606 19014
rect 17826 13082 17882 13084
rect 17906 13082 17962 13084
rect 17986 13082 18042 13084
rect 18066 13082 18122 13084
rect 17826 13030 17872 13082
rect 17872 13030 17882 13082
rect 17906 13030 17936 13082
rect 17936 13030 17948 13082
rect 17948 13030 17962 13082
rect 17986 13030 18000 13082
rect 18000 13030 18012 13082
rect 18012 13030 18042 13082
rect 18066 13030 18076 13082
rect 18076 13030 18122 13082
rect 17826 13028 17882 13030
rect 17906 13028 17962 13030
rect 17986 13028 18042 13030
rect 18066 13028 18122 13030
rect 17826 11994 17882 11996
rect 17906 11994 17962 11996
rect 17986 11994 18042 11996
rect 18066 11994 18122 11996
rect 17826 11942 17872 11994
rect 17872 11942 17882 11994
rect 17906 11942 17936 11994
rect 17936 11942 17948 11994
rect 17948 11942 17962 11994
rect 17986 11942 18000 11994
rect 18000 11942 18012 11994
rect 18012 11942 18042 11994
rect 18066 11942 18076 11994
rect 18076 11942 18122 11994
rect 17826 11940 17882 11942
rect 17906 11940 17962 11942
rect 17986 11940 18042 11942
rect 18066 11940 18122 11942
rect 21310 17978 21366 17980
rect 21390 17978 21446 17980
rect 21470 17978 21526 17980
rect 21550 17978 21606 17980
rect 21310 17926 21356 17978
rect 21356 17926 21366 17978
rect 21390 17926 21420 17978
rect 21420 17926 21432 17978
rect 21432 17926 21446 17978
rect 21470 17926 21484 17978
rect 21484 17926 21496 17978
rect 21496 17926 21526 17978
rect 21550 17926 21560 17978
rect 21560 17926 21606 17978
rect 21310 17924 21366 17926
rect 21390 17924 21446 17926
rect 21470 17924 21526 17926
rect 21550 17924 21606 17926
rect 21310 16890 21366 16892
rect 21390 16890 21446 16892
rect 21470 16890 21526 16892
rect 21550 16890 21606 16892
rect 21310 16838 21356 16890
rect 21356 16838 21366 16890
rect 21390 16838 21420 16890
rect 21420 16838 21432 16890
rect 21432 16838 21446 16890
rect 21470 16838 21484 16890
rect 21484 16838 21496 16890
rect 21496 16838 21526 16890
rect 21550 16838 21560 16890
rect 21560 16838 21606 16890
rect 21310 16836 21366 16838
rect 21390 16836 21446 16838
rect 21470 16836 21526 16838
rect 21550 16836 21606 16838
rect 21310 15802 21366 15804
rect 21390 15802 21446 15804
rect 21470 15802 21526 15804
rect 21550 15802 21606 15804
rect 21310 15750 21356 15802
rect 21356 15750 21366 15802
rect 21390 15750 21420 15802
rect 21420 15750 21432 15802
rect 21432 15750 21446 15802
rect 21470 15750 21484 15802
rect 21484 15750 21496 15802
rect 21496 15750 21526 15802
rect 21550 15750 21560 15802
rect 21560 15750 21606 15802
rect 21310 15748 21366 15750
rect 21390 15748 21446 15750
rect 21470 15748 21526 15750
rect 21550 15748 21606 15750
rect 21310 14714 21366 14716
rect 21390 14714 21446 14716
rect 21470 14714 21526 14716
rect 21550 14714 21606 14716
rect 21310 14662 21356 14714
rect 21356 14662 21366 14714
rect 21390 14662 21420 14714
rect 21420 14662 21432 14714
rect 21432 14662 21446 14714
rect 21470 14662 21484 14714
rect 21484 14662 21496 14714
rect 21496 14662 21526 14714
rect 21550 14662 21560 14714
rect 21560 14662 21606 14714
rect 21310 14660 21366 14662
rect 21390 14660 21446 14662
rect 21470 14660 21526 14662
rect 21550 14660 21606 14662
rect 21310 13626 21366 13628
rect 21390 13626 21446 13628
rect 21470 13626 21526 13628
rect 21550 13626 21606 13628
rect 21310 13574 21356 13626
rect 21356 13574 21366 13626
rect 21390 13574 21420 13626
rect 21420 13574 21432 13626
rect 21432 13574 21446 13626
rect 21470 13574 21484 13626
rect 21484 13574 21496 13626
rect 21496 13574 21526 13626
rect 21550 13574 21560 13626
rect 21560 13574 21606 13626
rect 21310 13572 21366 13574
rect 21390 13572 21446 13574
rect 21470 13572 21526 13574
rect 21550 13572 21606 13574
rect 23478 22092 23534 22128
rect 23478 22072 23480 22092
rect 23480 22072 23532 22092
rect 23532 22072 23534 22092
rect 24795 26138 24851 26140
rect 24875 26138 24931 26140
rect 24955 26138 25011 26140
rect 25035 26138 25091 26140
rect 24795 26086 24841 26138
rect 24841 26086 24851 26138
rect 24875 26086 24905 26138
rect 24905 26086 24917 26138
rect 24917 26086 24931 26138
rect 24955 26086 24969 26138
rect 24969 26086 24981 26138
rect 24981 26086 25011 26138
rect 25035 26086 25045 26138
rect 25045 26086 25091 26138
rect 24795 26084 24851 26086
rect 24875 26084 24931 26086
rect 24955 26084 25011 26086
rect 25035 26084 25091 26086
rect 24795 25050 24851 25052
rect 24875 25050 24931 25052
rect 24955 25050 25011 25052
rect 25035 25050 25091 25052
rect 24795 24998 24841 25050
rect 24841 24998 24851 25050
rect 24875 24998 24905 25050
rect 24905 24998 24917 25050
rect 24917 24998 24931 25050
rect 24955 24998 24969 25050
rect 24969 24998 24981 25050
rect 24981 24998 25011 25050
rect 25035 24998 25045 25050
rect 25045 24998 25091 25050
rect 24795 24996 24851 24998
rect 24875 24996 24931 24998
rect 24955 24996 25011 24998
rect 25035 24996 25091 24998
rect 24795 23962 24851 23964
rect 24875 23962 24931 23964
rect 24955 23962 25011 23964
rect 25035 23962 25091 23964
rect 24795 23910 24841 23962
rect 24841 23910 24851 23962
rect 24875 23910 24905 23962
rect 24905 23910 24917 23962
rect 24917 23910 24931 23962
rect 24955 23910 24969 23962
rect 24969 23910 24981 23962
rect 24981 23910 25011 23962
rect 25035 23910 25045 23962
rect 25045 23910 25091 23962
rect 24795 23908 24851 23910
rect 24875 23908 24931 23910
rect 24955 23908 25011 23910
rect 25035 23908 25091 23910
rect 24795 22874 24851 22876
rect 24875 22874 24931 22876
rect 24955 22874 25011 22876
rect 25035 22874 25091 22876
rect 24795 22822 24841 22874
rect 24841 22822 24851 22874
rect 24875 22822 24905 22874
rect 24905 22822 24917 22874
rect 24917 22822 24931 22874
rect 24955 22822 24969 22874
rect 24969 22822 24981 22874
rect 24981 22822 25011 22874
rect 25035 22822 25045 22874
rect 25045 22822 25091 22874
rect 24795 22820 24851 22822
rect 24875 22820 24931 22822
rect 24955 22820 25011 22822
rect 25035 22820 25091 22822
rect 24795 21786 24851 21788
rect 24875 21786 24931 21788
rect 24955 21786 25011 21788
rect 25035 21786 25091 21788
rect 24795 21734 24841 21786
rect 24841 21734 24851 21786
rect 24875 21734 24905 21786
rect 24905 21734 24917 21786
rect 24917 21734 24931 21786
rect 24955 21734 24969 21786
rect 24969 21734 24981 21786
rect 24981 21734 25011 21786
rect 25035 21734 25045 21786
rect 25045 21734 25091 21786
rect 24795 21732 24851 21734
rect 24875 21732 24931 21734
rect 24955 21732 25011 21734
rect 25035 21732 25091 21734
rect 24795 20698 24851 20700
rect 24875 20698 24931 20700
rect 24955 20698 25011 20700
rect 25035 20698 25091 20700
rect 24795 20646 24841 20698
rect 24841 20646 24851 20698
rect 24875 20646 24905 20698
rect 24905 20646 24917 20698
rect 24917 20646 24931 20698
rect 24955 20646 24969 20698
rect 24969 20646 24981 20698
rect 24981 20646 25011 20698
rect 25035 20646 25045 20698
rect 25045 20646 25091 20698
rect 24795 20644 24851 20646
rect 24875 20644 24931 20646
rect 24955 20644 25011 20646
rect 25035 20644 25091 20646
rect 24795 19610 24851 19612
rect 24875 19610 24931 19612
rect 24955 19610 25011 19612
rect 25035 19610 25091 19612
rect 24795 19558 24841 19610
rect 24841 19558 24851 19610
rect 24875 19558 24905 19610
rect 24905 19558 24917 19610
rect 24917 19558 24931 19610
rect 24955 19558 24969 19610
rect 24969 19558 24981 19610
rect 24981 19558 25011 19610
rect 25035 19558 25045 19610
rect 25045 19558 25091 19610
rect 24795 19556 24851 19558
rect 24875 19556 24931 19558
rect 24955 19556 25011 19558
rect 25035 19556 25091 19558
rect 28279 27770 28335 27772
rect 28359 27770 28415 27772
rect 28439 27770 28495 27772
rect 28519 27770 28575 27772
rect 28279 27718 28325 27770
rect 28325 27718 28335 27770
rect 28359 27718 28389 27770
rect 28389 27718 28401 27770
rect 28401 27718 28415 27770
rect 28439 27718 28453 27770
rect 28453 27718 28465 27770
rect 28465 27718 28495 27770
rect 28519 27718 28529 27770
rect 28529 27718 28575 27770
rect 28279 27716 28335 27718
rect 28359 27716 28415 27718
rect 28439 27716 28495 27718
rect 28519 27716 28575 27718
rect 28279 26682 28335 26684
rect 28359 26682 28415 26684
rect 28439 26682 28495 26684
rect 28519 26682 28575 26684
rect 28279 26630 28325 26682
rect 28325 26630 28335 26682
rect 28359 26630 28389 26682
rect 28389 26630 28401 26682
rect 28401 26630 28415 26682
rect 28439 26630 28453 26682
rect 28453 26630 28465 26682
rect 28465 26630 28495 26682
rect 28519 26630 28529 26682
rect 28529 26630 28575 26682
rect 28279 26628 28335 26630
rect 28359 26628 28415 26630
rect 28439 26628 28495 26630
rect 28519 26628 28575 26630
rect 28279 25594 28335 25596
rect 28359 25594 28415 25596
rect 28439 25594 28495 25596
rect 28519 25594 28575 25596
rect 28279 25542 28325 25594
rect 28325 25542 28335 25594
rect 28359 25542 28389 25594
rect 28389 25542 28401 25594
rect 28401 25542 28415 25594
rect 28439 25542 28453 25594
rect 28453 25542 28465 25594
rect 28465 25542 28495 25594
rect 28519 25542 28529 25594
rect 28529 25542 28575 25594
rect 28279 25540 28335 25542
rect 28359 25540 28415 25542
rect 28439 25540 28495 25542
rect 28519 25540 28575 25542
rect 28279 24506 28335 24508
rect 28359 24506 28415 24508
rect 28439 24506 28495 24508
rect 28519 24506 28575 24508
rect 28279 24454 28325 24506
rect 28325 24454 28335 24506
rect 28359 24454 28389 24506
rect 28389 24454 28401 24506
rect 28401 24454 28415 24506
rect 28439 24454 28453 24506
rect 28453 24454 28465 24506
rect 28465 24454 28495 24506
rect 28519 24454 28529 24506
rect 28529 24454 28575 24506
rect 28279 24452 28335 24454
rect 28359 24452 28415 24454
rect 28439 24452 28495 24454
rect 28519 24452 28575 24454
rect 28279 23418 28335 23420
rect 28359 23418 28415 23420
rect 28439 23418 28495 23420
rect 28519 23418 28575 23420
rect 28279 23366 28325 23418
rect 28325 23366 28335 23418
rect 28359 23366 28389 23418
rect 28389 23366 28401 23418
rect 28401 23366 28415 23418
rect 28439 23366 28453 23418
rect 28453 23366 28465 23418
rect 28465 23366 28495 23418
rect 28519 23366 28529 23418
rect 28529 23366 28575 23418
rect 28279 23364 28335 23366
rect 28359 23364 28415 23366
rect 28439 23364 28495 23366
rect 28519 23364 28575 23366
rect 28279 22330 28335 22332
rect 28359 22330 28415 22332
rect 28439 22330 28495 22332
rect 28519 22330 28575 22332
rect 28279 22278 28325 22330
rect 28325 22278 28335 22330
rect 28359 22278 28389 22330
rect 28389 22278 28401 22330
rect 28401 22278 28415 22330
rect 28439 22278 28453 22330
rect 28453 22278 28465 22330
rect 28465 22278 28495 22330
rect 28519 22278 28529 22330
rect 28529 22278 28575 22330
rect 28279 22276 28335 22278
rect 28359 22276 28415 22278
rect 28439 22276 28495 22278
rect 28519 22276 28575 22278
rect 28279 21242 28335 21244
rect 28359 21242 28415 21244
rect 28439 21242 28495 21244
rect 28519 21242 28575 21244
rect 28279 21190 28325 21242
rect 28325 21190 28335 21242
rect 28359 21190 28389 21242
rect 28389 21190 28401 21242
rect 28401 21190 28415 21242
rect 28439 21190 28453 21242
rect 28453 21190 28465 21242
rect 28465 21190 28495 21242
rect 28519 21190 28529 21242
rect 28529 21190 28575 21242
rect 28279 21188 28335 21190
rect 28359 21188 28415 21190
rect 28439 21188 28495 21190
rect 28519 21188 28575 21190
rect 28279 20154 28335 20156
rect 28359 20154 28415 20156
rect 28439 20154 28495 20156
rect 28519 20154 28575 20156
rect 28279 20102 28325 20154
rect 28325 20102 28335 20154
rect 28359 20102 28389 20154
rect 28389 20102 28401 20154
rect 28401 20102 28415 20154
rect 28439 20102 28453 20154
rect 28453 20102 28465 20154
rect 28465 20102 28495 20154
rect 28519 20102 28529 20154
rect 28529 20102 28575 20154
rect 28279 20100 28335 20102
rect 28359 20100 28415 20102
rect 28439 20100 28495 20102
rect 28519 20100 28575 20102
rect 27618 19216 27674 19272
rect 28279 19066 28335 19068
rect 28359 19066 28415 19068
rect 28439 19066 28495 19068
rect 28519 19066 28575 19068
rect 28279 19014 28325 19066
rect 28325 19014 28335 19066
rect 28359 19014 28389 19066
rect 28389 19014 28401 19066
rect 28401 19014 28415 19066
rect 28439 19014 28453 19066
rect 28453 19014 28465 19066
rect 28465 19014 28495 19066
rect 28519 19014 28529 19066
rect 28529 19014 28575 19066
rect 28279 19012 28335 19014
rect 28359 19012 28415 19014
rect 28439 19012 28495 19014
rect 28519 19012 28575 19014
rect 24795 18522 24851 18524
rect 24875 18522 24931 18524
rect 24955 18522 25011 18524
rect 25035 18522 25091 18524
rect 24795 18470 24841 18522
rect 24841 18470 24851 18522
rect 24875 18470 24905 18522
rect 24905 18470 24917 18522
rect 24917 18470 24931 18522
rect 24955 18470 24969 18522
rect 24969 18470 24981 18522
rect 24981 18470 25011 18522
rect 25035 18470 25045 18522
rect 25045 18470 25091 18522
rect 24795 18468 24851 18470
rect 24875 18468 24931 18470
rect 24955 18468 25011 18470
rect 25035 18468 25091 18470
rect 28279 17978 28335 17980
rect 28359 17978 28415 17980
rect 28439 17978 28495 17980
rect 28519 17978 28575 17980
rect 28279 17926 28325 17978
rect 28325 17926 28335 17978
rect 28359 17926 28389 17978
rect 28389 17926 28401 17978
rect 28401 17926 28415 17978
rect 28439 17926 28453 17978
rect 28453 17926 28465 17978
rect 28465 17926 28495 17978
rect 28519 17926 28529 17978
rect 28529 17926 28575 17978
rect 28279 17924 28335 17926
rect 28359 17924 28415 17926
rect 28439 17924 28495 17926
rect 28519 17924 28575 17926
rect 24795 17434 24851 17436
rect 24875 17434 24931 17436
rect 24955 17434 25011 17436
rect 25035 17434 25091 17436
rect 24795 17382 24841 17434
rect 24841 17382 24851 17434
rect 24875 17382 24905 17434
rect 24905 17382 24917 17434
rect 24917 17382 24931 17434
rect 24955 17382 24969 17434
rect 24969 17382 24981 17434
rect 24981 17382 25011 17434
rect 25035 17382 25045 17434
rect 25045 17382 25091 17434
rect 24795 17380 24851 17382
rect 24875 17380 24931 17382
rect 24955 17380 25011 17382
rect 25035 17380 25091 17382
rect 28279 16890 28335 16892
rect 28359 16890 28415 16892
rect 28439 16890 28495 16892
rect 28519 16890 28575 16892
rect 28279 16838 28325 16890
rect 28325 16838 28335 16890
rect 28359 16838 28389 16890
rect 28389 16838 28401 16890
rect 28401 16838 28415 16890
rect 28439 16838 28453 16890
rect 28453 16838 28465 16890
rect 28465 16838 28495 16890
rect 28519 16838 28529 16890
rect 28529 16838 28575 16890
rect 28279 16836 28335 16838
rect 28359 16836 28415 16838
rect 28439 16836 28495 16838
rect 28519 16836 28575 16838
rect 24795 16346 24851 16348
rect 24875 16346 24931 16348
rect 24955 16346 25011 16348
rect 25035 16346 25091 16348
rect 24795 16294 24841 16346
rect 24841 16294 24851 16346
rect 24875 16294 24905 16346
rect 24905 16294 24917 16346
rect 24917 16294 24931 16346
rect 24955 16294 24969 16346
rect 24969 16294 24981 16346
rect 24981 16294 25011 16346
rect 25035 16294 25045 16346
rect 25045 16294 25091 16346
rect 24795 16292 24851 16294
rect 24875 16292 24931 16294
rect 24955 16292 25011 16294
rect 25035 16292 25091 16294
rect 28279 15802 28335 15804
rect 28359 15802 28415 15804
rect 28439 15802 28495 15804
rect 28519 15802 28575 15804
rect 28279 15750 28325 15802
rect 28325 15750 28335 15802
rect 28359 15750 28389 15802
rect 28389 15750 28401 15802
rect 28401 15750 28415 15802
rect 28439 15750 28453 15802
rect 28453 15750 28465 15802
rect 28465 15750 28495 15802
rect 28519 15750 28529 15802
rect 28529 15750 28575 15802
rect 28279 15748 28335 15750
rect 28359 15748 28415 15750
rect 28439 15748 28495 15750
rect 28519 15748 28575 15750
rect 24795 15258 24851 15260
rect 24875 15258 24931 15260
rect 24955 15258 25011 15260
rect 25035 15258 25091 15260
rect 24795 15206 24841 15258
rect 24841 15206 24851 15258
rect 24875 15206 24905 15258
rect 24905 15206 24917 15258
rect 24917 15206 24931 15258
rect 24955 15206 24969 15258
rect 24969 15206 24981 15258
rect 24981 15206 25011 15258
rect 25035 15206 25045 15258
rect 25045 15206 25091 15258
rect 24795 15204 24851 15206
rect 24875 15204 24931 15206
rect 24955 15204 25011 15206
rect 25035 15204 25091 15206
rect 28279 14714 28335 14716
rect 28359 14714 28415 14716
rect 28439 14714 28495 14716
rect 28519 14714 28575 14716
rect 28279 14662 28325 14714
rect 28325 14662 28335 14714
rect 28359 14662 28389 14714
rect 28389 14662 28401 14714
rect 28401 14662 28415 14714
rect 28439 14662 28453 14714
rect 28453 14662 28465 14714
rect 28465 14662 28495 14714
rect 28519 14662 28529 14714
rect 28529 14662 28575 14714
rect 28279 14660 28335 14662
rect 28359 14660 28415 14662
rect 28439 14660 28495 14662
rect 28519 14660 28575 14662
rect 24795 14170 24851 14172
rect 24875 14170 24931 14172
rect 24955 14170 25011 14172
rect 25035 14170 25091 14172
rect 24795 14118 24841 14170
rect 24841 14118 24851 14170
rect 24875 14118 24905 14170
rect 24905 14118 24917 14170
rect 24917 14118 24931 14170
rect 24955 14118 24969 14170
rect 24969 14118 24981 14170
rect 24981 14118 25011 14170
rect 25035 14118 25045 14170
rect 25045 14118 25091 14170
rect 24795 14116 24851 14118
rect 24875 14116 24931 14118
rect 24955 14116 25011 14118
rect 25035 14116 25091 14118
rect 21310 12538 21366 12540
rect 21390 12538 21446 12540
rect 21470 12538 21526 12540
rect 21550 12538 21606 12540
rect 21310 12486 21356 12538
rect 21356 12486 21366 12538
rect 21390 12486 21420 12538
rect 21420 12486 21432 12538
rect 21432 12486 21446 12538
rect 21470 12486 21484 12538
rect 21484 12486 21496 12538
rect 21496 12486 21526 12538
rect 21550 12486 21560 12538
rect 21560 12486 21606 12538
rect 21310 12484 21366 12486
rect 21390 12484 21446 12486
rect 21470 12484 21526 12486
rect 21550 12484 21606 12486
rect 28279 13626 28335 13628
rect 28359 13626 28415 13628
rect 28439 13626 28495 13628
rect 28519 13626 28575 13628
rect 28279 13574 28325 13626
rect 28325 13574 28335 13626
rect 28359 13574 28389 13626
rect 28389 13574 28401 13626
rect 28401 13574 28415 13626
rect 28439 13574 28453 13626
rect 28453 13574 28465 13626
rect 28465 13574 28495 13626
rect 28519 13574 28529 13626
rect 28529 13574 28575 13626
rect 28279 13572 28335 13574
rect 28359 13572 28415 13574
rect 28439 13572 28495 13574
rect 28519 13572 28575 13574
rect 24795 13082 24851 13084
rect 24875 13082 24931 13084
rect 24955 13082 25011 13084
rect 25035 13082 25091 13084
rect 24795 13030 24841 13082
rect 24841 13030 24851 13082
rect 24875 13030 24905 13082
rect 24905 13030 24917 13082
rect 24917 13030 24931 13082
rect 24955 13030 24969 13082
rect 24969 13030 24981 13082
rect 24981 13030 25011 13082
rect 25035 13030 25045 13082
rect 25045 13030 25091 13082
rect 24795 13028 24851 13030
rect 24875 13028 24931 13030
rect 24955 13028 25011 13030
rect 25035 13028 25091 13030
rect 28279 12538 28335 12540
rect 28359 12538 28415 12540
rect 28439 12538 28495 12540
rect 28519 12538 28575 12540
rect 28279 12486 28325 12538
rect 28325 12486 28335 12538
rect 28359 12486 28389 12538
rect 28389 12486 28401 12538
rect 28401 12486 28415 12538
rect 28439 12486 28453 12538
rect 28453 12486 28465 12538
rect 28465 12486 28495 12538
rect 28519 12486 28529 12538
rect 28529 12486 28575 12538
rect 28279 12484 28335 12486
rect 28359 12484 28415 12486
rect 28439 12484 28495 12486
rect 28519 12484 28575 12486
rect 24795 11994 24851 11996
rect 24875 11994 24931 11996
rect 24955 11994 25011 11996
rect 25035 11994 25091 11996
rect 24795 11942 24841 11994
rect 24841 11942 24851 11994
rect 24875 11942 24905 11994
rect 24905 11942 24917 11994
rect 24917 11942 24931 11994
rect 24955 11942 24969 11994
rect 24969 11942 24981 11994
rect 24981 11942 25011 11994
rect 25035 11942 25045 11994
rect 25045 11942 25091 11994
rect 24795 11940 24851 11942
rect 24875 11940 24931 11942
rect 24955 11940 25011 11942
rect 25035 11940 25091 11942
rect 21310 11450 21366 11452
rect 21390 11450 21446 11452
rect 21470 11450 21526 11452
rect 21550 11450 21606 11452
rect 21310 11398 21356 11450
rect 21356 11398 21366 11450
rect 21390 11398 21420 11450
rect 21420 11398 21432 11450
rect 21432 11398 21446 11450
rect 21470 11398 21484 11450
rect 21484 11398 21496 11450
rect 21496 11398 21526 11450
rect 21550 11398 21560 11450
rect 21560 11398 21606 11450
rect 21310 11396 21366 11398
rect 21390 11396 21446 11398
rect 21470 11396 21526 11398
rect 21550 11396 21606 11398
rect 28279 11450 28335 11452
rect 28359 11450 28415 11452
rect 28439 11450 28495 11452
rect 28519 11450 28575 11452
rect 28279 11398 28325 11450
rect 28325 11398 28335 11450
rect 28359 11398 28389 11450
rect 28389 11398 28401 11450
rect 28401 11398 28415 11450
rect 28439 11398 28453 11450
rect 28453 11398 28465 11450
rect 28465 11398 28495 11450
rect 28519 11398 28529 11450
rect 28529 11398 28575 11450
rect 28279 11396 28335 11398
rect 28359 11396 28415 11398
rect 28439 11396 28495 11398
rect 28519 11396 28575 11398
rect 17826 10906 17882 10908
rect 17906 10906 17962 10908
rect 17986 10906 18042 10908
rect 18066 10906 18122 10908
rect 17826 10854 17872 10906
rect 17872 10854 17882 10906
rect 17906 10854 17936 10906
rect 17936 10854 17948 10906
rect 17948 10854 17962 10906
rect 17986 10854 18000 10906
rect 18000 10854 18012 10906
rect 18012 10854 18042 10906
rect 18066 10854 18076 10906
rect 18076 10854 18122 10906
rect 17826 10852 17882 10854
rect 17906 10852 17962 10854
rect 17986 10852 18042 10854
rect 18066 10852 18122 10854
rect 24795 10906 24851 10908
rect 24875 10906 24931 10908
rect 24955 10906 25011 10908
rect 25035 10906 25091 10908
rect 24795 10854 24841 10906
rect 24841 10854 24851 10906
rect 24875 10854 24905 10906
rect 24905 10854 24917 10906
rect 24917 10854 24931 10906
rect 24955 10854 24969 10906
rect 24969 10854 24981 10906
rect 24981 10854 25011 10906
rect 25035 10854 25045 10906
rect 25045 10854 25091 10906
rect 24795 10852 24851 10854
rect 24875 10852 24931 10854
rect 24955 10852 25011 10854
rect 25035 10852 25091 10854
rect 14341 10362 14397 10364
rect 14421 10362 14477 10364
rect 14501 10362 14557 10364
rect 14581 10362 14637 10364
rect 14341 10310 14387 10362
rect 14387 10310 14397 10362
rect 14421 10310 14451 10362
rect 14451 10310 14463 10362
rect 14463 10310 14477 10362
rect 14501 10310 14515 10362
rect 14515 10310 14527 10362
rect 14527 10310 14557 10362
rect 14581 10310 14591 10362
rect 14591 10310 14637 10362
rect 14341 10308 14397 10310
rect 14421 10308 14477 10310
rect 14501 10308 14557 10310
rect 14581 10308 14637 10310
rect 21310 10362 21366 10364
rect 21390 10362 21446 10364
rect 21470 10362 21526 10364
rect 21550 10362 21606 10364
rect 21310 10310 21356 10362
rect 21356 10310 21366 10362
rect 21390 10310 21420 10362
rect 21420 10310 21432 10362
rect 21432 10310 21446 10362
rect 21470 10310 21484 10362
rect 21484 10310 21496 10362
rect 21496 10310 21526 10362
rect 21550 10310 21560 10362
rect 21560 10310 21606 10362
rect 21310 10308 21366 10310
rect 21390 10308 21446 10310
rect 21470 10308 21526 10310
rect 21550 10308 21606 10310
rect 28279 10362 28335 10364
rect 28359 10362 28415 10364
rect 28439 10362 28495 10364
rect 28519 10362 28575 10364
rect 28279 10310 28325 10362
rect 28325 10310 28335 10362
rect 28359 10310 28389 10362
rect 28389 10310 28401 10362
rect 28401 10310 28415 10362
rect 28439 10310 28453 10362
rect 28453 10310 28465 10362
rect 28465 10310 28495 10362
rect 28519 10310 28529 10362
rect 28529 10310 28575 10362
rect 28279 10308 28335 10310
rect 28359 10308 28415 10310
rect 28439 10308 28495 10310
rect 28519 10308 28575 10310
rect 3888 9818 3944 9820
rect 3968 9818 4024 9820
rect 4048 9818 4104 9820
rect 4128 9818 4184 9820
rect 3888 9766 3934 9818
rect 3934 9766 3944 9818
rect 3968 9766 3998 9818
rect 3998 9766 4010 9818
rect 4010 9766 4024 9818
rect 4048 9766 4062 9818
rect 4062 9766 4074 9818
rect 4074 9766 4104 9818
rect 4128 9766 4138 9818
rect 4138 9766 4184 9818
rect 3888 9764 3944 9766
rect 3968 9764 4024 9766
rect 4048 9764 4104 9766
rect 4128 9764 4184 9766
rect 10857 9818 10913 9820
rect 10937 9818 10993 9820
rect 11017 9818 11073 9820
rect 11097 9818 11153 9820
rect 10857 9766 10903 9818
rect 10903 9766 10913 9818
rect 10937 9766 10967 9818
rect 10967 9766 10979 9818
rect 10979 9766 10993 9818
rect 11017 9766 11031 9818
rect 11031 9766 11043 9818
rect 11043 9766 11073 9818
rect 11097 9766 11107 9818
rect 11107 9766 11153 9818
rect 10857 9764 10913 9766
rect 10937 9764 10993 9766
rect 11017 9764 11073 9766
rect 11097 9764 11153 9766
rect 17826 9818 17882 9820
rect 17906 9818 17962 9820
rect 17986 9818 18042 9820
rect 18066 9818 18122 9820
rect 17826 9766 17872 9818
rect 17872 9766 17882 9818
rect 17906 9766 17936 9818
rect 17936 9766 17948 9818
rect 17948 9766 17962 9818
rect 17986 9766 18000 9818
rect 18000 9766 18012 9818
rect 18012 9766 18042 9818
rect 18066 9766 18076 9818
rect 18076 9766 18122 9818
rect 17826 9764 17882 9766
rect 17906 9764 17962 9766
rect 17986 9764 18042 9766
rect 18066 9764 18122 9766
rect 24795 9818 24851 9820
rect 24875 9818 24931 9820
rect 24955 9818 25011 9820
rect 25035 9818 25091 9820
rect 24795 9766 24841 9818
rect 24841 9766 24851 9818
rect 24875 9766 24905 9818
rect 24905 9766 24917 9818
rect 24917 9766 24931 9818
rect 24955 9766 24969 9818
rect 24969 9766 24981 9818
rect 24981 9766 25011 9818
rect 25035 9766 25045 9818
rect 25045 9766 25091 9818
rect 24795 9764 24851 9766
rect 24875 9764 24931 9766
rect 24955 9764 25011 9766
rect 25035 9764 25091 9766
rect 7372 9274 7428 9276
rect 7452 9274 7508 9276
rect 7532 9274 7588 9276
rect 7612 9274 7668 9276
rect 7372 9222 7418 9274
rect 7418 9222 7428 9274
rect 7452 9222 7482 9274
rect 7482 9222 7494 9274
rect 7494 9222 7508 9274
rect 7532 9222 7546 9274
rect 7546 9222 7558 9274
rect 7558 9222 7588 9274
rect 7612 9222 7622 9274
rect 7622 9222 7668 9274
rect 7372 9220 7428 9222
rect 7452 9220 7508 9222
rect 7532 9220 7588 9222
rect 7612 9220 7668 9222
rect 14341 9274 14397 9276
rect 14421 9274 14477 9276
rect 14501 9274 14557 9276
rect 14581 9274 14637 9276
rect 14341 9222 14387 9274
rect 14387 9222 14397 9274
rect 14421 9222 14451 9274
rect 14451 9222 14463 9274
rect 14463 9222 14477 9274
rect 14501 9222 14515 9274
rect 14515 9222 14527 9274
rect 14527 9222 14557 9274
rect 14581 9222 14591 9274
rect 14591 9222 14637 9274
rect 14341 9220 14397 9222
rect 14421 9220 14477 9222
rect 14501 9220 14557 9222
rect 14581 9220 14637 9222
rect 21310 9274 21366 9276
rect 21390 9274 21446 9276
rect 21470 9274 21526 9276
rect 21550 9274 21606 9276
rect 21310 9222 21356 9274
rect 21356 9222 21366 9274
rect 21390 9222 21420 9274
rect 21420 9222 21432 9274
rect 21432 9222 21446 9274
rect 21470 9222 21484 9274
rect 21484 9222 21496 9274
rect 21496 9222 21526 9274
rect 21550 9222 21560 9274
rect 21560 9222 21606 9274
rect 21310 9220 21366 9222
rect 21390 9220 21446 9222
rect 21470 9220 21526 9222
rect 21550 9220 21606 9222
rect 28279 9274 28335 9276
rect 28359 9274 28415 9276
rect 28439 9274 28495 9276
rect 28519 9274 28575 9276
rect 28279 9222 28325 9274
rect 28325 9222 28335 9274
rect 28359 9222 28389 9274
rect 28389 9222 28401 9274
rect 28401 9222 28415 9274
rect 28439 9222 28453 9274
rect 28453 9222 28465 9274
rect 28465 9222 28495 9274
rect 28519 9222 28529 9274
rect 28529 9222 28575 9274
rect 28279 9220 28335 9222
rect 28359 9220 28415 9222
rect 28439 9220 28495 9222
rect 28519 9220 28575 9222
rect 3888 8730 3944 8732
rect 3968 8730 4024 8732
rect 4048 8730 4104 8732
rect 4128 8730 4184 8732
rect 3888 8678 3934 8730
rect 3934 8678 3944 8730
rect 3968 8678 3998 8730
rect 3998 8678 4010 8730
rect 4010 8678 4024 8730
rect 4048 8678 4062 8730
rect 4062 8678 4074 8730
rect 4074 8678 4104 8730
rect 4128 8678 4138 8730
rect 4138 8678 4184 8730
rect 3888 8676 3944 8678
rect 3968 8676 4024 8678
rect 4048 8676 4104 8678
rect 4128 8676 4184 8678
rect 10857 8730 10913 8732
rect 10937 8730 10993 8732
rect 11017 8730 11073 8732
rect 11097 8730 11153 8732
rect 10857 8678 10903 8730
rect 10903 8678 10913 8730
rect 10937 8678 10967 8730
rect 10967 8678 10979 8730
rect 10979 8678 10993 8730
rect 11017 8678 11031 8730
rect 11031 8678 11043 8730
rect 11043 8678 11073 8730
rect 11097 8678 11107 8730
rect 11107 8678 11153 8730
rect 10857 8676 10913 8678
rect 10937 8676 10993 8678
rect 11017 8676 11073 8678
rect 11097 8676 11153 8678
rect 17826 8730 17882 8732
rect 17906 8730 17962 8732
rect 17986 8730 18042 8732
rect 18066 8730 18122 8732
rect 17826 8678 17872 8730
rect 17872 8678 17882 8730
rect 17906 8678 17936 8730
rect 17936 8678 17948 8730
rect 17948 8678 17962 8730
rect 17986 8678 18000 8730
rect 18000 8678 18012 8730
rect 18012 8678 18042 8730
rect 18066 8678 18076 8730
rect 18076 8678 18122 8730
rect 17826 8676 17882 8678
rect 17906 8676 17962 8678
rect 17986 8676 18042 8678
rect 18066 8676 18122 8678
rect 24795 8730 24851 8732
rect 24875 8730 24931 8732
rect 24955 8730 25011 8732
rect 25035 8730 25091 8732
rect 24795 8678 24841 8730
rect 24841 8678 24851 8730
rect 24875 8678 24905 8730
rect 24905 8678 24917 8730
rect 24917 8678 24931 8730
rect 24955 8678 24969 8730
rect 24969 8678 24981 8730
rect 24981 8678 25011 8730
rect 25035 8678 25045 8730
rect 25045 8678 25091 8730
rect 24795 8676 24851 8678
rect 24875 8676 24931 8678
rect 24955 8676 25011 8678
rect 25035 8676 25091 8678
rect 7372 8186 7428 8188
rect 7452 8186 7508 8188
rect 7532 8186 7588 8188
rect 7612 8186 7668 8188
rect 7372 8134 7418 8186
rect 7418 8134 7428 8186
rect 7452 8134 7482 8186
rect 7482 8134 7494 8186
rect 7494 8134 7508 8186
rect 7532 8134 7546 8186
rect 7546 8134 7558 8186
rect 7558 8134 7588 8186
rect 7612 8134 7622 8186
rect 7622 8134 7668 8186
rect 7372 8132 7428 8134
rect 7452 8132 7508 8134
rect 7532 8132 7588 8134
rect 7612 8132 7668 8134
rect 14341 8186 14397 8188
rect 14421 8186 14477 8188
rect 14501 8186 14557 8188
rect 14581 8186 14637 8188
rect 14341 8134 14387 8186
rect 14387 8134 14397 8186
rect 14421 8134 14451 8186
rect 14451 8134 14463 8186
rect 14463 8134 14477 8186
rect 14501 8134 14515 8186
rect 14515 8134 14527 8186
rect 14527 8134 14557 8186
rect 14581 8134 14591 8186
rect 14591 8134 14637 8186
rect 14341 8132 14397 8134
rect 14421 8132 14477 8134
rect 14501 8132 14557 8134
rect 14581 8132 14637 8134
rect 21310 8186 21366 8188
rect 21390 8186 21446 8188
rect 21470 8186 21526 8188
rect 21550 8186 21606 8188
rect 21310 8134 21356 8186
rect 21356 8134 21366 8186
rect 21390 8134 21420 8186
rect 21420 8134 21432 8186
rect 21432 8134 21446 8186
rect 21470 8134 21484 8186
rect 21484 8134 21496 8186
rect 21496 8134 21526 8186
rect 21550 8134 21560 8186
rect 21560 8134 21606 8186
rect 21310 8132 21366 8134
rect 21390 8132 21446 8134
rect 21470 8132 21526 8134
rect 21550 8132 21606 8134
rect 28279 8186 28335 8188
rect 28359 8186 28415 8188
rect 28439 8186 28495 8188
rect 28519 8186 28575 8188
rect 28279 8134 28325 8186
rect 28325 8134 28335 8186
rect 28359 8134 28389 8186
rect 28389 8134 28401 8186
rect 28401 8134 28415 8186
rect 28439 8134 28453 8186
rect 28453 8134 28465 8186
rect 28465 8134 28495 8186
rect 28519 8134 28529 8186
rect 28529 8134 28575 8186
rect 28279 8132 28335 8134
rect 28359 8132 28415 8134
rect 28439 8132 28495 8134
rect 28519 8132 28575 8134
rect 3888 7642 3944 7644
rect 3968 7642 4024 7644
rect 4048 7642 4104 7644
rect 4128 7642 4184 7644
rect 3888 7590 3934 7642
rect 3934 7590 3944 7642
rect 3968 7590 3998 7642
rect 3998 7590 4010 7642
rect 4010 7590 4024 7642
rect 4048 7590 4062 7642
rect 4062 7590 4074 7642
rect 4074 7590 4104 7642
rect 4128 7590 4138 7642
rect 4138 7590 4184 7642
rect 3888 7588 3944 7590
rect 3968 7588 4024 7590
rect 4048 7588 4104 7590
rect 4128 7588 4184 7590
rect 10857 7642 10913 7644
rect 10937 7642 10993 7644
rect 11017 7642 11073 7644
rect 11097 7642 11153 7644
rect 10857 7590 10903 7642
rect 10903 7590 10913 7642
rect 10937 7590 10967 7642
rect 10967 7590 10979 7642
rect 10979 7590 10993 7642
rect 11017 7590 11031 7642
rect 11031 7590 11043 7642
rect 11043 7590 11073 7642
rect 11097 7590 11107 7642
rect 11107 7590 11153 7642
rect 10857 7588 10913 7590
rect 10937 7588 10993 7590
rect 11017 7588 11073 7590
rect 11097 7588 11153 7590
rect 17826 7642 17882 7644
rect 17906 7642 17962 7644
rect 17986 7642 18042 7644
rect 18066 7642 18122 7644
rect 17826 7590 17872 7642
rect 17872 7590 17882 7642
rect 17906 7590 17936 7642
rect 17936 7590 17948 7642
rect 17948 7590 17962 7642
rect 17986 7590 18000 7642
rect 18000 7590 18012 7642
rect 18012 7590 18042 7642
rect 18066 7590 18076 7642
rect 18076 7590 18122 7642
rect 17826 7588 17882 7590
rect 17906 7588 17962 7590
rect 17986 7588 18042 7590
rect 18066 7588 18122 7590
rect 24795 7642 24851 7644
rect 24875 7642 24931 7644
rect 24955 7642 25011 7644
rect 25035 7642 25091 7644
rect 24795 7590 24841 7642
rect 24841 7590 24851 7642
rect 24875 7590 24905 7642
rect 24905 7590 24917 7642
rect 24917 7590 24931 7642
rect 24955 7590 24969 7642
rect 24969 7590 24981 7642
rect 24981 7590 25011 7642
rect 25035 7590 25045 7642
rect 25045 7590 25091 7642
rect 24795 7588 24851 7590
rect 24875 7588 24931 7590
rect 24955 7588 25011 7590
rect 25035 7588 25091 7590
rect 7372 7098 7428 7100
rect 7452 7098 7508 7100
rect 7532 7098 7588 7100
rect 7612 7098 7668 7100
rect 7372 7046 7418 7098
rect 7418 7046 7428 7098
rect 7452 7046 7482 7098
rect 7482 7046 7494 7098
rect 7494 7046 7508 7098
rect 7532 7046 7546 7098
rect 7546 7046 7558 7098
rect 7558 7046 7588 7098
rect 7612 7046 7622 7098
rect 7622 7046 7668 7098
rect 7372 7044 7428 7046
rect 7452 7044 7508 7046
rect 7532 7044 7588 7046
rect 7612 7044 7668 7046
rect 14341 7098 14397 7100
rect 14421 7098 14477 7100
rect 14501 7098 14557 7100
rect 14581 7098 14637 7100
rect 14341 7046 14387 7098
rect 14387 7046 14397 7098
rect 14421 7046 14451 7098
rect 14451 7046 14463 7098
rect 14463 7046 14477 7098
rect 14501 7046 14515 7098
rect 14515 7046 14527 7098
rect 14527 7046 14557 7098
rect 14581 7046 14591 7098
rect 14591 7046 14637 7098
rect 14341 7044 14397 7046
rect 14421 7044 14477 7046
rect 14501 7044 14557 7046
rect 14581 7044 14637 7046
rect 21310 7098 21366 7100
rect 21390 7098 21446 7100
rect 21470 7098 21526 7100
rect 21550 7098 21606 7100
rect 21310 7046 21356 7098
rect 21356 7046 21366 7098
rect 21390 7046 21420 7098
rect 21420 7046 21432 7098
rect 21432 7046 21446 7098
rect 21470 7046 21484 7098
rect 21484 7046 21496 7098
rect 21496 7046 21526 7098
rect 21550 7046 21560 7098
rect 21560 7046 21606 7098
rect 21310 7044 21366 7046
rect 21390 7044 21446 7046
rect 21470 7044 21526 7046
rect 21550 7044 21606 7046
rect 28279 7098 28335 7100
rect 28359 7098 28415 7100
rect 28439 7098 28495 7100
rect 28519 7098 28575 7100
rect 28279 7046 28325 7098
rect 28325 7046 28335 7098
rect 28359 7046 28389 7098
rect 28389 7046 28401 7098
rect 28401 7046 28415 7098
rect 28439 7046 28453 7098
rect 28453 7046 28465 7098
rect 28465 7046 28495 7098
rect 28519 7046 28529 7098
rect 28529 7046 28575 7098
rect 28279 7044 28335 7046
rect 28359 7044 28415 7046
rect 28439 7044 28495 7046
rect 28519 7044 28575 7046
rect 3888 6554 3944 6556
rect 3968 6554 4024 6556
rect 4048 6554 4104 6556
rect 4128 6554 4184 6556
rect 3888 6502 3934 6554
rect 3934 6502 3944 6554
rect 3968 6502 3998 6554
rect 3998 6502 4010 6554
rect 4010 6502 4024 6554
rect 4048 6502 4062 6554
rect 4062 6502 4074 6554
rect 4074 6502 4104 6554
rect 4128 6502 4138 6554
rect 4138 6502 4184 6554
rect 3888 6500 3944 6502
rect 3968 6500 4024 6502
rect 4048 6500 4104 6502
rect 4128 6500 4184 6502
rect 10857 6554 10913 6556
rect 10937 6554 10993 6556
rect 11017 6554 11073 6556
rect 11097 6554 11153 6556
rect 10857 6502 10903 6554
rect 10903 6502 10913 6554
rect 10937 6502 10967 6554
rect 10967 6502 10979 6554
rect 10979 6502 10993 6554
rect 11017 6502 11031 6554
rect 11031 6502 11043 6554
rect 11043 6502 11073 6554
rect 11097 6502 11107 6554
rect 11107 6502 11153 6554
rect 10857 6500 10913 6502
rect 10937 6500 10993 6502
rect 11017 6500 11073 6502
rect 11097 6500 11153 6502
rect 17826 6554 17882 6556
rect 17906 6554 17962 6556
rect 17986 6554 18042 6556
rect 18066 6554 18122 6556
rect 17826 6502 17872 6554
rect 17872 6502 17882 6554
rect 17906 6502 17936 6554
rect 17936 6502 17948 6554
rect 17948 6502 17962 6554
rect 17986 6502 18000 6554
rect 18000 6502 18012 6554
rect 18012 6502 18042 6554
rect 18066 6502 18076 6554
rect 18076 6502 18122 6554
rect 17826 6500 17882 6502
rect 17906 6500 17962 6502
rect 17986 6500 18042 6502
rect 18066 6500 18122 6502
rect 24795 6554 24851 6556
rect 24875 6554 24931 6556
rect 24955 6554 25011 6556
rect 25035 6554 25091 6556
rect 24795 6502 24841 6554
rect 24841 6502 24851 6554
rect 24875 6502 24905 6554
rect 24905 6502 24917 6554
rect 24917 6502 24931 6554
rect 24955 6502 24969 6554
rect 24969 6502 24981 6554
rect 24981 6502 25011 6554
rect 25035 6502 25045 6554
rect 25045 6502 25091 6554
rect 24795 6500 24851 6502
rect 24875 6500 24931 6502
rect 24955 6500 25011 6502
rect 25035 6500 25091 6502
rect 7372 6010 7428 6012
rect 7452 6010 7508 6012
rect 7532 6010 7588 6012
rect 7612 6010 7668 6012
rect 7372 5958 7418 6010
rect 7418 5958 7428 6010
rect 7452 5958 7482 6010
rect 7482 5958 7494 6010
rect 7494 5958 7508 6010
rect 7532 5958 7546 6010
rect 7546 5958 7558 6010
rect 7558 5958 7588 6010
rect 7612 5958 7622 6010
rect 7622 5958 7668 6010
rect 7372 5956 7428 5958
rect 7452 5956 7508 5958
rect 7532 5956 7588 5958
rect 7612 5956 7668 5958
rect 14341 6010 14397 6012
rect 14421 6010 14477 6012
rect 14501 6010 14557 6012
rect 14581 6010 14637 6012
rect 14341 5958 14387 6010
rect 14387 5958 14397 6010
rect 14421 5958 14451 6010
rect 14451 5958 14463 6010
rect 14463 5958 14477 6010
rect 14501 5958 14515 6010
rect 14515 5958 14527 6010
rect 14527 5958 14557 6010
rect 14581 5958 14591 6010
rect 14591 5958 14637 6010
rect 14341 5956 14397 5958
rect 14421 5956 14477 5958
rect 14501 5956 14557 5958
rect 14581 5956 14637 5958
rect 21310 6010 21366 6012
rect 21390 6010 21446 6012
rect 21470 6010 21526 6012
rect 21550 6010 21606 6012
rect 21310 5958 21356 6010
rect 21356 5958 21366 6010
rect 21390 5958 21420 6010
rect 21420 5958 21432 6010
rect 21432 5958 21446 6010
rect 21470 5958 21484 6010
rect 21484 5958 21496 6010
rect 21496 5958 21526 6010
rect 21550 5958 21560 6010
rect 21560 5958 21606 6010
rect 21310 5956 21366 5958
rect 21390 5956 21446 5958
rect 21470 5956 21526 5958
rect 21550 5956 21606 5958
rect 28279 6010 28335 6012
rect 28359 6010 28415 6012
rect 28439 6010 28495 6012
rect 28519 6010 28575 6012
rect 28279 5958 28325 6010
rect 28325 5958 28335 6010
rect 28359 5958 28389 6010
rect 28389 5958 28401 6010
rect 28401 5958 28415 6010
rect 28439 5958 28453 6010
rect 28453 5958 28465 6010
rect 28465 5958 28495 6010
rect 28519 5958 28529 6010
rect 28529 5958 28575 6010
rect 28279 5956 28335 5958
rect 28359 5956 28415 5958
rect 28439 5956 28495 5958
rect 28519 5956 28575 5958
rect 3888 5466 3944 5468
rect 3968 5466 4024 5468
rect 4048 5466 4104 5468
rect 4128 5466 4184 5468
rect 3888 5414 3934 5466
rect 3934 5414 3944 5466
rect 3968 5414 3998 5466
rect 3998 5414 4010 5466
rect 4010 5414 4024 5466
rect 4048 5414 4062 5466
rect 4062 5414 4074 5466
rect 4074 5414 4104 5466
rect 4128 5414 4138 5466
rect 4138 5414 4184 5466
rect 3888 5412 3944 5414
rect 3968 5412 4024 5414
rect 4048 5412 4104 5414
rect 4128 5412 4184 5414
rect 10857 5466 10913 5468
rect 10937 5466 10993 5468
rect 11017 5466 11073 5468
rect 11097 5466 11153 5468
rect 10857 5414 10903 5466
rect 10903 5414 10913 5466
rect 10937 5414 10967 5466
rect 10967 5414 10979 5466
rect 10979 5414 10993 5466
rect 11017 5414 11031 5466
rect 11031 5414 11043 5466
rect 11043 5414 11073 5466
rect 11097 5414 11107 5466
rect 11107 5414 11153 5466
rect 10857 5412 10913 5414
rect 10937 5412 10993 5414
rect 11017 5412 11073 5414
rect 11097 5412 11153 5414
rect 17826 5466 17882 5468
rect 17906 5466 17962 5468
rect 17986 5466 18042 5468
rect 18066 5466 18122 5468
rect 17826 5414 17872 5466
rect 17872 5414 17882 5466
rect 17906 5414 17936 5466
rect 17936 5414 17948 5466
rect 17948 5414 17962 5466
rect 17986 5414 18000 5466
rect 18000 5414 18012 5466
rect 18012 5414 18042 5466
rect 18066 5414 18076 5466
rect 18076 5414 18122 5466
rect 17826 5412 17882 5414
rect 17906 5412 17962 5414
rect 17986 5412 18042 5414
rect 18066 5412 18122 5414
rect 24795 5466 24851 5468
rect 24875 5466 24931 5468
rect 24955 5466 25011 5468
rect 25035 5466 25091 5468
rect 24795 5414 24841 5466
rect 24841 5414 24851 5466
rect 24875 5414 24905 5466
rect 24905 5414 24917 5466
rect 24917 5414 24931 5466
rect 24955 5414 24969 5466
rect 24969 5414 24981 5466
rect 24981 5414 25011 5466
rect 25035 5414 25045 5466
rect 25045 5414 25091 5466
rect 24795 5412 24851 5414
rect 24875 5412 24931 5414
rect 24955 5412 25011 5414
rect 25035 5412 25091 5414
rect 7372 4922 7428 4924
rect 7452 4922 7508 4924
rect 7532 4922 7588 4924
rect 7612 4922 7668 4924
rect 7372 4870 7418 4922
rect 7418 4870 7428 4922
rect 7452 4870 7482 4922
rect 7482 4870 7494 4922
rect 7494 4870 7508 4922
rect 7532 4870 7546 4922
rect 7546 4870 7558 4922
rect 7558 4870 7588 4922
rect 7612 4870 7622 4922
rect 7622 4870 7668 4922
rect 7372 4868 7428 4870
rect 7452 4868 7508 4870
rect 7532 4868 7588 4870
rect 7612 4868 7668 4870
rect 14341 4922 14397 4924
rect 14421 4922 14477 4924
rect 14501 4922 14557 4924
rect 14581 4922 14637 4924
rect 14341 4870 14387 4922
rect 14387 4870 14397 4922
rect 14421 4870 14451 4922
rect 14451 4870 14463 4922
rect 14463 4870 14477 4922
rect 14501 4870 14515 4922
rect 14515 4870 14527 4922
rect 14527 4870 14557 4922
rect 14581 4870 14591 4922
rect 14591 4870 14637 4922
rect 14341 4868 14397 4870
rect 14421 4868 14477 4870
rect 14501 4868 14557 4870
rect 14581 4868 14637 4870
rect 21310 4922 21366 4924
rect 21390 4922 21446 4924
rect 21470 4922 21526 4924
rect 21550 4922 21606 4924
rect 21310 4870 21356 4922
rect 21356 4870 21366 4922
rect 21390 4870 21420 4922
rect 21420 4870 21432 4922
rect 21432 4870 21446 4922
rect 21470 4870 21484 4922
rect 21484 4870 21496 4922
rect 21496 4870 21526 4922
rect 21550 4870 21560 4922
rect 21560 4870 21606 4922
rect 21310 4868 21366 4870
rect 21390 4868 21446 4870
rect 21470 4868 21526 4870
rect 21550 4868 21606 4870
rect 28279 4922 28335 4924
rect 28359 4922 28415 4924
rect 28439 4922 28495 4924
rect 28519 4922 28575 4924
rect 28279 4870 28325 4922
rect 28325 4870 28335 4922
rect 28359 4870 28389 4922
rect 28389 4870 28401 4922
rect 28401 4870 28415 4922
rect 28439 4870 28453 4922
rect 28453 4870 28465 4922
rect 28465 4870 28495 4922
rect 28519 4870 28529 4922
rect 28529 4870 28575 4922
rect 28279 4868 28335 4870
rect 28359 4868 28415 4870
rect 28439 4868 28495 4870
rect 28519 4868 28575 4870
rect 3888 4378 3944 4380
rect 3968 4378 4024 4380
rect 4048 4378 4104 4380
rect 4128 4378 4184 4380
rect 3888 4326 3934 4378
rect 3934 4326 3944 4378
rect 3968 4326 3998 4378
rect 3998 4326 4010 4378
rect 4010 4326 4024 4378
rect 4048 4326 4062 4378
rect 4062 4326 4074 4378
rect 4074 4326 4104 4378
rect 4128 4326 4138 4378
rect 4138 4326 4184 4378
rect 3888 4324 3944 4326
rect 3968 4324 4024 4326
rect 4048 4324 4104 4326
rect 4128 4324 4184 4326
rect 10857 4378 10913 4380
rect 10937 4378 10993 4380
rect 11017 4378 11073 4380
rect 11097 4378 11153 4380
rect 10857 4326 10903 4378
rect 10903 4326 10913 4378
rect 10937 4326 10967 4378
rect 10967 4326 10979 4378
rect 10979 4326 10993 4378
rect 11017 4326 11031 4378
rect 11031 4326 11043 4378
rect 11043 4326 11073 4378
rect 11097 4326 11107 4378
rect 11107 4326 11153 4378
rect 10857 4324 10913 4326
rect 10937 4324 10993 4326
rect 11017 4324 11073 4326
rect 11097 4324 11153 4326
rect 17826 4378 17882 4380
rect 17906 4378 17962 4380
rect 17986 4378 18042 4380
rect 18066 4378 18122 4380
rect 17826 4326 17872 4378
rect 17872 4326 17882 4378
rect 17906 4326 17936 4378
rect 17936 4326 17948 4378
rect 17948 4326 17962 4378
rect 17986 4326 18000 4378
rect 18000 4326 18012 4378
rect 18012 4326 18042 4378
rect 18066 4326 18076 4378
rect 18076 4326 18122 4378
rect 17826 4324 17882 4326
rect 17906 4324 17962 4326
rect 17986 4324 18042 4326
rect 18066 4324 18122 4326
rect 24795 4378 24851 4380
rect 24875 4378 24931 4380
rect 24955 4378 25011 4380
rect 25035 4378 25091 4380
rect 24795 4326 24841 4378
rect 24841 4326 24851 4378
rect 24875 4326 24905 4378
rect 24905 4326 24917 4378
rect 24917 4326 24931 4378
rect 24955 4326 24969 4378
rect 24969 4326 24981 4378
rect 24981 4326 25011 4378
rect 25035 4326 25045 4378
rect 25045 4326 25091 4378
rect 24795 4324 24851 4326
rect 24875 4324 24931 4326
rect 24955 4324 25011 4326
rect 25035 4324 25091 4326
rect 7372 3834 7428 3836
rect 7452 3834 7508 3836
rect 7532 3834 7588 3836
rect 7612 3834 7668 3836
rect 7372 3782 7418 3834
rect 7418 3782 7428 3834
rect 7452 3782 7482 3834
rect 7482 3782 7494 3834
rect 7494 3782 7508 3834
rect 7532 3782 7546 3834
rect 7546 3782 7558 3834
rect 7558 3782 7588 3834
rect 7612 3782 7622 3834
rect 7622 3782 7668 3834
rect 7372 3780 7428 3782
rect 7452 3780 7508 3782
rect 7532 3780 7588 3782
rect 7612 3780 7668 3782
rect 14341 3834 14397 3836
rect 14421 3834 14477 3836
rect 14501 3834 14557 3836
rect 14581 3834 14637 3836
rect 14341 3782 14387 3834
rect 14387 3782 14397 3834
rect 14421 3782 14451 3834
rect 14451 3782 14463 3834
rect 14463 3782 14477 3834
rect 14501 3782 14515 3834
rect 14515 3782 14527 3834
rect 14527 3782 14557 3834
rect 14581 3782 14591 3834
rect 14591 3782 14637 3834
rect 14341 3780 14397 3782
rect 14421 3780 14477 3782
rect 14501 3780 14557 3782
rect 14581 3780 14637 3782
rect 21310 3834 21366 3836
rect 21390 3834 21446 3836
rect 21470 3834 21526 3836
rect 21550 3834 21606 3836
rect 21310 3782 21356 3834
rect 21356 3782 21366 3834
rect 21390 3782 21420 3834
rect 21420 3782 21432 3834
rect 21432 3782 21446 3834
rect 21470 3782 21484 3834
rect 21484 3782 21496 3834
rect 21496 3782 21526 3834
rect 21550 3782 21560 3834
rect 21560 3782 21606 3834
rect 21310 3780 21366 3782
rect 21390 3780 21446 3782
rect 21470 3780 21526 3782
rect 21550 3780 21606 3782
rect 28279 3834 28335 3836
rect 28359 3834 28415 3836
rect 28439 3834 28495 3836
rect 28519 3834 28575 3836
rect 28279 3782 28325 3834
rect 28325 3782 28335 3834
rect 28359 3782 28389 3834
rect 28389 3782 28401 3834
rect 28401 3782 28415 3834
rect 28439 3782 28453 3834
rect 28453 3782 28465 3834
rect 28465 3782 28495 3834
rect 28519 3782 28529 3834
rect 28529 3782 28575 3834
rect 28279 3780 28335 3782
rect 28359 3780 28415 3782
rect 28439 3780 28495 3782
rect 28519 3780 28575 3782
rect 3888 3290 3944 3292
rect 3968 3290 4024 3292
rect 4048 3290 4104 3292
rect 4128 3290 4184 3292
rect 3888 3238 3934 3290
rect 3934 3238 3944 3290
rect 3968 3238 3998 3290
rect 3998 3238 4010 3290
rect 4010 3238 4024 3290
rect 4048 3238 4062 3290
rect 4062 3238 4074 3290
rect 4074 3238 4104 3290
rect 4128 3238 4138 3290
rect 4138 3238 4184 3290
rect 3888 3236 3944 3238
rect 3968 3236 4024 3238
rect 4048 3236 4104 3238
rect 4128 3236 4184 3238
rect 10857 3290 10913 3292
rect 10937 3290 10993 3292
rect 11017 3290 11073 3292
rect 11097 3290 11153 3292
rect 10857 3238 10903 3290
rect 10903 3238 10913 3290
rect 10937 3238 10967 3290
rect 10967 3238 10979 3290
rect 10979 3238 10993 3290
rect 11017 3238 11031 3290
rect 11031 3238 11043 3290
rect 11043 3238 11073 3290
rect 11097 3238 11107 3290
rect 11107 3238 11153 3290
rect 10857 3236 10913 3238
rect 10937 3236 10993 3238
rect 11017 3236 11073 3238
rect 11097 3236 11153 3238
rect 17826 3290 17882 3292
rect 17906 3290 17962 3292
rect 17986 3290 18042 3292
rect 18066 3290 18122 3292
rect 17826 3238 17872 3290
rect 17872 3238 17882 3290
rect 17906 3238 17936 3290
rect 17936 3238 17948 3290
rect 17948 3238 17962 3290
rect 17986 3238 18000 3290
rect 18000 3238 18012 3290
rect 18012 3238 18042 3290
rect 18066 3238 18076 3290
rect 18076 3238 18122 3290
rect 17826 3236 17882 3238
rect 17906 3236 17962 3238
rect 17986 3236 18042 3238
rect 18066 3236 18122 3238
rect 24795 3290 24851 3292
rect 24875 3290 24931 3292
rect 24955 3290 25011 3292
rect 25035 3290 25091 3292
rect 24795 3238 24841 3290
rect 24841 3238 24851 3290
rect 24875 3238 24905 3290
rect 24905 3238 24917 3290
rect 24917 3238 24931 3290
rect 24955 3238 24969 3290
rect 24969 3238 24981 3290
rect 24981 3238 25011 3290
rect 25035 3238 25045 3290
rect 25045 3238 25091 3290
rect 24795 3236 24851 3238
rect 24875 3236 24931 3238
rect 24955 3236 25011 3238
rect 25035 3236 25091 3238
rect 7372 2746 7428 2748
rect 7452 2746 7508 2748
rect 7532 2746 7588 2748
rect 7612 2746 7668 2748
rect 7372 2694 7418 2746
rect 7418 2694 7428 2746
rect 7452 2694 7482 2746
rect 7482 2694 7494 2746
rect 7494 2694 7508 2746
rect 7532 2694 7546 2746
rect 7546 2694 7558 2746
rect 7558 2694 7588 2746
rect 7612 2694 7622 2746
rect 7622 2694 7668 2746
rect 7372 2692 7428 2694
rect 7452 2692 7508 2694
rect 7532 2692 7588 2694
rect 7612 2692 7668 2694
rect 14341 2746 14397 2748
rect 14421 2746 14477 2748
rect 14501 2746 14557 2748
rect 14581 2746 14637 2748
rect 14341 2694 14387 2746
rect 14387 2694 14397 2746
rect 14421 2694 14451 2746
rect 14451 2694 14463 2746
rect 14463 2694 14477 2746
rect 14501 2694 14515 2746
rect 14515 2694 14527 2746
rect 14527 2694 14557 2746
rect 14581 2694 14591 2746
rect 14591 2694 14637 2746
rect 14341 2692 14397 2694
rect 14421 2692 14477 2694
rect 14501 2692 14557 2694
rect 14581 2692 14637 2694
rect 21310 2746 21366 2748
rect 21390 2746 21446 2748
rect 21470 2746 21526 2748
rect 21550 2746 21606 2748
rect 21310 2694 21356 2746
rect 21356 2694 21366 2746
rect 21390 2694 21420 2746
rect 21420 2694 21432 2746
rect 21432 2694 21446 2746
rect 21470 2694 21484 2746
rect 21484 2694 21496 2746
rect 21496 2694 21526 2746
rect 21550 2694 21560 2746
rect 21560 2694 21606 2746
rect 21310 2692 21366 2694
rect 21390 2692 21446 2694
rect 21470 2692 21526 2694
rect 21550 2692 21606 2694
rect 28279 2746 28335 2748
rect 28359 2746 28415 2748
rect 28439 2746 28495 2748
rect 28519 2746 28575 2748
rect 28279 2694 28325 2746
rect 28325 2694 28335 2746
rect 28359 2694 28389 2746
rect 28389 2694 28401 2746
rect 28401 2694 28415 2746
rect 28439 2694 28453 2746
rect 28453 2694 28465 2746
rect 28465 2694 28495 2746
rect 28519 2694 28529 2746
rect 28529 2694 28575 2746
rect 28279 2692 28335 2694
rect 28359 2692 28415 2694
rect 28439 2692 28495 2694
rect 28519 2692 28575 2694
rect 3888 2202 3944 2204
rect 3968 2202 4024 2204
rect 4048 2202 4104 2204
rect 4128 2202 4184 2204
rect 3888 2150 3934 2202
rect 3934 2150 3944 2202
rect 3968 2150 3998 2202
rect 3998 2150 4010 2202
rect 4010 2150 4024 2202
rect 4048 2150 4062 2202
rect 4062 2150 4074 2202
rect 4074 2150 4104 2202
rect 4128 2150 4138 2202
rect 4138 2150 4184 2202
rect 3888 2148 3944 2150
rect 3968 2148 4024 2150
rect 4048 2148 4104 2150
rect 4128 2148 4184 2150
rect 10857 2202 10913 2204
rect 10937 2202 10993 2204
rect 11017 2202 11073 2204
rect 11097 2202 11153 2204
rect 10857 2150 10903 2202
rect 10903 2150 10913 2202
rect 10937 2150 10967 2202
rect 10967 2150 10979 2202
rect 10979 2150 10993 2202
rect 11017 2150 11031 2202
rect 11031 2150 11043 2202
rect 11043 2150 11073 2202
rect 11097 2150 11107 2202
rect 11107 2150 11153 2202
rect 10857 2148 10913 2150
rect 10937 2148 10993 2150
rect 11017 2148 11073 2150
rect 11097 2148 11153 2150
rect 17826 2202 17882 2204
rect 17906 2202 17962 2204
rect 17986 2202 18042 2204
rect 18066 2202 18122 2204
rect 17826 2150 17872 2202
rect 17872 2150 17882 2202
rect 17906 2150 17936 2202
rect 17936 2150 17948 2202
rect 17948 2150 17962 2202
rect 17986 2150 18000 2202
rect 18000 2150 18012 2202
rect 18012 2150 18042 2202
rect 18066 2150 18076 2202
rect 18076 2150 18122 2202
rect 17826 2148 17882 2150
rect 17906 2148 17962 2150
rect 17986 2148 18042 2150
rect 18066 2148 18122 2150
rect 24795 2202 24851 2204
rect 24875 2202 24931 2204
rect 24955 2202 25011 2204
rect 25035 2202 25091 2204
rect 24795 2150 24841 2202
rect 24841 2150 24851 2202
rect 24875 2150 24905 2202
rect 24905 2150 24917 2202
rect 24917 2150 24931 2202
rect 24955 2150 24969 2202
rect 24969 2150 24981 2202
rect 24981 2150 25011 2202
rect 25035 2150 25045 2202
rect 25045 2150 25091 2202
rect 24795 2148 24851 2150
rect 24875 2148 24931 2150
rect 24955 2148 25011 2150
rect 25035 2148 25091 2150
rect 7372 1658 7428 1660
rect 7452 1658 7508 1660
rect 7532 1658 7588 1660
rect 7612 1658 7668 1660
rect 7372 1606 7418 1658
rect 7418 1606 7428 1658
rect 7452 1606 7482 1658
rect 7482 1606 7494 1658
rect 7494 1606 7508 1658
rect 7532 1606 7546 1658
rect 7546 1606 7558 1658
rect 7558 1606 7588 1658
rect 7612 1606 7622 1658
rect 7622 1606 7668 1658
rect 7372 1604 7428 1606
rect 7452 1604 7508 1606
rect 7532 1604 7588 1606
rect 7612 1604 7668 1606
rect 14341 1658 14397 1660
rect 14421 1658 14477 1660
rect 14501 1658 14557 1660
rect 14581 1658 14637 1660
rect 14341 1606 14387 1658
rect 14387 1606 14397 1658
rect 14421 1606 14451 1658
rect 14451 1606 14463 1658
rect 14463 1606 14477 1658
rect 14501 1606 14515 1658
rect 14515 1606 14527 1658
rect 14527 1606 14557 1658
rect 14581 1606 14591 1658
rect 14591 1606 14637 1658
rect 14341 1604 14397 1606
rect 14421 1604 14477 1606
rect 14501 1604 14557 1606
rect 14581 1604 14637 1606
rect 21310 1658 21366 1660
rect 21390 1658 21446 1660
rect 21470 1658 21526 1660
rect 21550 1658 21606 1660
rect 21310 1606 21356 1658
rect 21356 1606 21366 1658
rect 21390 1606 21420 1658
rect 21420 1606 21432 1658
rect 21432 1606 21446 1658
rect 21470 1606 21484 1658
rect 21484 1606 21496 1658
rect 21496 1606 21526 1658
rect 21550 1606 21560 1658
rect 21560 1606 21606 1658
rect 21310 1604 21366 1606
rect 21390 1604 21446 1606
rect 21470 1604 21526 1606
rect 21550 1604 21606 1606
rect 28279 1658 28335 1660
rect 28359 1658 28415 1660
rect 28439 1658 28495 1660
rect 28519 1658 28575 1660
rect 28279 1606 28325 1658
rect 28325 1606 28335 1658
rect 28359 1606 28389 1658
rect 28389 1606 28401 1658
rect 28401 1606 28415 1658
rect 28439 1606 28453 1658
rect 28453 1606 28465 1658
rect 28465 1606 28495 1658
rect 28519 1606 28529 1658
rect 28529 1606 28575 1658
rect 28279 1604 28335 1606
rect 28359 1604 28415 1606
rect 28439 1604 28495 1606
rect 28519 1604 28575 1606
rect 3888 1114 3944 1116
rect 3968 1114 4024 1116
rect 4048 1114 4104 1116
rect 4128 1114 4184 1116
rect 3888 1062 3934 1114
rect 3934 1062 3944 1114
rect 3968 1062 3998 1114
rect 3998 1062 4010 1114
rect 4010 1062 4024 1114
rect 4048 1062 4062 1114
rect 4062 1062 4074 1114
rect 4074 1062 4104 1114
rect 4128 1062 4138 1114
rect 4138 1062 4184 1114
rect 3888 1060 3944 1062
rect 3968 1060 4024 1062
rect 4048 1060 4104 1062
rect 4128 1060 4184 1062
rect 10857 1114 10913 1116
rect 10937 1114 10993 1116
rect 11017 1114 11073 1116
rect 11097 1114 11153 1116
rect 10857 1062 10903 1114
rect 10903 1062 10913 1114
rect 10937 1062 10967 1114
rect 10967 1062 10979 1114
rect 10979 1062 10993 1114
rect 11017 1062 11031 1114
rect 11031 1062 11043 1114
rect 11043 1062 11073 1114
rect 11097 1062 11107 1114
rect 11107 1062 11153 1114
rect 10857 1060 10913 1062
rect 10937 1060 10993 1062
rect 11017 1060 11073 1062
rect 11097 1060 11153 1062
rect 17826 1114 17882 1116
rect 17906 1114 17962 1116
rect 17986 1114 18042 1116
rect 18066 1114 18122 1116
rect 17826 1062 17872 1114
rect 17872 1062 17882 1114
rect 17906 1062 17936 1114
rect 17936 1062 17948 1114
rect 17948 1062 17962 1114
rect 17986 1062 18000 1114
rect 18000 1062 18012 1114
rect 18012 1062 18042 1114
rect 18066 1062 18076 1114
rect 18076 1062 18122 1114
rect 17826 1060 17882 1062
rect 17906 1060 17962 1062
rect 17986 1060 18042 1062
rect 18066 1060 18122 1062
rect 24795 1114 24851 1116
rect 24875 1114 24931 1116
rect 24955 1114 25011 1116
rect 25035 1114 25091 1116
rect 24795 1062 24841 1114
rect 24841 1062 24851 1114
rect 24875 1062 24905 1114
rect 24905 1062 24917 1114
rect 24917 1062 24931 1114
rect 24955 1062 24969 1114
rect 24969 1062 24981 1114
rect 24981 1062 25011 1114
rect 25035 1062 25045 1114
rect 25045 1062 25091 1114
rect 24795 1060 24851 1062
rect 24875 1060 24931 1062
rect 24955 1060 25011 1062
rect 25035 1060 25091 1062
rect 7372 570 7428 572
rect 7452 570 7508 572
rect 7532 570 7588 572
rect 7612 570 7668 572
rect 7372 518 7418 570
rect 7418 518 7428 570
rect 7452 518 7482 570
rect 7482 518 7494 570
rect 7494 518 7508 570
rect 7532 518 7546 570
rect 7546 518 7558 570
rect 7558 518 7588 570
rect 7612 518 7622 570
rect 7622 518 7668 570
rect 7372 516 7428 518
rect 7452 516 7508 518
rect 7532 516 7588 518
rect 7612 516 7668 518
rect 14341 570 14397 572
rect 14421 570 14477 572
rect 14501 570 14557 572
rect 14581 570 14637 572
rect 14341 518 14387 570
rect 14387 518 14397 570
rect 14421 518 14451 570
rect 14451 518 14463 570
rect 14463 518 14477 570
rect 14501 518 14515 570
rect 14515 518 14527 570
rect 14527 518 14557 570
rect 14581 518 14591 570
rect 14591 518 14637 570
rect 14341 516 14397 518
rect 14421 516 14477 518
rect 14501 516 14557 518
rect 14581 516 14637 518
rect 21310 570 21366 572
rect 21390 570 21446 572
rect 21470 570 21526 572
rect 21550 570 21606 572
rect 21310 518 21356 570
rect 21356 518 21366 570
rect 21390 518 21420 570
rect 21420 518 21432 570
rect 21432 518 21446 570
rect 21470 518 21484 570
rect 21484 518 21496 570
rect 21496 518 21526 570
rect 21550 518 21560 570
rect 21560 518 21606 570
rect 21310 516 21366 518
rect 21390 516 21446 518
rect 21470 516 21526 518
rect 21550 516 21606 518
rect 28279 570 28335 572
rect 28359 570 28415 572
rect 28439 570 28495 572
rect 28519 570 28575 572
rect 28279 518 28325 570
rect 28325 518 28335 570
rect 28359 518 28389 570
rect 28389 518 28401 570
rect 28401 518 28415 570
rect 28439 518 28453 570
rect 28453 518 28465 570
rect 28465 518 28495 570
rect 28519 518 28529 570
rect 28529 518 28575 570
rect 28279 516 28335 518
rect 28359 516 28415 518
rect 28439 516 28495 518
rect 28519 516 28575 518
<< metal3 >>
rect 3878 28320 4194 28321
rect 3878 28256 3884 28320
rect 3948 28256 3964 28320
rect 4028 28256 4044 28320
rect 4108 28256 4124 28320
rect 4188 28256 4194 28320
rect 3878 28255 4194 28256
rect 10847 28320 11163 28321
rect 10847 28256 10853 28320
rect 10917 28256 10933 28320
rect 10997 28256 11013 28320
rect 11077 28256 11093 28320
rect 11157 28256 11163 28320
rect 10847 28255 11163 28256
rect 17816 28320 18132 28321
rect 17816 28256 17822 28320
rect 17886 28256 17902 28320
rect 17966 28256 17982 28320
rect 18046 28256 18062 28320
rect 18126 28256 18132 28320
rect 17816 28255 18132 28256
rect 24785 28320 25101 28321
rect 24785 28256 24791 28320
rect 24855 28256 24871 28320
rect 24935 28256 24951 28320
rect 25015 28256 25031 28320
rect 25095 28256 25101 28320
rect 24785 28255 25101 28256
rect 7362 27776 7678 27777
rect 7362 27712 7368 27776
rect 7432 27712 7448 27776
rect 7512 27712 7528 27776
rect 7592 27712 7608 27776
rect 7672 27712 7678 27776
rect 7362 27711 7678 27712
rect 14331 27776 14647 27777
rect 14331 27712 14337 27776
rect 14401 27712 14417 27776
rect 14481 27712 14497 27776
rect 14561 27712 14577 27776
rect 14641 27712 14647 27776
rect 14331 27711 14647 27712
rect 21300 27776 21616 27777
rect 21300 27712 21306 27776
rect 21370 27712 21386 27776
rect 21450 27712 21466 27776
rect 21530 27712 21546 27776
rect 21610 27712 21616 27776
rect 21300 27711 21616 27712
rect 28269 27776 28585 27777
rect 28269 27712 28275 27776
rect 28339 27712 28355 27776
rect 28419 27712 28435 27776
rect 28499 27712 28515 27776
rect 28579 27712 28585 27776
rect 28269 27711 28585 27712
rect 3878 27232 4194 27233
rect 3878 27168 3884 27232
rect 3948 27168 3964 27232
rect 4028 27168 4044 27232
rect 4108 27168 4124 27232
rect 4188 27168 4194 27232
rect 3878 27167 4194 27168
rect 10847 27232 11163 27233
rect 10847 27168 10853 27232
rect 10917 27168 10933 27232
rect 10997 27168 11013 27232
rect 11077 27168 11093 27232
rect 11157 27168 11163 27232
rect 10847 27167 11163 27168
rect 17816 27232 18132 27233
rect 17816 27168 17822 27232
rect 17886 27168 17902 27232
rect 17966 27168 17982 27232
rect 18046 27168 18062 27232
rect 18126 27168 18132 27232
rect 17816 27167 18132 27168
rect 24785 27232 25101 27233
rect 24785 27168 24791 27232
rect 24855 27168 24871 27232
rect 24935 27168 24951 27232
rect 25015 27168 25031 27232
rect 25095 27168 25101 27232
rect 24785 27167 25101 27168
rect 7362 26688 7678 26689
rect 7362 26624 7368 26688
rect 7432 26624 7448 26688
rect 7512 26624 7528 26688
rect 7592 26624 7608 26688
rect 7672 26624 7678 26688
rect 7362 26623 7678 26624
rect 14331 26688 14647 26689
rect 14331 26624 14337 26688
rect 14401 26624 14417 26688
rect 14481 26624 14497 26688
rect 14561 26624 14577 26688
rect 14641 26624 14647 26688
rect 14331 26623 14647 26624
rect 21300 26688 21616 26689
rect 21300 26624 21306 26688
rect 21370 26624 21386 26688
rect 21450 26624 21466 26688
rect 21530 26624 21546 26688
rect 21610 26624 21616 26688
rect 21300 26623 21616 26624
rect 28269 26688 28585 26689
rect 28269 26624 28275 26688
rect 28339 26624 28355 26688
rect 28419 26624 28435 26688
rect 28499 26624 28515 26688
rect 28579 26624 28585 26688
rect 28269 26623 28585 26624
rect 3878 26144 4194 26145
rect 3878 26080 3884 26144
rect 3948 26080 3964 26144
rect 4028 26080 4044 26144
rect 4108 26080 4124 26144
rect 4188 26080 4194 26144
rect 3878 26079 4194 26080
rect 10847 26144 11163 26145
rect 10847 26080 10853 26144
rect 10917 26080 10933 26144
rect 10997 26080 11013 26144
rect 11077 26080 11093 26144
rect 11157 26080 11163 26144
rect 10847 26079 11163 26080
rect 17816 26144 18132 26145
rect 17816 26080 17822 26144
rect 17886 26080 17902 26144
rect 17966 26080 17982 26144
rect 18046 26080 18062 26144
rect 18126 26080 18132 26144
rect 17816 26079 18132 26080
rect 24785 26144 25101 26145
rect 24785 26080 24791 26144
rect 24855 26080 24871 26144
rect 24935 26080 24951 26144
rect 25015 26080 25031 26144
rect 25095 26080 25101 26144
rect 24785 26079 25101 26080
rect 7362 25600 7678 25601
rect 7362 25536 7368 25600
rect 7432 25536 7448 25600
rect 7512 25536 7528 25600
rect 7592 25536 7608 25600
rect 7672 25536 7678 25600
rect 7362 25535 7678 25536
rect 14331 25600 14647 25601
rect 14331 25536 14337 25600
rect 14401 25536 14417 25600
rect 14481 25536 14497 25600
rect 14561 25536 14577 25600
rect 14641 25536 14647 25600
rect 14331 25535 14647 25536
rect 21300 25600 21616 25601
rect 21300 25536 21306 25600
rect 21370 25536 21386 25600
rect 21450 25536 21466 25600
rect 21530 25536 21546 25600
rect 21610 25536 21616 25600
rect 21300 25535 21616 25536
rect 28269 25600 28585 25601
rect 28269 25536 28275 25600
rect 28339 25536 28355 25600
rect 28419 25536 28435 25600
rect 28499 25536 28515 25600
rect 28579 25536 28585 25600
rect 28269 25535 28585 25536
rect 13721 25394 13787 25397
rect 18597 25394 18663 25397
rect 13721 25392 18663 25394
rect 13721 25336 13726 25392
rect 13782 25336 18602 25392
rect 18658 25336 18663 25392
rect 13721 25334 18663 25336
rect 13721 25331 13787 25334
rect 18597 25331 18663 25334
rect 3878 25056 4194 25057
rect 3878 24992 3884 25056
rect 3948 24992 3964 25056
rect 4028 24992 4044 25056
rect 4108 24992 4124 25056
rect 4188 24992 4194 25056
rect 3878 24991 4194 24992
rect 10847 25056 11163 25057
rect 10847 24992 10853 25056
rect 10917 24992 10933 25056
rect 10997 24992 11013 25056
rect 11077 24992 11093 25056
rect 11157 24992 11163 25056
rect 10847 24991 11163 24992
rect 17816 25056 18132 25057
rect 17816 24992 17822 25056
rect 17886 24992 17902 25056
rect 17966 24992 17982 25056
rect 18046 24992 18062 25056
rect 18126 24992 18132 25056
rect 17816 24991 18132 24992
rect 24785 25056 25101 25057
rect 24785 24992 24791 25056
rect 24855 24992 24871 25056
rect 24935 24992 24951 25056
rect 25015 24992 25031 25056
rect 25095 24992 25101 25056
rect 24785 24991 25101 24992
rect 7362 24512 7678 24513
rect 7362 24448 7368 24512
rect 7432 24448 7448 24512
rect 7512 24448 7528 24512
rect 7592 24448 7608 24512
rect 7672 24448 7678 24512
rect 7362 24447 7678 24448
rect 14331 24512 14647 24513
rect 14331 24448 14337 24512
rect 14401 24448 14417 24512
rect 14481 24448 14497 24512
rect 14561 24448 14577 24512
rect 14641 24448 14647 24512
rect 14331 24447 14647 24448
rect 21300 24512 21616 24513
rect 21300 24448 21306 24512
rect 21370 24448 21386 24512
rect 21450 24448 21466 24512
rect 21530 24448 21546 24512
rect 21610 24448 21616 24512
rect 21300 24447 21616 24448
rect 28269 24512 28585 24513
rect 28269 24448 28275 24512
rect 28339 24448 28355 24512
rect 28419 24448 28435 24512
rect 28499 24448 28515 24512
rect 28579 24448 28585 24512
rect 28269 24447 28585 24448
rect 3878 23968 4194 23969
rect 3878 23904 3884 23968
rect 3948 23904 3964 23968
rect 4028 23904 4044 23968
rect 4108 23904 4124 23968
rect 4188 23904 4194 23968
rect 3878 23903 4194 23904
rect 10847 23968 11163 23969
rect 10847 23904 10853 23968
rect 10917 23904 10933 23968
rect 10997 23904 11013 23968
rect 11077 23904 11093 23968
rect 11157 23904 11163 23968
rect 10847 23903 11163 23904
rect 17816 23968 18132 23969
rect 17816 23904 17822 23968
rect 17886 23904 17902 23968
rect 17966 23904 17982 23968
rect 18046 23904 18062 23968
rect 18126 23904 18132 23968
rect 17816 23903 18132 23904
rect 24785 23968 25101 23969
rect 24785 23904 24791 23968
rect 24855 23904 24871 23968
rect 24935 23904 24951 23968
rect 25015 23904 25031 23968
rect 25095 23904 25101 23968
rect 24785 23903 25101 23904
rect 7362 23424 7678 23425
rect 7362 23360 7368 23424
rect 7432 23360 7448 23424
rect 7512 23360 7528 23424
rect 7592 23360 7608 23424
rect 7672 23360 7678 23424
rect 7362 23359 7678 23360
rect 14331 23424 14647 23425
rect 14331 23360 14337 23424
rect 14401 23360 14417 23424
rect 14481 23360 14497 23424
rect 14561 23360 14577 23424
rect 14641 23360 14647 23424
rect 14331 23359 14647 23360
rect 21300 23424 21616 23425
rect 21300 23360 21306 23424
rect 21370 23360 21386 23424
rect 21450 23360 21466 23424
rect 21530 23360 21546 23424
rect 21610 23360 21616 23424
rect 21300 23359 21616 23360
rect 28269 23424 28585 23425
rect 28269 23360 28275 23424
rect 28339 23360 28355 23424
rect 28419 23360 28435 23424
rect 28499 23360 28515 23424
rect 28579 23360 28585 23424
rect 28269 23359 28585 23360
rect 15009 23218 15075 23221
rect 22921 23218 22987 23221
rect 15009 23216 22987 23218
rect 15009 23160 15014 23216
rect 15070 23160 22926 23216
rect 22982 23160 22987 23216
rect 15009 23158 22987 23160
rect 15009 23155 15075 23158
rect 22921 23155 22987 23158
rect 2221 23082 2287 23085
rect 13169 23082 13235 23085
rect 2221 23080 13235 23082
rect 2221 23024 2226 23080
rect 2282 23024 13174 23080
rect 13230 23024 13235 23080
rect 2221 23022 13235 23024
rect 2221 23019 2287 23022
rect 13169 23019 13235 23022
rect 13721 23082 13787 23085
rect 17309 23082 17375 23085
rect 18781 23082 18847 23085
rect 13721 23080 17375 23082
rect 13721 23024 13726 23080
rect 13782 23024 17314 23080
rect 17370 23024 17375 23080
rect 13721 23022 17375 23024
rect 13721 23019 13787 23022
rect 17309 23019 17375 23022
rect 17542 23080 18847 23082
rect 17542 23024 18786 23080
rect 18842 23024 18847 23080
rect 17542 23022 18847 23024
rect 12341 22946 12407 22949
rect 15837 22946 15903 22949
rect 17542 22946 17602 23022
rect 18781 23019 18847 23022
rect 12341 22944 17602 22946
rect 12341 22888 12346 22944
rect 12402 22888 15842 22944
rect 15898 22888 17602 22944
rect 12341 22886 17602 22888
rect 12341 22883 12407 22886
rect 15837 22883 15903 22886
rect 3878 22880 4194 22881
rect 3878 22816 3884 22880
rect 3948 22816 3964 22880
rect 4028 22816 4044 22880
rect 4108 22816 4124 22880
rect 4188 22816 4194 22880
rect 3878 22815 4194 22816
rect 10847 22880 11163 22881
rect 10847 22816 10853 22880
rect 10917 22816 10933 22880
rect 10997 22816 11013 22880
rect 11077 22816 11093 22880
rect 11157 22816 11163 22880
rect 10847 22815 11163 22816
rect 17816 22880 18132 22881
rect 17816 22816 17822 22880
rect 17886 22816 17902 22880
rect 17966 22816 17982 22880
rect 18046 22816 18062 22880
rect 18126 22816 18132 22880
rect 17816 22815 18132 22816
rect 24785 22880 25101 22881
rect 24785 22816 24791 22880
rect 24855 22816 24871 22880
rect 24935 22816 24951 22880
rect 25015 22816 25031 22880
rect 25095 22816 25101 22880
rect 24785 22815 25101 22816
rect 4337 22538 4403 22541
rect 5349 22538 5415 22541
rect 4337 22536 5415 22538
rect 4337 22480 4342 22536
rect 4398 22480 5354 22536
rect 5410 22480 5415 22536
rect 4337 22478 5415 22480
rect 4337 22475 4403 22478
rect 5349 22475 5415 22478
rect 7362 22336 7678 22337
rect 7362 22272 7368 22336
rect 7432 22272 7448 22336
rect 7512 22272 7528 22336
rect 7592 22272 7608 22336
rect 7672 22272 7678 22336
rect 7362 22271 7678 22272
rect 14331 22336 14647 22337
rect 14331 22272 14337 22336
rect 14401 22272 14417 22336
rect 14481 22272 14497 22336
rect 14561 22272 14577 22336
rect 14641 22272 14647 22336
rect 14331 22271 14647 22272
rect 21300 22336 21616 22337
rect 21300 22272 21306 22336
rect 21370 22272 21386 22336
rect 21450 22272 21466 22336
rect 21530 22272 21546 22336
rect 21610 22272 21616 22336
rect 21300 22271 21616 22272
rect 28269 22336 28585 22337
rect 28269 22272 28275 22336
rect 28339 22272 28355 22336
rect 28419 22272 28435 22336
rect 28499 22272 28515 22336
rect 28579 22272 28585 22336
rect 28269 22271 28585 22272
rect 21081 22130 21147 22133
rect 23473 22130 23539 22133
rect 21081 22128 23539 22130
rect 21081 22072 21086 22128
rect 21142 22072 23478 22128
rect 23534 22072 23539 22128
rect 21081 22070 23539 22072
rect 21081 22067 21147 22070
rect 23473 22067 23539 22070
rect 7741 21994 7807 21997
rect 13721 21994 13787 21997
rect 7741 21992 13787 21994
rect 7741 21936 7746 21992
rect 7802 21936 13726 21992
rect 13782 21936 13787 21992
rect 7741 21934 13787 21936
rect 7741 21931 7807 21934
rect 13721 21931 13787 21934
rect 3878 21792 4194 21793
rect 3878 21728 3884 21792
rect 3948 21728 3964 21792
rect 4028 21728 4044 21792
rect 4108 21728 4124 21792
rect 4188 21728 4194 21792
rect 3878 21727 4194 21728
rect 10847 21792 11163 21793
rect 10847 21728 10853 21792
rect 10917 21728 10933 21792
rect 10997 21728 11013 21792
rect 11077 21728 11093 21792
rect 11157 21728 11163 21792
rect 10847 21727 11163 21728
rect 17816 21792 18132 21793
rect 17816 21728 17822 21792
rect 17886 21728 17902 21792
rect 17966 21728 17982 21792
rect 18046 21728 18062 21792
rect 18126 21728 18132 21792
rect 17816 21727 18132 21728
rect 24785 21792 25101 21793
rect 24785 21728 24791 21792
rect 24855 21728 24871 21792
rect 24935 21728 24951 21792
rect 25015 21728 25031 21792
rect 25095 21728 25101 21792
rect 24785 21727 25101 21728
rect 11605 21450 11671 21453
rect 11881 21450 11947 21453
rect 16757 21450 16823 21453
rect 11605 21448 16823 21450
rect 11605 21392 11610 21448
rect 11666 21392 11886 21448
rect 11942 21392 16762 21448
rect 16818 21392 16823 21448
rect 11605 21390 16823 21392
rect 11605 21387 11671 21390
rect 11881 21387 11947 21390
rect 16757 21387 16823 21390
rect 7362 21248 7678 21249
rect 7362 21184 7368 21248
rect 7432 21184 7448 21248
rect 7512 21184 7528 21248
rect 7592 21184 7608 21248
rect 7672 21184 7678 21248
rect 7362 21183 7678 21184
rect 14331 21248 14647 21249
rect 14331 21184 14337 21248
rect 14401 21184 14417 21248
rect 14481 21184 14497 21248
rect 14561 21184 14577 21248
rect 14641 21184 14647 21248
rect 14331 21183 14647 21184
rect 21300 21248 21616 21249
rect 21300 21184 21306 21248
rect 21370 21184 21386 21248
rect 21450 21184 21466 21248
rect 21530 21184 21546 21248
rect 21610 21184 21616 21248
rect 21300 21183 21616 21184
rect 28269 21248 28585 21249
rect 28269 21184 28275 21248
rect 28339 21184 28355 21248
rect 28419 21184 28435 21248
rect 28499 21184 28515 21248
rect 28579 21184 28585 21248
rect 28269 21183 28585 21184
rect 9857 20906 9923 20909
rect 9857 20904 12450 20906
rect 9857 20848 9862 20904
rect 9918 20848 12450 20904
rect 9857 20846 12450 20848
rect 9857 20843 9923 20846
rect 12390 20770 12450 20846
rect 13486 20770 13492 20772
rect 12390 20710 13492 20770
rect 13486 20708 13492 20710
rect 13556 20770 13562 20772
rect 14089 20770 14155 20773
rect 13556 20768 14155 20770
rect 13556 20712 14094 20768
rect 14150 20712 14155 20768
rect 13556 20710 14155 20712
rect 13556 20708 13562 20710
rect 14089 20707 14155 20710
rect 3878 20704 4194 20705
rect 3878 20640 3884 20704
rect 3948 20640 3964 20704
rect 4028 20640 4044 20704
rect 4108 20640 4124 20704
rect 4188 20640 4194 20704
rect 3878 20639 4194 20640
rect 10847 20704 11163 20705
rect 10847 20640 10853 20704
rect 10917 20640 10933 20704
rect 10997 20640 11013 20704
rect 11077 20640 11093 20704
rect 11157 20640 11163 20704
rect 10847 20639 11163 20640
rect 17816 20704 18132 20705
rect 17816 20640 17822 20704
rect 17886 20640 17902 20704
rect 17966 20640 17982 20704
rect 18046 20640 18062 20704
rect 18126 20640 18132 20704
rect 17816 20639 18132 20640
rect 24785 20704 25101 20705
rect 24785 20640 24791 20704
rect 24855 20640 24871 20704
rect 24935 20640 24951 20704
rect 25015 20640 25031 20704
rect 25095 20640 25101 20704
rect 24785 20639 25101 20640
rect 5717 20498 5783 20501
rect 11053 20498 11119 20501
rect 5717 20496 11119 20498
rect 5717 20440 5722 20496
rect 5778 20440 11058 20496
rect 11114 20440 11119 20496
rect 5717 20438 11119 20440
rect 5717 20435 5783 20438
rect 11053 20435 11119 20438
rect 7362 20160 7678 20161
rect 7362 20096 7368 20160
rect 7432 20096 7448 20160
rect 7512 20096 7528 20160
rect 7592 20096 7608 20160
rect 7672 20096 7678 20160
rect 7362 20095 7678 20096
rect 14331 20160 14647 20161
rect 14331 20096 14337 20160
rect 14401 20096 14417 20160
rect 14481 20096 14497 20160
rect 14561 20096 14577 20160
rect 14641 20096 14647 20160
rect 14331 20095 14647 20096
rect 21300 20160 21616 20161
rect 21300 20096 21306 20160
rect 21370 20096 21386 20160
rect 21450 20096 21466 20160
rect 21530 20096 21546 20160
rect 21610 20096 21616 20160
rect 21300 20095 21616 20096
rect 28269 20160 28585 20161
rect 28269 20096 28275 20160
rect 28339 20096 28355 20160
rect 28419 20096 28435 20160
rect 28499 20096 28515 20160
rect 28579 20096 28585 20160
rect 28269 20095 28585 20096
rect 3878 19616 4194 19617
rect 3878 19552 3884 19616
rect 3948 19552 3964 19616
rect 4028 19552 4044 19616
rect 4108 19552 4124 19616
rect 4188 19552 4194 19616
rect 3878 19551 4194 19552
rect 10847 19616 11163 19617
rect 10847 19552 10853 19616
rect 10917 19552 10933 19616
rect 10997 19552 11013 19616
rect 11077 19552 11093 19616
rect 11157 19552 11163 19616
rect 10847 19551 11163 19552
rect 17816 19616 18132 19617
rect 17816 19552 17822 19616
rect 17886 19552 17902 19616
rect 17966 19552 17982 19616
rect 18046 19552 18062 19616
rect 18126 19552 18132 19616
rect 17816 19551 18132 19552
rect 24785 19616 25101 19617
rect 24785 19552 24791 19616
rect 24855 19552 24871 19616
rect 24935 19552 24951 19616
rect 25015 19552 25031 19616
rect 25095 19552 25101 19616
rect 24785 19551 25101 19552
rect 3601 19410 3667 19413
rect 6177 19410 6243 19413
rect 3601 19408 6243 19410
rect 3601 19352 3606 19408
rect 3662 19352 6182 19408
rect 6238 19352 6243 19408
rect 3601 19350 6243 19352
rect 3601 19347 3667 19350
rect 6177 19347 6243 19350
rect 21541 19274 21607 19277
rect 27613 19274 27679 19277
rect 21541 19272 27679 19274
rect 21541 19216 21546 19272
rect 21602 19216 27618 19272
rect 27674 19216 27679 19272
rect 21541 19214 27679 19216
rect 21541 19211 21607 19214
rect 27613 19211 27679 19214
rect 7362 19072 7678 19073
rect 7362 19008 7368 19072
rect 7432 19008 7448 19072
rect 7512 19008 7528 19072
rect 7592 19008 7608 19072
rect 7672 19008 7678 19072
rect 7362 19007 7678 19008
rect 14331 19072 14647 19073
rect 14331 19008 14337 19072
rect 14401 19008 14417 19072
rect 14481 19008 14497 19072
rect 14561 19008 14577 19072
rect 14641 19008 14647 19072
rect 14331 19007 14647 19008
rect 21300 19072 21616 19073
rect 21300 19008 21306 19072
rect 21370 19008 21386 19072
rect 21450 19008 21466 19072
rect 21530 19008 21546 19072
rect 21610 19008 21616 19072
rect 21300 19007 21616 19008
rect 28269 19072 28585 19073
rect 28269 19008 28275 19072
rect 28339 19008 28355 19072
rect 28419 19008 28435 19072
rect 28499 19008 28515 19072
rect 28579 19008 28585 19072
rect 28269 19007 28585 19008
rect 3878 18528 4194 18529
rect 3878 18464 3884 18528
rect 3948 18464 3964 18528
rect 4028 18464 4044 18528
rect 4108 18464 4124 18528
rect 4188 18464 4194 18528
rect 3878 18463 4194 18464
rect 10847 18528 11163 18529
rect 10847 18464 10853 18528
rect 10917 18464 10933 18528
rect 10997 18464 11013 18528
rect 11077 18464 11093 18528
rect 11157 18464 11163 18528
rect 10847 18463 11163 18464
rect 17816 18528 18132 18529
rect 17816 18464 17822 18528
rect 17886 18464 17902 18528
rect 17966 18464 17982 18528
rect 18046 18464 18062 18528
rect 18126 18464 18132 18528
rect 17816 18463 18132 18464
rect 24785 18528 25101 18529
rect 24785 18464 24791 18528
rect 24855 18464 24871 18528
rect 24935 18464 24951 18528
rect 25015 18464 25031 18528
rect 25095 18464 25101 18528
rect 24785 18463 25101 18464
rect 7362 17984 7678 17985
rect 7362 17920 7368 17984
rect 7432 17920 7448 17984
rect 7512 17920 7528 17984
rect 7592 17920 7608 17984
rect 7672 17920 7678 17984
rect 7362 17919 7678 17920
rect 14331 17984 14647 17985
rect 14331 17920 14337 17984
rect 14401 17920 14417 17984
rect 14481 17920 14497 17984
rect 14561 17920 14577 17984
rect 14641 17920 14647 17984
rect 14331 17919 14647 17920
rect 21300 17984 21616 17985
rect 21300 17920 21306 17984
rect 21370 17920 21386 17984
rect 21450 17920 21466 17984
rect 21530 17920 21546 17984
rect 21610 17920 21616 17984
rect 21300 17919 21616 17920
rect 28269 17984 28585 17985
rect 28269 17920 28275 17984
rect 28339 17920 28355 17984
rect 28419 17920 28435 17984
rect 28499 17920 28515 17984
rect 28579 17920 28585 17984
rect 28269 17919 28585 17920
rect 13353 17642 13419 17645
rect 14641 17642 14707 17645
rect 13353 17640 14707 17642
rect 13353 17584 13358 17640
rect 13414 17584 14646 17640
rect 14702 17584 14707 17640
rect 13353 17582 14707 17584
rect 13353 17579 13419 17582
rect 14641 17579 14707 17582
rect 3878 17440 4194 17441
rect 3878 17376 3884 17440
rect 3948 17376 3964 17440
rect 4028 17376 4044 17440
rect 4108 17376 4124 17440
rect 4188 17376 4194 17440
rect 3878 17375 4194 17376
rect 10847 17440 11163 17441
rect 10847 17376 10853 17440
rect 10917 17376 10933 17440
rect 10997 17376 11013 17440
rect 11077 17376 11093 17440
rect 11157 17376 11163 17440
rect 10847 17375 11163 17376
rect 17816 17440 18132 17441
rect 17816 17376 17822 17440
rect 17886 17376 17902 17440
rect 17966 17376 17982 17440
rect 18046 17376 18062 17440
rect 18126 17376 18132 17440
rect 17816 17375 18132 17376
rect 24785 17440 25101 17441
rect 24785 17376 24791 17440
rect 24855 17376 24871 17440
rect 24935 17376 24951 17440
rect 25015 17376 25031 17440
rect 25095 17376 25101 17440
rect 24785 17375 25101 17376
rect 12985 17098 13051 17101
rect 16849 17098 16915 17101
rect 12985 17096 16915 17098
rect 12985 17040 12990 17096
rect 13046 17040 16854 17096
rect 16910 17040 16915 17096
rect 12985 17038 16915 17040
rect 12985 17035 13051 17038
rect 16849 17035 16915 17038
rect 7362 16896 7678 16897
rect 7362 16832 7368 16896
rect 7432 16832 7448 16896
rect 7512 16832 7528 16896
rect 7592 16832 7608 16896
rect 7672 16832 7678 16896
rect 7362 16831 7678 16832
rect 14331 16896 14647 16897
rect 14331 16832 14337 16896
rect 14401 16832 14417 16896
rect 14481 16832 14497 16896
rect 14561 16832 14577 16896
rect 14641 16832 14647 16896
rect 14331 16831 14647 16832
rect 21300 16896 21616 16897
rect 21300 16832 21306 16896
rect 21370 16832 21386 16896
rect 21450 16832 21466 16896
rect 21530 16832 21546 16896
rect 21610 16832 21616 16896
rect 21300 16831 21616 16832
rect 28269 16896 28585 16897
rect 28269 16832 28275 16896
rect 28339 16832 28355 16896
rect 28419 16832 28435 16896
rect 28499 16832 28515 16896
rect 28579 16832 28585 16896
rect 28269 16831 28585 16832
rect 13445 16420 13511 16421
rect 13445 16416 13492 16420
rect 13556 16418 13562 16420
rect 13445 16360 13450 16416
rect 13445 16356 13492 16360
rect 13556 16358 13602 16418
rect 13556 16356 13562 16358
rect 13445 16355 13511 16356
rect 3878 16352 4194 16353
rect 3878 16288 3884 16352
rect 3948 16288 3964 16352
rect 4028 16288 4044 16352
rect 4108 16288 4124 16352
rect 4188 16288 4194 16352
rect 3878 16287 4194 16288
rect 10847 16352 11163 16353
rect 10847 16288 10853 16352
rect 10917 16288 10933 16352
rect 10997 16288 11013 16352
rect 11077 16288 11093 16352
rect 11157 16288 11163 16352
rect 10847 16287 11163 16288
rect 17816 16352 18132 16353
rect 17816 16288 17822 16352
rect 17886 16288 17902 16352
rect 17966 16288 17982 16352
rect 18046 16288 18062 16352
rect 18126 16288 18132 16352
rect 17816 16287 18132 16288
rect 24785 16352 25101 16353
rect 24785 16288 24791 16352
rect 24855 16288 24871 16352
rect 24935 16288 24951 16352
rect 25015 16288 25031 16352
rect 25095 16288 25101 16352
rect 24785 16287 25101 16288
rect 15745 16146 15811 16149
rect 17769 16146 17835 16149
rect 15745 16144 17835 16146
rect 15745 16088 15750 16144
rect 15806 16088 17774 16144
rect 17830 16088 17835 16144
rect 15745 16086 17835 16088
rect 15745 16083 15811 16086
rect 17769 16083 17835 16086
rect 15929 16010 15995 16013
rect 17861 16010 17927 16013
rect 15929 16008 17927 16010
rect 15929 15952 15934 16008
rect 15990 15952 17866 16008
rect 17922 15952 17927 16008
rect 15929 15950 17927 15952
rect 15929 15947 15995 15950
rect 17861 15947 17927 15950
rect 7362 15808 7678 15809
rect 7362 15744 7368 15808
rect 7432 15744 7448 15808
rect 7512 15744 7528 15808
rect 7592 15744 7608 15808
rect 7672 15744 7678 15808
rect 7362 15743 7678 15744
rect 14331 15808 14647 15809
rect 14331 15744 14337 15808
rect 14401 15744 14417 15808
rect 14481 15744 14497 15808
rect 14561 15744 14577 15808
rect 14641 15744 14647 15808
rect 14331 15743 14647 15744
rect 21300 15808 21616 15809
rect 21300 15744 21306 15808
rect 21370 15744 21386 15808
rect 21450 15744 21466 15808
rect 21530 15744 21546 15808
rect 21610 15744 21616 15808
rect 21300 15743 21616 15744
rect 28269 15808 28585 15809
rect 28269 15744 28275 15808
rect 28339 15744 28355 15808
rect 28419 15744 28435 15808
rect 28499 15744 28515 15808
rect 28579 15744 28585 15808
rect 28269 15743 28585 15744
rect 3878 15264 4194 15265
rect 3878 15200 3884 15264
rect 3948 15200 3964 15264
rect 4028 15200 4044 15264
rect 4108 15200 4124 15264
rect 4188 15200 4194 15264
rect 3878 15199 4194 15200
rect 10847 15264 11163 15265
rect 10847 15200 10853 15264
rect 10917 15200 10933 15264
rect 10997 15200 11013 15264
rect 11077 15200 11093 15264
rect 11157 15200 11163 15264
rect 10847 15199 11163 15200
rect 17816 15264 18132 15265
rect 17816 15200 17822 15264
rect 17886 15200 17902 15264
rect 17966 15200 17982 15264
rect 18046 15200 18062 15264
rect 18126 15200 18132 15264
rect 17816 15199 18132 15200
rect 24785 15264 25101 15265
rect 24785 15200 24791 15264
rect 24855 15200 24871 15264
rect 24935 15200 24951 15264
rect 25015 15200 25031 15264
rect 25095 15200 25101 15264
rect 24785 15199 25101 15200
rect 10317 14922 10383 14925
rect 11697 14922 11763 14925
rect 10317 14920 11763 14922
rect 10317 14864 10322 14920
rect 10378 14864 11702 14920
rect 11758 14864 11763 14920
rect 10317 14862 11763 14864
rect 10317 14859 10383 14862
rect 11697 14859 11763 14862
rect 7362 14720 7678 14721
rect 7362 14656 7368 14720
rect 7432 14656 7448 14720
rect 7512 14656 7528 14720
rect 7592 14656 7608 14720
rect 7672 14656 7678 14720
rect 7362 14655 7678 14656
rect 14331 14720 14647 14721
rect 14331 14656 14337 14720
rect 14401 14656 14417 14720
rect 14481 14656 14497 14720
rect 14561 14656 14577 14720
rect 14641 14656 14647 14720
rect 14331 14655 14647 14656
rect 21300 14720 21616 14721
rect 21300 14656 21306 14720
rect 21370 14656 21386 14720
rect 21450 14656 21466 14720
rect 21530 14656 21546 14720
rect 21610 14656 21616 14720
rect 21300 14655 21616 14656
rect 28269 14720 28585 14721
rect 28269 14656 28275 14720
rect 28339 14656 28355 14720
rect 28419 14656 28435 14720
rect 28499 14656 28515 14720
rect 28579 14656 28585 14720
rect 28269 14655 28585 14656
rect 3878 14176 4194 14177
rect 3878 14112 3884 14176
rect 3948 14112 3964 14176
rect 4028 14112 4044 14176
rect 4108 14112 4124 14176
rect 4188 14112 4194 14176
rect 3878 14111 4194 14112
rect 10847 14176 11163 14177
rect 10847 14112 10853 14176
rect 10917 14112 10933 14176
rect 10997 14112 11013 14176
rect 11077 14112 11093 14176
rect 11157 14112 11163 14176
rect 10847 14111 11163 14112
rect 17816 14176 18132 14177
rect 17816 14112 17822 14176
rect 17886 14112 17902 14176
rect 17966 14112 17982 14176
rect 18046 14112 18062 14176
rect 18126 14112 18132 14176
rect 17816 14111 18132 14112
rect 24785 14176 25101 14177
rect 24785 14112 24791 14176
rect 24855 14112 24871 14176
rect 24935 14112 24951 14176
rect 25015 14112 25031 14176
rect 25095 14112 25101 14176
rect 24785 14111 25101 14112
rect 7362 13632 7678 13633
rect 7362 13568 7368 13632
rect 7432 13568 7448 13632
rect 7512 13568 7528 13632
rect 7592 13568 7608 13632
rect 7672 13568 7678 13632
rect 7362 13567 7678 13568
rect 14331 13632 14647 13633
rect 14331 13568 14337 13632
rect 14401 13568 14417 13632
rect 14481 13568 14497 13632
rect 14561 13568 14577 13632
rect 14641 13568 14647 13632
rect 14331 13567 14647 13568
rect 21300 13632 21616 13633
rect 21300 13568 21306 13632
rect 21370 13568 21386 13632
rect 21450 13568 21466 13632
rect 21530 13568 21546 13632
rect 21610 13568 21616 13632
rect 21300 13567 21616 13568
rect 28269 13632 28585 13633
rect 28269 13568 28275 13632
rect 28339 13568 28355 13632
rect 28419 13568 28435 13632
rect 28499 13568 28515 13632
rect 28579 13568 28585 13632
rect 28269 13567 28585 13568
rect 3878 13088 4194 13089
rect 3878 13024 3884 13088
rect 3948 13024 3964 13088
rect 4028 13024 4044 13088
rect 4108 13024 4124 13088
rect 4188 13024 4194 13088
rect 3878 13023 4194 13024
rect 10847 13088 11163 13089
rect 10847 13024 10853 13088
rect 10917 13024 10933 13088
rect 10997 13024 11013 13088
rect 11077 13024 11093 13088
rect 11157 13024 11163 13088
rect 10847 13023 11163 13024
rect 17816 13088 18132 13089
rect 17816 13024 17822 13088
rect 17886 13024 17902 13088
rect 17966 13024 17982 13088
rect 18046 13024 18062 13088
rect 18126 13024 18132 13088
rect 17816 13023 18132 13024
rect 24785 13088 25101 13089
rect 24785 13024 24791 13088
rect 24855 13024 24871 13088
rect 24935 13024 24951 13088
rect 25015 13024 25031 13088
rect 25095 13024 25101 13088
rect 24785 13023 25101 13024
rect 13445 12882 13511 12885
rect 16297 12882 16363 12885
rect 13445 12880 16363 12882
rect 13445 12824 13450 12880
rect 13506 12824 16302 12880
rect 16358 12824 16363 12880
rect 13445 12822 16363 12824
rect 13445 12819 13511 12822
rect 16297 12819 16363 12822
rect 13905 12746 13971 12749
rect 13905 12744 15026 12746
rect 13905 12688 13910 12744
rect 13966 12688 15026 12744
rect 13905 12686 15026 12688
rect 13905 12683 13971 12686
rect 14966 12613 15026 12686
rect 14966 12608 15075 12613
rect 14966 12552 15014 12608
rect 15070 12552 15075 12608
rect 14966 12550 15075 12552
rect 15009 12547 15075 12550
rect 7362 12544 7678 12545
rect 7362 12480 7368 12544
rect 7432 12480 7448 12544
rect 7512 12480 7528 12544
rect 7592 12480 7608 12544
rect 7672 12480 7678 12544
rect 7362 12479 7678 12480
rect 14331 12544 14647 12545
rect 14331 12480 14337 12544
rect 14401 12480 14417 12544
rect 14481 12480 14497 12544
rect 14561 12480 14577 12544
rect 14641 12480 14647 12544
rect 14331 12479 14647 12480
rect 21300 12544 21616 12545
rect 21300 12480 21306 12544
rect 21370 12480 21386 12544
rect 21450 12480 21466 12544
rect 21530 12480 21546 12544
rect 21610 12480 21616 12544
rect 21300 12479 21616 12480
rect 28269 12544 28585 12545
rect 28269 12480 28275 12544
rect 28339 12480 28355 12544
rect 28419 12480 28435 12544
rect 28499 12480 28515 12544
rect 28579 12480 28585 12544
rect 28269 12479 28585 12480
rect 3878 12000 4194 12001
rect 3878 11936 3884 12000
rect 3948 11936 3964 12000
rect 4028 11936 4044 12000
rect 4108 11936 4124 12000
rect 4188 11936 4194 12000
rect 3878 11935 4194 11936
rect 10847 12000 11163 12001
rect 10847 11936 10853 12000
rect 10917 11936 10933 12000
rect 10997 11936 11013 12000
rect 11077 11936 11093 12000
rect 11157 11936 11163 12000
rect 10847 11935 11163 11936
rect 17816 12000 18132 12001
rect 17816 11936 17822 12000
rect 17886 11936 17902 12000
rect 17966 11936 17982 12000
rect 18046 11936 18062 12000
rect 18126 11936 18132 12000
rect 17816 11935 18132 11936
rect 24785 12000 25101 12001
rect 24785 11936 24791 12000
rect 24855 11936 24871 12000
rect 24935 11936 24951 12000
rect 25015 11936 25031 12000
rect 25095 11936 25101 12000
rect 24785 11935 25101 11936
rect 7362 11456 7678 11457
rect 7362 11392 7368 11456
rect 7432 11392 7448 11456
rect 7512 11392 7528 11456
rect 7592 11392 7608 11456
rect 7672 11392 7678 11456
rect 7362 11391 7678 11392
rect 14331 11456 14647 11457
rect 14331 11392 14337 11456
rect 14401 11392 14417 11456
rect 14481 11392 14497 11456
rect 14561 11392 14577 11456
rect 14641 11392 14647 11456
rect 14331 11391 14647 11392
rect 21300 11456 21616 11457
rect 21300 11392 21306 11456
rect 21370 11392 21386 11456
rect 21450 11392 21466 11456
rect 21530 11392 21546 11456
rect 21610 11392 21616 11456
rect 21300 11391 21616 11392
rect 28269 11456 28585 11457
rect 28269 11392 28275 11456
rect 28339 11392 28355 11456
rect 28419 11392 28435 11456
rect 28499 11392 28515 11456
rect 28579 11392 28585 11456
rect 28269 11391 28585 11392
rect 3878 10912 4194 10913
rect 3878 10848 3884 10912
rect 3948 10848 3964 10912
rect 4028 10848 4044 10912
rect 4108 10848 4124 10912
rect 4188 10848 4194 10912
rect 3878 10847 4194 10848
rect 10847 10912 11163 10913
rect 10847 10848 10853 10912
rect 10917 10848 10933 10912
rect 10997 10848 11013 10912
rect 11077 10848 11093 10912
rect 11157 10848 11163 10912
rect 10847 10847 11163 10848
rect 17816 10912 18132 10913
rect 17816 10848 17822 10912
rect 17886 10848 17902 10912
rect 17966 10848 17982 10912
rect 18046 10848 18062 10912
rect 18126 10848 18132 10912
rect 17816 10847 18132 10848
rect 24785 10912 25101 10913
rect 24785 10848 24791 10912
rect 24855 10848 24871 10912
rect 24935 10848 24951 10912
rect 25015 10848 25031 10912
rect 25095 10848 25101 10912
rect 24785 10847 25101 10848
rect 7362 10368 7678 10369
rect 7362 10304 7368 10368
rect 7432 10304 7448 10368
rect 7512 10304 7528 10368
rect 7592 10304 7608 10368
rect 7672 10304 7678 10368
rect 7362 10303 7678 10304
rect 14331 10368 14647 10369
rect 14331 10304 14337 10368
rect 14401 10304 14417 10368
rect 14481 10304 14497 10368
rect 14561 10304 14577 10368
rect 14641 10304 14647 10368
rect 14331 10303 14647 10304
rect 21300 10368 21616 10369
rect 21300 10304 21306 10368
rect 21370 10304 21386 10368
rect 21450 10304 21466 10368
rect 21530 10304 21546 10368
rect 21610 10304 21616 10368
rect 21300 10303 21616 10304
rect 28269 10368 28585 10369
rect 28269 10304 28275 10368
rect 28339 10304 28355 10368
rect 28419 10304 28435 10368
rect 28499 10304 28515 10368
rect 28579 10304 28585 10368
rect 28269 10303 28585 10304
rect 3878 9824 4194 9825
rect 3878 9760 3884 9824
rect 3948 9760 3964 9824
rect 4028 9760 4044 9824
rect 4108 9760 4124 9824
rect 4188 9760 4194 9824
rect 3878 9759 4194 9760
rect 10847 9824 11163 9825
rect 10847 9760 10853 9824
rect 10917 9760 10933 9824
rect 10997 9760 11013 9824
rect 11077 9760 11093 9824
rect 11157 9760 11163 9824
rect 10847 9759 11163 9760
rect 17816 9824 18132 9825
rect 17816 9760 17822 9824
rect 17886 9760 17902 9824
rect 17966 9760 17982 9824
rect 18046 9760 18062 9824
rect 18126 9760 18132 9824
rect 17816 9759 18132 9760
rect 24785 9824 25101 9825
rect 24785 9760 24791 9824
rect 24855 9760 24871 9824
rect 24935 9760 24951 9824
rect 25015 9760 25031 9824
rect 25095 9760 25101 9824
rect 24785 9759 25101 9760
rect 7362 9280 7678 9281
rect 7362 9216 7368 9280
rect 7432 9216 7448 9280
rect 7512 9216 7528 9280
rect 7592 9216 7608 9280
rect 7672 9216 7678 9280
rect 7362 9215 7678 9216
rect 14331 9280 14647 9281
rect 14331 9216 14337 9280
rect 14401 9216 14417 9280
rect 14481 9216 14497 9280
rect 14561 9216 14577 9280
rect 14641 9216 14647 9280
rect 14331 9215 14647 9216
rect 21300 9280 21616 9281
rect 21300 9216 21306 9280
rect 21370 9216 21386 9280
rect 21450 9216 21466 9280
rect 21530 9216 21546 9280
rect 21610 9216 21616 9280
rect 21300 9215 21616 9216
rect 28269 9280 28585 9281
rect 28269 9216 28275 9280
rect 28339 9216 28355 9280
rect 28419 9216 28435 9280
rect 28499 9216 28515 9280
rect 28579 9216 28585 9280
rect 28269 9215 28585 9216
rect 3878 8736 4194 8737
rect 3878 8672 3884 8736
rect 3948 8672 3964 8736
rect 4028 8672 4044 8736
rect 4108 8672 4124 8736
rect 4188 8672 4194 8736
rect 3878 8671 4194 8672
rect 10847 8736 11163 8737
rect 10847 8672 10853 8736
rect 10917 8672 10933 8736
rect 10997 8672 11013 8736
rect 11077 8672 11093 8736
rect 11157 8672 11163 8736
rect 10847 8671 11163 8672
rect 17816 8736 18132 8737
rect 17816 8672 17822 8736
rect 17886 8672 17902 8736
rect 17966 8672 17982 8736
rect 18046 8672 18062 8736
rect 18126 8672 18132 8736
rect 17816 8671 18132 8672
rect 24785 8736 25101 8737
rect 24785 8672 24791 8736
rect 24855 8672 24871 8736
rect 24935 8672 24951 8736
rect 25015 8672 25031 8736
rect 25095 8672 25101 8736
rect 24785 8671 25101 8672
rect 7362 8192 7678 8193
rect 7362 8128 7368 8192
rect 7432 8128 7448 8192
rect 7512 8128 7528 8192
rect 7592 8128 7608 8192
rect 7672 8128 7678 8192
rect 7362 8127 7678 8128
rect 14331 8192 14647 8193
rect 14331 8128 14337 8192
rect 14401 8128 14417 8192
rect 14481 8128 14497 8192
rect 14561 8128 14577 8192
rect 14641 8128 14647 8192
rect 14331 8127 14647 8128
rect 21300 8192 21616 8193
rect 21300 8128 21306 8192
rect 21370 8128 21386 8192
rect 21450 8128 21466 8192
rect 21530 8128 21546 8192
rect 21610 8128 21616 8192
rect 21300 8127 21616 8128
rect 28269 8192 28585 8193
rect 28269 8128 28275 8192
rect 28339 8128 28355 8192
rect 28419 8128 28435 8192
rect 28499 8128 28515 8192
rect 28579 8128 28585 8192
rect 28269 8127 28585 8128
rect 3878 7648 4194 7649
rect 3878 7584 3884 7648
rect 3948 7584 3964 7648
rect 4028 7584 4044 7648
rect 4108 7584 4124 7648
rect 4188 7584 4194 7648
rect 3878 7583 4194 7584
rect 10847 7648 11163 7649
rect 10847 7584 10853 7648
rect 10917 7584 10933 7648
rect 10997 7584 11013 7648
rect 11077 7584 11093 7648
rect 11157 7584 11163 7648
rect 10847 7583 11163 7584
rect 17816 7648 18132 7649
rect 17816 7584 17822 7648
rect 17886 7584 17902 7648
rect 17966 7584 17982 7648
rect 18046 7584 18062 7648
rect 18126 7584 18132 7648
rect 17816 7583 18132 7584
rect 24785 7648 25101 7649
rect 24785 7584 24791 7648
rect 24855 7584 24871 7648
rect 24935 7584 24951 7648
rect 25015 7584 25031 7648
rect 25095 7584 25101 7648
rect 24785 7583 25101 7584
rect 7362 7104 7678 7105
rect 7362 7040 7368 7104
rect 7432 7040 7448 7104
rect 7512 7040 7528 7104
rect 7592 7040 7608 7104
rect 7672 7040 7678 7104
rect 7362 7039 7678 7040
rect 14331 7104 14647 7105
rect 14331 7040 14337 7104
rect 14401 7040 14417 7104
rect 14481 7040 14497 7104
rect 14561 7040 14577 7104
rect 14641 7040 14647 7104
rect 14331 7039 14647 7040
rect 21300 7104 21616 7105
rect 21300 7040 21306 7104
rect 21370 7040 21386 7104
rect 21450 7040 21466 7104
rect 21530 7040 21546 7104
rect 21610 7040 21616 7104
rect 21300 7039 21616 7040
rect 28269 7104 28585 7105
rect 28269 7040 28275 7104
rect 28339 7040 28355 7104
rect 28419 7040 28435 7104
rect 28499 7040 28515 7104
rect 28579 7040 28585 7104
rect 28269 7039 28585 7040
rect 3878 6560 4194 6561
rect 3878 6496 3884 6560
rect 3948 6496 3964 6560
rect 4028 6496 4044 6560
rect 4108 6496 4124 6560
rect 4188 6496 4194 6560
rect 3878 6495 4194 6496
rect 10847 6560 11163 6561
rect 10847 6496 10853 6560
rect 10917 6496 10933 6560
rect 10997 6496 11013 6560
rect 11077 6496 11093 6560
rect 11157 6496 11163 6560
rect 10847 6495 11163 6496
rect 17816 6560 18132 6561
rect 17816 6496 17822 6560
rect 17886 6496 17902 6560
rect 17966 6496 17982 6560
rect 18046 6496 18062 6560
rect 18126 6496 18132 6560
rect 17816 6495 18132 6496
rect 24785 6560 25101 6561
rect 24785 6496 24791 6560
rect 24855 6496 24871 6560
rect 24935 6496 24951 6560
rect 25015 6496 25031 6560
rect 25095 6496 25101 6560
rect 24785 6495 25101 6496
rect 7362 6016 7678 6017
rect 7362 5952 7368 6016
rect 7432 5952 7448 6016
rect 7512 5952 7528 6016
rect 7592 5952 7608 6016
rect 7672 5952 7678 6016
rect 7362 5951 7678 5952
rect 14331 6016 14647 6017
rect 14331 5952 14337 6016
rect 14401 5952 14417 6016
rect 14481 5952 14497 6016
rect 14561 5952 14577 6016
rect 14641 5952 14647 6016
rect 14331 5951 14647 5952
rect 21300 6016 21616 6017
rect 21300 5952 21306 6016
rect 21370 5952 21386 6016
rect 21450 5952 21466 6016
rect 21530 5952 21546 6016
rect 21610 5952 21616 6016
rect 21300 5951 21616 5952
rect 28269 6016 28585 6017
rect 28269 5952 28275 6016
rect 28339 5952 28355 6016
rect 28419 5952 28435 6016
rect 28499 5952 28515 6016
rect 28579 5952 28585 6016
rect 28269 5951 28585 5952
rect 3878 5472 4194 5473
rect 3878 5408 3884 5472
rect 3948 5408 3964 5472
rect 4028 5408 4044 5472
rect 4108 5408 4124 5472
rect 4188 5408 4194 5472
rect 3878 5407 4194 5408
rect 10847 5472 11163 5473
rect 10847 5408 10853 5472
rect 10917 5408 10933 5472
rect 10997 5408 11013 5472
rect 11077 5408 11093 5472
rect 11157 5408 11163 5472
rect 10847 5407 11163 5408
rect 17816 5472 18132 5473
rect 17816 5408 17822 5472
rect 17886 5408 17902 5472
rect 17966 5408 17982 5472
rect 18046 5408 18062 5472
rect 18126 5408 18132 5472
rect 17816 5407 18132 5408
rect 24785 5472 25101 5473
rect 24785 5408 24791 5472
rect 24855 5408 24871 5472
rect 24935 5408 24951 5472
rect 25015 5408 25031 5472
rect 25095 5408 25101 5472
rect 24785 5407 25101 5408
rect 7362 4928 7678 4929
rect 7362 4864 7368 4928
rect 7432 4864 7448 4928
rect 7512 4864 7528 4928
rect 7592 4864 7608 4928
rect 7672 4864 7678 4928
rect 7362 4863 7678 4864
rect 14331 4928 14647 4929
rect 14331 4864 14337 4928
rect 14401 4864 14417 4928
rect 14481 4864 14497 4928
rect 14561 4864 14577 4928
rect 14641 4864 14647 4928
rect 14331 4863 14647 4864
rect 21300 4928 21616 4929
rect 21300 4864 21306 4928
rect 21370 4864 21386 4928
rect 21450 4864 21466 4928
rect 21530 4864 21546 4928
rect 21610 4864 21616 4928
rect 21300 4863 21616 4864
rect 28269 4928 28585 4929
rect 28269 4864 28275 4928
rect 28339 4864 28355 4928
rect 28419 4864 28435 4928
rect 28499 4864 28515 4928
rect 28579 4864 28585 4928
rect 28269 4863 28585 4864
rect 3878 4384 4194 4385
rect 3878 4320 3884 4384
rect 3948 4320 3964 4384
rect 4028 4320 4044 4384
rect 4108 4320 4124 4384
rect 4188 4320 4194 4384
rect 3878 4319 4194 4320
rect 10847 4384 11163 4385
rect 10847 4320 10853 4384
rect 10917 4320 10933 4384
rect 10997 4320 11013 4384
rect 11077 4320 11093 4384
rect 11157 4320 11163 4384
rect 10847 4319 11163 4320
rect 17816 4384 18132 4385
rect 17816 4320 17822 4384
rect 17886 4320 17902 4384
rect 17966 4320 17982 4384
rect 18046 4320 18062 4384
rect 18126 4320 18132 4384
rect 17816 4319 18132 4320
rect 24785 4384 25101 4385
rect 24785 4320 24791 4384
rect 24855 4320 24871 4384
rect 24935 4320 24951 4384
rect 25015 4320 25031 4384
rect 25095 4320 25101 4384
rect 24785 4319 25101 4320
rect 7362 3840 7678 3841
rect 7362 3776 7368 3840
rect 7432 3776 7448 3840
rect 7512 3776 7528 3840
rect 7592 3776 7608 3840
rect 7672 3776 7678 3840
rect 7362 3775 7678 3776
rect 14331 3840 14647 3841
rect 14331 3776 14337 3840
rect 14401 3776 14417 3840
rect 14481 3776 14497 3840
rect 14561 3776 14577 3840
rect 14641 3776 14647 3840
rect 14331 3775 14647 3776
rect 21300 3840 21616 3841
rect 21300 3776 21306 3840
rect 21370 3776 21386 3840
rect 21450 3776 21466 3840
rect 21530 3776 21546 3840
rect 21610 3776 21616 3840
rect 21300 3775 21616 3776
rect 28269 3840 28585 3841
rect 28269 3776 28275 3840
rect 28339 3776 28355 3840
rect 28419 3776 28435 3840
rect 28499 3776 28515 3840
rect 28579 3776 28585 3840
rect 28269 3775 28585 3776
rect 3878 3296 4194 3297
rect 3878 3232 3884 3296
rect 3948 3232 3964 3296
rect 4028 3232 4044 3296
rect 4108 3232 4124 3296
rect 4188 3232 4194 3296
rect 3878 3231 4194 3232
rect 10847 3296 11163 3297
rect 10847 3232 10853 3296
rect 10917 3232 10933 3296
rect 10997 3232 11013 3296
rect 11077 3232 11093 3296
rect 11157 3232 11163 3296
rect 10847 3231 11163 3232
rect 17816 3296 18132 3297
rect 17816 3232 17822 3296
rect 17886 3232 17902 3296
rect 17966 3232 17982 3296
rect 18046 3232 18062 3296
rect 18126 3232 18132 3296
rect 17816 3231 18132 3232
rect 24785 3296 25101 3297
rect 24785 3232 24791 3296
rect 24855 3232 24871 3296
rect 24935 3232 24951 3296
rect 25015 3232 25031 3296
rect 25095 3232 25101 3296
rect 24785 3231 25101 3232
rect 7362 2752 7678 2753
rect 7362 2688 7368 2752
rect 7432 2688 7448 2752
rect 7512 2688 7528 2752
rect 7592 2688 7608 2752
rect 7672 2688 7678 2752
rect 7362 2687 7678 2688
rect 14331 2752 14647 2753
rect 14331 2688 14337 2752
rect 14401 2688 14417 2752
rect 14481 2688 14497 2752
rect 14561 2688 14577 2752
rect 14641 2688 14647 2752
rect 14331 2687 14647 2688
rect 21300 2752 21616 2753
rect 21300 2688 21306 2752
rect 21370 2688 21386 2752
rect 21450 2688 21466 2752
rect 21530 2688 21546 2752
rect 21610 2688 21616 2752
rect 21300 2687 21616 2688
rect 28269 2752 28585 2753
rect 28269 2688 28275 2752
rect 28339 2688 28355 2752
rect 28419 2688 28435 2752
rect 28499 2688 28515 2752
rect 28579 2688 28585 2752
rect 28269 2687 28585 2688
rect 3878 2208 4194 2209
rect 3878 2144 3884 2208
rect 3948 2144 3964 2208
rect 4028 2144 4044 2208
rect 4108 2144 4124 2208
rect 4188 2144 4194 2208
rect 3878 2143 4194 2144
rect 10847 2208 11163 2209
rect 10847 2144 10853 2208
rect 10917 2144 10933 2208
rect 10997 2144 11013 2208
rect 11077 2144 11093 2208
rect 11157 2144 11163 2208
rect 10847 2143 11163 2144
rect 17816 2208 18132 2209
rect 17816 2144 17822 2208
rect 17886 2144 17902 2208
rect 17966 2144 17982 2208
rect 18046 2144 18062 2208
rect 18126 2144 18132 2208
rect 17816 2143 18132 2144
rect 24785 2208 25101 2209
rect 24785 2144 24791 2208
rect 24855 2144 24871 2208
rect 24935 2144 24951 2208
rect 25015 2144 25031 2208
rect 25095 2144 25101 2208
rect 24785 2143 25101 2144
rect 7362 1664 7678 1665
rect 7362 1600 7368 1664
rect 7432 1600 7448 1664
rect 7512 1600 7528 1664
rect 7592 1600 7608 1664
rect 7672 1600 7678 1664
rect 7362 1599 7678 1600
rect 14331 1664 14647 1665
rect 14331 1600 14337 1664
rect 14401 1600 14417 1664
rect 14481 1600 14497 1664
rect 14561 1600 14577 1664
rect 14641 1600 14647 1664
rect 14331 1599 14647 1600
rect 21300 1664 21616 1665
rect 21300 1600 21306 1664
rect 21370 1600 21386 1664
rect 21450 1600 21466 1664
rect 21530 1600 21546 1664
rect 21610 1600 21616 1664
rect 21300 1599 21616 1600
rect 28269 1664 28585 1665
rect 28269 1600 28275 1664
rect 28339 1600 28355 1664
rect 28419 1600 28435 1664
rect 28499 1600 28515 1664
rect 28579 1600 28585 1664
rect 28269 1599 28585 1600
rect 3878 1120 4194 1121
rect 3878 1056 3884 1120
rect 3948 1056 3964 1120
rect 4028 1056 4044 1120
rect 4108 1056 4124 1120
rect 4188 1056 4194 1120
rect 3878 1055 4194 1056
rect 10847 1120 11163 1121
rect 10847 1056 10853 1120
rect 10917 1056 10933 1120
rect 10997 1056 11013 1120
rect 11077 1056 11093 1120
rect 11157 1056 11163 1120
rect 10847 1055 11163 1056
rect 17816 1120 18132 1121
rect 17816 1056 17822 1120
rect 17886 1056 17902 1120
rect 17966 1056 17982 1120
rect 18046 1056 18062 1120
rect 18126 1056 18132 1120
rect 17816 1055 18132 1056
rect 24785 1120 25101 1121
rect 24785 1056 24791 1120
rect 24855 1056 24871 1120
rect 24935 1056 24951 1120
rect 25015 1056 25031 1120
rect 25095 1056 25101 1120
rect 24785 1055 25101 1056
rect 7362 576 7678 577
rect 7362 512 7368 576
rect 7432 512 7448 576
rect 7512 512 7528 576
rect 7592 512 7608 576
rect 7672 512 7678 576
rect 7362 511 7678 512
rect 14331 576 14647 577
rect 14331 512 14337 576
rect 14401 512 14417 576
rect 14481 512 14497 576
rect 14561 512 14577 576
rect 14641 512 14647 576
rect 14331 511 14647 512
rect 21300 576 21616 577
rect 21300 512 21306 576
rect 21370 512 21386 576
rect 21450 512 21466 576
rect 21530 512 21546 576
rect 21610 512 21616 576
rect 21300 511 21616 512
rect 28269 576 28585 577
rect 28269 512 28275 576
rect 28339 512 28355 576
rect 28419 512 28435 576
rect 28499 512 28515 576
rect 28579 512 28585 576
rect 28269 511 28585 512
<< via3 >>
rect 3884 28316 3948 28320
rect 3884 28260 3888 28316
rect 3888 28260 3944 28316
rect 3944 28260 3948 28316
rect 3884 28256 3948 28260
rect 3964 28316 4028 28320
rect 3964 28260 3968 28316
rect 3968 28260 4024 28316
rect 4024 28260 4028 28316
rect 3964 28256 4028 28260
rect 4044 28316 4108 28320
rect 4044 28260 4048 28316
rect 4048 28260 4104 28316
rect 4104 28260 4108 28316
rect 4044 28256 4108 28260
rect 4124 28316 4188 28320
rect 4124 28260 4128 28316
rect 4128 28260 4184 28316
rect 4184 28260 4188 28316
rect 4124 28256 4188 28260
rect 10853 28316 10917 28320
rect 10853 28260 10857 28316
rect 10857 28260 10913 28316
rect 10913 28260 10917 28316
rect 10853 28256 10917 28260
rect 10933 28316 10997 28320
rect 10933 28260 10937 28316
rect 10937 28260 10993 28316
rect 10993 28260 10997 28316
rect 10933 28256 10997 28260
rect 11013 28316 11077 28320
rect 11013 28260 11017 28316
rect 11017 28260 11073 28316
rect 11073 28260 11077 28316
rect 11013 28256 11077 28260
rect 11093 28316 11157 28320
rect 11093 28260 11097 28316
rect 11097 28260 11153 28316
rect 11153 28260 11157 28316
rect 11093 28256 11157 28260
rect 17822 28316 17886 28320
rect 17822 28260 17826 28316
rect 17826 28260 17882 28316
rect 17882 28260 17886 28316
rect 17822 28256 17886 28260
rect 17902 28316 17966 28320
rect 17902 28260 17906 28316
rect 17906 28260 17962 28316
rect 17962 28260 17966 28316
rect 17902 28256 17966 28260
rect 17982 28316 18046 28320
rect 17982 28260 17986 28316
rect 17986 28260 18042 28316
rect 18042 28260 18046 28316
rect 17982 28256 18046 28260
rect 18062 28316 18126 28320
rect 18062 28260 18066 28316
rect 18066 28260 18122 28316
rect 18122 28260 18126 28316
rect 18062 28256 18126 28260
rect 24791 28316 24855 28320
rect 24791 28260 24795 28316
rect 24795 28260 24851 28316
rect 24851 28260 24855 28316
rect 24791 28256 24855 28260
rect 24871 28316 24935 28320
rect 24871 28260 24875 28316
rect 24875 28260 24931 28316
rect 24931 28260 24935 28316
rect 24871 28256 24935 28260
rect 24951 28316 25015 28320
rect 24951 28260 24955 28316
rect 24955 28260 25011 28316
rect 25011 28260 25015 28316
rect 24951 28256 25015 28260
rect 25031 28316 25095 28320
rect 25031 28260 25035 28316
rect 25035 28260 25091 28316
rect 25091 28260 25095 28316
rect 25031 28256 25095 28260
rect 7368 27772 7432 27776
rect 7368 27716 7372 27772
rect 7372 27716 7428 27772
rect 7428 27716 7432 27772
rect 7368 27712 7432 27716
rect 7448 27772 7512 27776
rect 7448 27716 7452 27772
rect 7452 27716 7508 27772
rect 7508 27716 7512 27772
rect 7448 27712 7512 27716
rect 7528 27772 7592 27776
rect 7528 27716 7532 27772
rect 7532 27716 7588 27772
rect 7588 27716 7592 27772
rect 7528 27712 7592 27716
rect 7608 27772 7672 27776
rect 7608 27716 7612 27772
rect 7612 27716 7668 27772
rect 7668 27716 7672 27772
rect 7608 27712 7672 27716
rect 14337 27772 14401 27776
rect 14337 27716 14341 27772
rect 14341 27716 14397 27772
rect 14397 27716 14401 27772
rect 14337 27712 14401 27716
rect 14417 27772 14481 27776
rect 14417 27716 14421 27772
rect 14421 27716 14477 27772
rect 14477 27716 14481 27772
rect 14417 27712 14481 27716
rect 14497 27772 14561 27776
rect 14497 27716 14501 27772
rect 14501 27716 14557 27772
rect 14557 27716 14561 27772
rect 14497 27712 14561 27716
rect 14577 27772 14641 27776
rect 14577 27716 14581 27772
rect 14581 27716 14637 27772
rect 14637 27716 14641 27772
rect 14577 27712 14641 27716
rect 21306 27772 21370 27776
rect 21306 27716 21310 27772
rect 21310 27716 21366 27772
rect 21366 27716 21370 27772
rect 21306 27712 21370 27716
rect 21386 27772 21450 27776
rect 21386 27716 21390 27772
rect 21390 27716 21446 27772
rect 21446 27716 21450 27772
rect 21386 27712 21450 27716
rect 21466 27772 21530 27776
rect 21466 27716 21470 27772
rect 21470 27716 21526 27772
rect 21526 27716 21530 27772
rect 21466 27712 21530 27716
rect 21546 27772 21610 27776
rect 21546 27716 21550 27772
rect 21550 27716 21606 27772
rect 21606 27716 21610 27772
rect 21546 27712 21610 27716
rect 28275 27772 28339 27776
rect 28275 27716 28279 27772
rect 28279 27716 28335 27772
rect 28335 27716 28339 27772
rect 28275 27712 28339 27716
rect 28355 27772 28419 27776
rect 28355 27716 28359 27772
rect 28359 27716 28415 27772
rect 28415 27716 28419 27772
rect 28355 27712 28419 27716
rect 28435 27772 28499 27776
rect 28435 27716 28439 27772
rect 28439 27716 28495 27772
rect 28495 27716 28499 27772
rect 28435 27712 28499 27716
rect 28515 27772 28579 27776
rect 28515 27716 28519 27772
rect 28519 27716 28575 27772
rect 28575 27716 28579 27772
rect 28515 27712 28579 27716
rect 3884 27228 3948 27232
rect 3884 27172 3888 27228
rect 3888 27172 3944 27228
rect 3944 27172 3948 27228
rect 3884 27168 3948 27172
rect 3964 27228 4028 27232
rect 3964 27172 3968 27228
rect 3968 27172 4024 27228
rect 4024 27172 4028 27228
rect 3964 27168 4028 27172
rect 4044 27228 4108 27232
rect 4044 27172 4048 27228
rect 4048 27172 4104 27228
rect 4104 27172 4108 27228
rect 4044 27168 4108 27172
rect 4124 27228 4188 27232
rect 4124 27172 4128 27228
rect 4128 27172 4184 27228
rect 4184 27172 4188 27228
rect 4124 27168 4188 27172
rect 10853 27228 10917 27232
rect 10853 27172 10857 27228
rect 10857 27172 10913 27228
rect 10913 27172 10917 27228
rect 10853 27168 10917 27172
rect 10933 27228 10997 27232
rect 10933 27172 10937 27228
rect 10937 27172 10993 27228
rect 10993 27172 10997 27228
rect 10933 27168 10997 27172
rect 11013 27228 11077 27232
rect 11013 27172 11017 27228
rect 11017 27172 11073 27228
rect 11073 27172 11077 27228
rect 11013 27168 11077 27172
rect 11093 27228 11157 27232
rect 11093 27172 11097 27228
rect 11097 27172 11153 27228
rect 11153 27172 11157 27228
rect 11093 27168 11157 27172
rect 17822 27228 17886 27232
rect 17822 27172 17826 27228
rect 17826 27172 17882 27228
rect 17882 27172 17886 27228
rect 17822 27168 17886 27172
rect 17902 27228 17966 27232
rect 17902 27172 17906 27228
rect 17906 27172 17962 27228
rect 17962 27172 17966 27228
rect 17902 27168 17966 27172
rect 17982 27228 18046 27232
rect 17982 27172 17986 27228
rect 17986 27172 18042 27228
rect 18042 27172 18046 27228
rect 17982 27168 18046 27172
rect 18062 27228 18126 27232
rect 18062 27172 18066 27228
rect 18066 27172 18122 27228
rect 18122 27172 18126 27228
rect 18062 27168 18126 27172
rect 24791 27228 24855 27232
rect 24791 27172 24795 27228
rect 24795 27172 24851 27228
rect 24851 27172 24855 27228
rect 24791 27168 24855 27172
rect 24871 27228 24935 27232
rect 24871 27172 24875 27228
rect 24875 27172 24931 27228
rect 24931 27172 24935 27228
rect 24871 27168 24935 27172
rect 24951 27228 25015 27232
rect 24951 27172 24955 27228
rect 24955 27172 25011 27228
rect 25011 27172 25015 27228
rect 24951 27168 25015 27172
rect 25031 27228 25095 27232
rect 25031 27172 25035 27228
rect 25035 27172 25091 27228
rect 25091 27172 25095 27228
rect 25031 27168 25095 27172
rect 7368 26684 7432 26688
rect 7368 26628 7372 26684
rect 7372 26628 7428 26684
rect 7428 26628 7432 26684
rect 7368 26624 7432 26628
rect 7448 26684 7512 26688
rect 7448 26628 7452 26684
rect 7452 26628 7508 26684
rect 7508 26628 7512 26684
rect 7448 26624 7512 26628
rect 7528 26684 7592 26688
rect 7528 26628 7532 26684
rect 7532 26628 7588 26684
rect 7588 26628 7592 26684
rect 7528 26624 7592 26628
rect 7608 26684 7672 26688
rect 7608 26628 7612 26684
rect 7612 26628 7668 26684
rect 7668 26628 7672 26684
rect 7608 26624 7672 26628
rect 14337 26684 14401 26688
rect 14337 26628 14341 26684
rect 14341 26628 14397 26684
rect 14397 26628 14401 26684
rect 14337 26624 14401 26628
rect 14417 26684 14481 26688
rect 14417 26628 14421 26684
rect 14421 26628 14477 26684
rect 14477 26628 14481 26684
rect 14417 26624 14481 26628
rect 14497 26684 14561 26688
rect 14497 26628 14501 26684
rect 14501 26628 14557 26684
rect 14557 26628 14561 26684
rect 14497 26624 14561 26628
rect 14577 26684 14641 26688
rect 14577 26628 14581 26684
rect 14581 26628 14637 26684
rect 14637 26628 14641 26684
rect 14577 26624 14641 26628
rect 21306 26684 21370 26688
rect 21306 26628 21310 26684
rect 21310 26628 21366 26684
rect 21366 26628 21370 26684
rect 21306 26624 21370 26628
rect 21386 26684 21450 26688
rect 21386 26628 21390 26684
rect 21390 26628 21446 26684
rect 21446 26628 21450 26684
rect 21386 26624 21450 26628
rect 21466 26684 21530 26688
rect 21466 26628 21470 26684
rect 21470 26628 21526 26684
rect 21526 26628 21530 26684
rect 21466 26624 21530 26628
rect 21546 26684 21610 26688
rect 21546 26628 21550 26684
rect 21550 26628 21606 26684
rect 21606 26628 21610 26684
rect 21546 26624 21610 26628
rect 28275 26684 28339 26688
rect 28275 26628 28279 26684
rect 28279 26628 28335 26684
rect 28335 26628 28339 26684
rect 28275 26624 28339 26628
rect 28355 26684 28419 26688
rect 28355 26628 28359 26684
rect 28359 26628 28415 26684
rect 28415 26628 28419 26684
rect 28355 26624 28419 26628
rect 28435 26684 28499 26688
rect 28435 26628 28439 26684
rect 28439 26628 28495 26684
rect 28495 26628 28499 26684
rect 28435 26624 28499 26628
rect 28515 26684 28579 26688
rect 28515 26628 28519 26684
rect 28519 26628 28575 26684
rect 28575 26628 28579 26684
rect 28515 26624 28579 26628
rect 3884 26140 3948 26144
rect 3884 26084 3888 26140
rect 3888 26084 3944 26140
rect 3944 26084 3948 26140
rect 3884 26080 3948 26084
rect 3964 26140 4028 26144
rect 3964 26084 3968 26140
rect 3968 26084 4024 26140
rect 4024 26084 4028 26140
rect 3964 26080 4028 26084
rect 4044 26140 4108 26144
rect 4044 26084 4048 26140
rect 4048 26084 4104 26140
rect 4104 26084 4108 26140
rect 4044 26080 4108 26084
rect 4124 26140 4188 26144
rect 4124 26084 4128 26140
rect 4128 26084 4184 26140
rect 4184 26084 4188 26140
rect 4124 26080 4188 26084
rect 10853 26140 10917 26144
rect 10853 26084 10857 26140
rect 10857 26084 10913 26140
rect 10913 26084 10917 26140
rect 10853 26080 10917 26084
rect 10933 26140 10997 26144
rect 10933 26084 10937 26140
rect 10937 26084 10993 26140
rect 10993 26084 10997 26140
rect 10933 26080 10997 26084
rect 11013 26140 11077 26144
rect 11013 26084 11017 26140
rect 11017 26084 11073 26140
rect 11073 26084 11077 26140
rect 11013 26080 11077 26084
rect 11093 26140 11157 26144
rect 11093 26084 11097 26140
rect 11097 26084 11153 26140
rect 11153 26084 11157 26140
rect 11093 26080 11157 26084
rect 17822 26140 17886 26144
rect 17822 26084 17826 26140
rect 17826 26084 17882 26140
rect 17882 26084 17886 26140
rect 17822 26080 17886 26084
rect 17902 26140 17966 26144
rect 17902 26084 17906 26140
rect 17906 26084 17962 26140
rect 17962 26084 17966 26140
rect 17902 26080 17966 26084
rect 17982 26140 18046 26144
rect 17982 26084 17986 26140
rect 17986 26084 18042 26140
rect 18042 26084 18046 26140
rect 17982 26080 18046 26084
rect 18062 26140 18126 26144
rect 18062 26084 18066 26140
rect 18066 26084 18122 26140
rect 18122 26084 18126 26140
rect 18062 26080 18126 26084
rect 24791 26140 24855 26144
rect 24791 26084 24795 26140
rect 24795 26084 24851 26140
rect 24851 26084 24855 26140
rect 24791 26080 24855 26084
rect 24871 26140 24935 26144
rect 24871 26084 24875 26140
rect 24875 26084 24931 26140
rect 24931 26084 24935 26140
rect 24871 26080 24935 26084
rect 24951 26140 25015 26144
rect 24951 26084 24955 26140
rect 24955 26084 25011 26140
rect 25011 26084 25015 26140
rect 24951 26080 25015 26084
rect 25031 26140 25095 26144
rect 25031 26084 25035 26140
rect 25035 26084 25091 26140
rect 25091 26084 25095 26140
rect 25031 26080 25095 26084
rect 7368 25596 7432 25600
rect 7368 25540 7372 25596
rect 7372 25540 7428 25596
rect 7428 25540 7432 25596
rect 7368 25536 7432 25540
rect 7448 25596 7512 25600
rect 7448 25540 7452 25596
rect 7452 25540 7508 25596
rect 7508 25540 7512 25596
rect 7448 25536 7512 25540
rect 7528 25596 7592 25600
rect 7528 25540 7532 25596
rect 7532 25540 7588 25596
rect 7588 25540 7592 25596
rect 7528 25536 7592 25540
rect 7608 25596 7672 25600
rect 7608 25540 7612 25596
rect 7612 25540 7668 25596
rect 7668 25540 7672 25596
rect 7608 25536 7672 25540
rect 14337 25596 14401 25600
rect 14337 25540 14341 25596
rect 14341 25540 14397 25596
rect 14397 25540 14401 25596
rect 14337 25536 14401 25540
rect 14417 25596 14481 25600
rect 14417 25540 14421 25596
rect 14421 25540 14477 25596
rect 14477 25540 14481 25596
rect 14417 25536 14481 25540
rect 14497 25596 14561 25600
rect 14497 25540 14501 25596
rect 14501 25540 14557 25596
rect 14557 25540 14561 25596
rect 14497 25536 14561 25540
rect 14577 25596 14641 25600
rect 14577 25540 14581 25596
rect 14581 25540 14637 25596
rect 14637 25540 14641 25596
rect 14577 25536 14641 25540
rect 21306 25596 21370 25600
rect 21306 25540 21310 25596
rect 21310 25540 21366 25596
rect 21366 25540 21370 25596
rect 21306 25536 21370 25540
rect 21386 25596 21450 25600
rect 21386 25540 21390 25596
rect 21390 25540 21446 25596
rect 21446 25540 21450 25596
rect 21386 25536 21450 25540
rect 21466 25596 21530 25600
rect 21466 25540 21470 25596
rect 21470 25540 21526 25596
rect 21526 25540 21530 25596
rect 21466 25536 21530 25540
rect 21546 25596 21610 25600
rect 21546 25540 21550 25596
rect 21550 25540 21606 25596
rect 21606 25540 21610 25596
rect 21546 25536 21610 25540
rect 28275 25596 28339 25600
rect 28275 25540 28279 25596
rect 28279 25540 28335 25596
rect 28335 25540 28339 25596
rect 28275 25536 28339 25540
rect 28355 25596 28419 25600
rect 28355 25540 28359 25596
rect 28359 25540 28415 25596
rect 28415 25540 28419 25596
rect 28355 25536 28419 25540
rect 28435 25596 28499 25600
rect 28435 25540 28439 25596
rect 28439 25540 28495 25596
rect 28495 25540 28499 25596
rect 28435 25536 28499 25540
rect 28515 25596 28579 25600
rect 28515 25540 28519 25596
rect 28519 25540 28575 25596
rect 28575 25540 28579 25596
rect 28515 25536 28579 25540
rect 3884 25052 3948 25056
rect 3884 24996 3888 25052
rect 3888 24996 3944 25052
rect 3944 24996 3948 25052
rect 3884 24992 3948 24996
rect 3964 25052 4028 25056
rect 3964 24996 3968 25052
rect 3968 24996 4024 25052
rect 4024 24996 4028 25052
rect 3964 24992 4028 24996
rect 4044 25052 4108 25056
rect 4044 24996 4048 25052
rect 4048 24996 4104 25052
rect 4104 24996 4108 25052
rect 4044 24992 4108 24996
rect 4124 25052 4188 25056
rect 4124 24996 4128 25052
rect 4128 24996 4184 25052
rect 4184 24996 4188 25052
rect 4124 24992 4188 24996
rect 10853 25052 10917 25056
rect 10853 24996 10857 25052
rect 10857 24996 10913 25052
rect 10913 24996 10917 25052
rect 10853 24992 10917 24996
rect 10933 25052 10997 25056
rect 10933 24996 10937 25052
rect 10937 24996 10993 25052
rect 10993 24996 10997 25052
rect 10933 24992 10997 24996
rect 11013 25052 11077 25056
rect 11013 24996 11017 25052
rect 11017 24996 11073 25052
rect 11073 24996 11077 25052
rect 11013 24992 11077 24996
rect 11093 25052 11157 25056
rect 11093 24996 11097 25052
rect 11097 24996 11153 25052
rect 11153 24996 11157 25052
rect 11093 24992 11157 24996
rect 17822 25052 17886 25056
rect 17822 24996 17826 25052
rect 17826 24996 17882 25052
rect 17882 24996 17886 25052
rect 17822 24992 17886 24996
rect 17902 25052 17966 25056
rect 17902 24996 17906 25052
rect 17906 24996 17962 25052
rect 17962 24996 17966 25052
rect 17902 24992 17966 24996
rect 17982 25052 18046 25056
rect 17982 24996 17986 25052
rect 17986 24996 18042 25052
rect 18042 24996 18046 25052
rect 17982 24992 18046 24996
rect 18062 25052 18126 25056
rect 18062 24996 18066 25052
rect 18066 24996 18122 25052
rect 18122 24996 18126 25052
rect 18062 24992 18126 24996
rect 24791 25052 24855 25056
rect 24791 24996 24795 25052
rect 24795 24996 24851 25052
rect 24851 24996 24855 25052
rect 24791 24992 24855 24996
rect 24871 25052 24935 25056
rect 24871 24996 24875 25052
rect 24875 24996 24931 25052
rect 24931 24996 24935 25052
rect 24871 24992 24935 24996
rect 24951 25052 25015 25056
rect 24951 24996 24955 25052
rect 24955 24996 25011 25052
rect 25011 24996 25015 25052
rect 24951 24992 25015 24996
rect 25031 25052 25095 25056
rect 25031 24996 25035 25052
rect 25035 24996 25091 25052
rect 25091 24996 25095 25052
rect 25031 24992 25095 24996
rect 7368 24508 7432 24512
rect 7368 24452 7372 24508
rect 7372 24452 7428 24508
rect 7428 24452 7432 24508
rect 7368 24448 7432 24452
rect 7448 24508 7512 24512
rect 7448 24452 7452 24508
rect 7452 24452 7508 24508
rect 7508 24452 7512 24508
rect 7448 24448 7512 24452
rect 7528 24508 7592 24512
rect 7528 24452 7532 24508
rect 7532 24452 7588 24508
rect 7588 24452 7592 24508
rect 7528 24448 7592 24452
rect 7608 24508 7672 24512
rect 7608 24452 7612 24508
rect 7612 24452 7668 24508
rect 7668 24452 7672 24508
rect 7608 24448 7672 24452
rect 14337 24508 14401 24512
rect 14337 24452 14341 24508
rect 14341 24452 14397 24508
rect 14397 24452 14401 24508
rect 14337 24448 14401 24452
rect 14417 24508 14481 24512
rect 14417 24452 14421 24508
rect 14421 24452 14477 24508
rect 14477 24452 14481 24508
rect 14417 24448 14481 24452
rect 14497 24508 14561 24512
rect 14497 24452 14501 24508
rect 14501 24452 14557 24508
rect 14557 24452 14561 24508
rect 14497 24448 14561 24452
rect 14577 24508 14641 24512
rect 14577 24452 14581 24508
rect 14581 24452 14637 24508
rect 14637 24452 14641 24508
rect 14577 24448 14641 24452
rect 21306 24508 21370 24512
rect 21306 24452 21310 24508
rect 21310 24452 21366 24508
rect 21366 24452 21370 24508
rect 21306 24448 21370 24452
rect 21386 24508 21450 24512
rect 21386 24452 21390 24508
rect 21390 24452 21446 24508
rect 21446 24452 21450 24508
rect 21386 24448 21450 24452
rect 21466 24508 21530 24512
rect 21466 24452 21470 24508
rect 21470 24452 21526 24508
rect 21526 24452 21530 24508
rect 21466 24448 21530 24452
rect 21546 24508 21610 24512
rect 21546 24452 21550 24508
rect 21550 24452 21606 24508
rect 21606 24452 21610 24508
rect 21546 24448 21610 24452
rect 28275 24508 28339 24512
rect 28275 24452 28279 24508
rect 28279 24452 28335 24508
rect 28335 24452 28339 24508
rect 28275 24448 28339 24452
rect 28355 24508 28419 24512
rect 28355 24452 28359 24508
rect 28359 24452 28415 24508
rect 28415 24452 28419 24508
rect 28355 24448 28419 24452
rect 28435 24508 28499 24512
rect 28435 24452 28439 24508
rect 28439 24452 28495 24508
rect 28495 24452 28499 24508
rect 28435 24448 28499 24452
rect 28515 24508 28579 24512
rect 28515 24452 28519 24508
rect 28519 24452 28575 24508
rect 28575 24452 28579 24508
rect 28515 24448 28579 24452
rect 3884 23964 3948 23968
rect 3884 23908 3888 23964
rect 3888 23908 3944 23964
rect 3944 23908 3948 23964
rect 3884 23904 3948 23908
rect 3964 23964 4028 23968
rect 3964 23908 3968 23964
rect 3968 23908 4024 23964
rect 4024 23908 4028 23964
rect 3964 23904 4028 23908
rect 4044 23964 4108 23968
rect 4044 23908 4048 23964
rect 4048 23908 4104 23964
rect 4104 23908 4108 23964
rect 4044 23904 4108 23908
rect 4124 23964 4188 23968
rect 4124 23908 4128 23964
rect 4128 23908 4184 23964
rect 4184 23908 4188 23964
rect 4124 23904 4188 23908
rect 10853 23964 10917 23968
rect 10853 23908 10857 23964
rect 10857 23908 10913 23964
rect 10913 23908 10917 23964
rect 10853 23904 10917 23908
rect 10933 23964 10997 23968
rect 10933 23908 10937 23964
rect 10937 23908 10993 23964
rect 10993 23908 10997 23964
rect 10933 23904 10997 23908
rect 11013 23964 11077 23968
rect 11013 23908 11017 23964
rect 11017 23908 11073 23964
rect 11073 23908 11077 23964
rect 11013 23904 11077 23908
rect 11093 23964 11157 23968
rect 11093 23908 11097 23964
rect 11097 23908 11153 23964
rect 11153 23908 11157 23964
rect 11093 23904 11157 23908
rect 17822 23964 17886 23968
rect 17822 23908 17826 23964
rect 17826 23908 17882 23964
rect 17882 23908 17886 23964
rect 17822 23904 17886 23908
rect 17902 23964 17966 23968
rect 17902 23908 17906 23964
rect 17906 23908 17962 23964
rect 17962 23908 17966 23964
rect 17902 23904 17966 23908
rect 17982 23964 18046 23968
rect 17982 23908 17986 23964
rect 17986 23908 18042 23964
rect 18042 23908 18046 23964
rect 17982 23904 18046 23908
rect 18062 23964 18126 23968
rect 18062 23908 18066 23964
rect 18066 23908 18122 23964
rect 18122 23908 18126 23964
rect 18062 23904 18126 23908
rect 24791 23964 24855 23968
rect 24791 23908 24795 23964
rect 24795 23908 24851 23964
rect 24851 23908 24855 23964
rect 24791 23904 24855 23908
rect 24871 23964 24935 23968
rect 24871 23908 24875 23964
rect 24875 23908 24931 23964
rect 24931 23908 24935 23964
rect 24871 23904 24935 23908
rect 24951 23964 25015 23968
rect 24951 23908 24955 23964
rect 24955 23908 25011 23964
rect 25011 23908 25015 23964
rect 24951 23904 25015 23908
rect 25031 23964 25095 23968
rect 25031 23908 25035 23964
rect 25035 23908 25091 23964
rect 25091 23908 25095 23964
rect 25031 23904 25095 23908
rect 7368 23420 7432 23424
rect 7368 23364 7372 23420
rect 7372 23364 7428 23420
rect 7428 23364 7432 23420
rect 7368 23360 7432 23364
rect 7448 23420 7512 23424
rect 7448 23364 7452 23420
rect 7452 23364 7508 23420
rect 7508 23364 7512 23420
rect 7448 23360 7512 23364
rect 7528 23420 7592 23424
rect 7528 23364 7532 23420
rect 7532 23364 7588 23420
rect 7588 23364 7592 23420
rect 7528 23360 7592 23364
rect 7608 23420 7672 23424
rect 7608 23364 7612 23420
rect 7612 23364 7668 23420
rect 7668 23364 7672 23420
rect 7608 23360 7672 23364
rect 14337 23420 14401 23424
rect 14337 23364 14341 23420
rect 14341 23364 14397 23420
rect 14397 23364 14401 23420
rect 14337 23360 14401 23364
rect 14417 23420 14481 23424
rect 14417 23364 14421 23420
rect 14421 23364 14477 23420
rect 14477 23364 14481 23420
rect 14417 23360 14481 23364
rect 14497 23420 14561 23424
rect 14497 23364 14501 23420
rect 14501 23364 14557 23420
rect 14557 23364 14561 23420
rect 14497 23360 14561 23364
rect 14577 23420 14641 23424
rect 14577 23364 14581 23420
rect 14581 23364 14637 23420
rect 14637 23364 14641 23420
rect 14577 23360 14641 23364
rect 21306 23420 21370 23424
rect 21306 23364 21310 23420
rect 21310 23364 21366 23420
rect 21366 23364 21370 23420
rect 21306 23360 21370 23364
rect 21386 23420 21450 23424
rect 21386 23364 21390 23420
rect 21390 23364 21446 23420
rect 21446 23364 21450 23420
rect 21386 23360 21450 23364
rect 21466 23420 21530 23424
rect 21466 23364 21470 23420
rect 21470 23364 21526 23420
rect 21526 23364 21530 23420
rect 21466 23360 21530 23364
rect 21546 23420 21610 23424
rect 21546 23364 21550 23420
rect 21550 23364 21606 23420
rect 21606 23364 21610 23420
rect 21546 23360 21610 23364
rect 28275 23420 28339 23424
rect 28275 23364 28279 23420
rect 28279 23364 28335 23420
rect 28335 23364 28339 23420
rect 28275 23360 28339 23364
rect 28355 23420 28419 23424
rect 28355 23364 28359 23420
rect 28359 23364 28415 23420
rect 28415 23364 28419 23420
rect 28355 23360 28419 23364
rect 28435 23420 28499 23424
rect 28435 23364 28439 23420
rect 28439 23364 28495 23420
rect 28495 23364 28499 23420
rect 28435 23360 28499 23364
rect 28515 23420 28579 23424
rect 28515 23364 28519 23420
rect 28519 23364 28575 23420
rect 28575 23364 28579 23420
rect 28515 23360 28579 23364
rect 3884 22876 3948 22880
rect 3884 22820 3888 22876
rect 3888 22820 3944 22876
rect 3944 22820 3948 22876
rect 3884 22816 3948 22820
rect 3964 22876 4028 22880
rect 3964 22820 3968 22876
rect 3968 22820 4024 22876
rect 4024 22820 4028 22876
rect 3964 22816 4028 22820
rect 4044 22876 4108 22880
rect 4044 22820 4048 22876
rect 4048 22820 4104 22876
rect 4104 22820 4108 22876
rect 4044 22816 4108 22820
rect 4124 22876 4188 22880
rect 4124 22820 4128 22876
rect 4128 22820 4184 22876
rect 4184 22820 4188 22876
rect 4124 22816 4188 22820
rect 10853 22876 10917 22880
rect 10853 22820 10857 22876
rect 10857 22820 10913 22876
rect 10913 22820 10917 22876
rect 10853 22816 10917 22820
rect 10933 22876 10997 22880
rect 10933 22820 10937 22876
rect 10937 22820 10993 22876
rect 10993 22820 10997 22876
rect 10933 22816 10997 22820
rect 11013 22876 11077 22880
rect 11013 22820 11017 22876
rect 11017 22820 11073 22876
rect 11073 22820 11077 22876
rect 11013 22816 11077 22820
rect 11093 22876 11157 22880
rect 11093 22820 11097 22876
rect 11097 22820 11153 22876
rect 11153 22820 11157 22876
rect 11093 22816 11157 22820
rect 17822 22876 17886 22880
rect 17822 22820 17826 22876
rect 17826 22820 17882 22876
rect 17882 22820 17886 22876
rect 17822 22816 17886 22820
rect 17902 22876 17966 22880
rect 17902 22820 17906 22876
rect 17906 22820 17962 22876
rect 17962 22820 17966 22876
rect 17902 22816 17966 22820
rect 17982 22876 18046 22880
rect 17982 22820 17986 22876
rect 17986 22820 18042 22876
rect 18042 22820 18046 22876
rect 17982 22816 18046 22820
rect 18062 22876 18126 22880
rect 18062 22820 18066 22876
rect 18066 22820 18122 22876
rect 18122 22820 18126 22876
rect 18062 22816 18126 22820
rect 24791 22876 24855 22880
rect 24791 22820 24795 22876
rect 24795 22820 24851 22876
rect 24851 22820 24855 22876
rect 24791 22816 24855 22820
rect 24871 22876 24935 22880
rect 24871 22820 24875 22876
rect 24875 22820 24931 22876
rect 24931 22820 24935 22876
rect 24871 22816 24935 22820
rect 24951 22876 25015 22880
rect 24951 22820 24955 22876
rect 24955 22820 25011 22876
rect 25011 22820 25015 22876
rect 24951 22816 25015 22820
rect 25031 22876 25095 22880
rect 25031 22820 25035 22876
rect 25035 22820 25091 22876
rect 25091 22820 25095 22876
rect 25031 22816 25095 22820
rect 7368 22332 7432 22336
rect 7368 22276 7372 22332
rect 7372 22276 7428 22332
rect 7428 22276 7432 22332
rect 7368 22272 7432 22276
rect 7448 22332 7512 22336
rect 7448 22276 7452 22332
rect 7452 22276 7508 22332
rect 7508 22276 7512 22332
rect 7448 22272 7512 22276
rect 7528 22332 7592 22336
rect 7528 22276 7532 22332
rect 7532 22276 7588 22332
rect 7588 22276 7592 22332
rect 7528 22272 7592 22276
rect 7608 22332 7672 22336
rect 7608 22276 7612 22332
rect 7612 22276 7668 22332
rect 7668 22276 7672 22332
rect 7608 22272 7672 22276
rect 14337 22332 14401 22336
rect 14337 22276 14341 22332
rect 14341 22276 14397 22332
rect 14397 22276 14401 22332
rect 14337 22272 14401 22276
rect 14417 22332 14481 22336
rect 14417 22276 14421 22332
rect 14421 22276 14477 22332
rect 14477 22276 14481 22332
rect 14417 22272 14481 22276
rect 14497 22332 14561 22336
rect 14497 22276 14501 22332
rect 14501 22276 14557 22332
rect 14557 22276 14561 22332
rect 14497 22272 14561 22276
rect 14577 22332 14641 22336
rect 14577 22276 14581 22332
rect 14581 22276 14637 22332
rect 14637 22276 14641 22332
rect 14577 22272 14641 22276
rect 21306 22332 21370 22336
rect 21306 22276 21310 22332
rect 21310 22276 21366 22332
rect 21366 22276 21370 22332
rect 21306 22272 21370 22276
rect 21386 22332 21450 22336
rect 21386 22276 21390 22332
rect 21390 22276 21446 22332
rect 21446 22276 21450 22332
rect 21386 22272 21450 22276
rect 21466 22332 21530 22336
rect 21466 22276 21470 22332
rect 21470 22276 21526 22332
rect 21526 22276 21530 22332
rect 21466 22272 21530 22276
rect 21546 22332 21610 22336
rect 21546 22276 21550 22332
rect 21550 22276 21606 22332
rect 21606 22276 21610 22332
rect 21546 22272 21610 22276
rect 28275 22332 28339 22336
rect 28275 22276 28279 22332
rect 28279 22276 28335 22332
rect 28335 22276 28339 22332
rect 28275 22272 28339 22276
rect 28355 22332 28419 22336
rect 28355 22276 28359 22332
rect 28359 22276 28415 22332
rect 28415 22276 28419 22332
rect 28355 22272 28419 22276
rect 28435 22332 28499 22336
rect 28435 22276 28439 22332
rect 28439 22276 28495 22332
rect 28495 22276 28499 22332
rect 28435 22272 28499 22276
rect 28515 22332 28579 22336
rect 28515 22276 28519 22332
rect 28519 22276 28575 22332
rect 28575 22276 28579 22332
rect 28515 22272 28579 22276
rect 3884 21788 3948 21792
rect 3884 21732 3888 21788
rect 3888 21732 3944 21788
rect 3944 21732 3948 21788
rect 3884 21728 3948 21732
rect 3964 21788 4028 21792
rect 3964 21732 3968 21788
rect 3968 21732 4024 21788
rect 4024 21732 4028 21788
rect 3964 21728 4028 21732
rect 4044 21788 4108 21792
rect 4044 21732 4048 21788
rect 4048 21732 4104 21788
rect 4104 21732 4108 21788
rect 4044 21728 4108 21732
rect 4124 21788 4188 21792
rect 4124 21732 4128 21788
rect 4128 21732 4184 21788
rect 4184 21732 4188 21788
rect 4124 21728 4188 21732
rect 10853 21788 10917 21792
rect 10853 21732 10857 21788
rect 10857 21732 10913 21788
rect 10913 21732 10917 21788
rect 10853 21728 10917 21732
rect 10933 21788 10997 21792
rect 10933 21732 10937 21788
rect 10937 21732 10993 21788
rect 10993 21732 10997 21788
rect 10933 21728 10997 21732
rect 11013 21788 11077 21792
rect 11013 21732 11017 21788
rect 11017 21732 11073 21788
rect 11073 21732 11077 21788
rect 11013 21728 11077 21732
rect 11093 21788 11157 21792
rect 11093 21732 11097 21788
rect 11097 21732 11153 21788
rect 11153 21732 11157 21788
rect 11093 21728 11157 21732
rect 17822 21788 17886 21792
rect 17822 21732 17826 21788
rect 17826 21732 17882 21788
rect 17882 21732 17886 21788
rect 17822 21728 17886 21732
rect 17902 21788 17966 21792
rect 17902 21732 17906 21788
rect 17906 21732 17962 21788
rect 17962 21732 17966 21788
rect 17902 21728 17966 21732
rect 17982 21788 18046 21792
rect 17982 21732 17986 21788
rect 17986 21732 18042 21788
rect 18042 21732 18046 21788
rect 17982 21728 18046 21732
rect 18062 21788 18126 21792
rect 18062 21732 18066 21788
rect 18066 21732 18122 21788
rect 18122 21732 18126 21788
rect 18062 21728 18126 21732
rect 24791 21788 24855 21792
rect 24791 21732 24795 21788
rect 24795 21732 24851 21788
rect 24851 21732 24855 21788
rect 24791 21728 24855 21732
rect 24871 21788 24935 21792
rect 24871 21732 24875 21788
rect 24875 21732 24931 21788
rect 24931 21732 24935 21788
rect 24871 21728 24935 21732
rect 24951 21788 25015 21792
rect 24951 21732 24955 21788
rect 24955 21732 25011 21788
rect 25011 21732 25015 21788
rect 24951 21728 25015 21732
rect 25031 21788 25095 21792
rect 25031 21732 25035 21788
rect 25035 21732 25091 21788
rect 25091 21732 25095 21788
rect 25031 21728 25095 21732
rect 7368 21244 7432 21248
rect 7368 21188 7372 21244
rect 7372 21188 7428 21244
rect 7428 21188 7432 21244
rect 7368 21184 7432 21188
rect 7448 21244 7512 21248
rect 7448 21188 7452 21244
rect 7452 21188 7508 21244
rect 7508 21188 7512 21244
rect 7448 21184 7512 21188
rect 7528 21244 7592 21248
rect 7528 21188 7532 21244
rect 7532 21188 7588 21244
rect 7588 21188 7592 21244
rect 7528 21184 7592 21188
rect 7608 21244 7672 21248
rect 7608 21188 7612 21244
rect 7612 21188 7668 21244
rect 7668 21188 7672 21244
rect 7608 21184 7672 21188
rect 14337 21244 14401 21248
rect 14337 21188 14341 21244
rect 14341 21188 14397 21244
rect 14397 21188 14401 21244
rect 14337 21184 14401 21188
rect 14417 21244 14481 21248
rect 14417 21188 14421 21244
rect 14421 21188 14477 21244
rect 14477 21188 14481 21244
rect 14417 21184 14481 21188
rect 14497 21244 14561 21248
rect 14497 21188 14501 21244
rect 14501 21188 14557 21244
rect 14557 21188 14561 21244
rect 14497 21184 14561 21188
rect 14577 21244 14641 21248
rect 14577 21188 14581 21244
rect 14581 21188 14637 21244
rect 14637 21188 14641 21244
rect 14577 21184 14641 21188
rect 21306 21244 21370 21248
rect 21306 21188 21310 21244
rect 21310 21188 21366 21244
rect 21366 21188 21370 21244
rect 21306 21184 21370 21188
rect 21386 21244 21450 21248
rect 21386 21188 21390 21244
rect 21390 21188 21446 21244
rect 21446 21188 21450 21244
rect 21386 21184 21450 21188
rect 21466 21244 21530 21248
rect 21466 21188 21470 21244
rect 21470 21188 21526 21244
rect 21526 21188 21530 21244
rect 21466 21184 21530 21188
rect 21546 21244 21610 21248
rect 21546 21188 21550 21244
rect 21550 21188 21606 21244
rect 21606 21188 21610 21244
rect 21546 21184 21610 21188
rect 28275 21244 28339 21248
rect 28275 21188 28279 21244
rect 28279 21188 28335 21244
rect 28335 21188 28339 21244
rect 28275 21184 28339 21188
rect 28355 21244 28419 21248
rect 28355 21188 28359 21244
rect 28359 21188 28415 21244
rect 28415 21188 28419 21244
rect 28355 21184 28419 21188
rect 28435 21244 28499 21248
rect 28435 21188 28439 21244
rect 28439 21188 28495 21244
rect 28495 21188 28499 21244
rect 28435 21184 28499 21188
rect 28515 21244 28579 21248
rect 28515 21188 28519 21244
rect 28519 21188 28575 21244
rect 28575 21188 28579 21244
rect 28515 21184 28579 21188
rect 13492 20708 13556 20772
rect 3884 20700 3948 20704
rect 3884 20644 3888 20700
rect 3888 20644 3944 20700
rect 3944 20644 3948 20700
rect 3884 20640 3948 20644
rect 3964 20700 4028 20704
rect 3964 20644 3968 20700
rect 3968 20644 4024 20700
rect 4024 20644 4028 20700
rect 3964 20640 4028 20644
rect 4044 20700 4108 20704
rect 4044 20644 4048 20700
rect 4048 20644 4104 20700
rect 4104 20644 4108 20700
rect 4044 20640 4108 20644
rect 4124 20700 4188 20704
rect 4124 20644 4128 20700
rect 4128 20644 4184 20700
rect 4184 20644 4188 20700
rect 4124 20640 4188 20644
rect 10853 20700 10917 20704
rect 10853 20644 10857 20700
rect 10857 20644 10913 20700
rect 10913 20644 10917 20700
rect 10853 20640 10917 20644
rect 10933 20700 10997 20704
rect 10933 20644 10937 20700
rect 10937 20644 10993 20700
rect 10993 20644 10997 20700
rect 10933 20640 10997 20644
rect 11013 20700 11077 20704
rect 11013 20644 11017 20700
rect 11017 20644 11073 20700
rect 11073 20644 11077 20700
rect 11013 20640 11077 20644
rect 11093 20700 11157 20704
rect 11093 20644 11097 20700
rect 11097 20644 11153 20700
rect 11153 20644 11157 20700
rect 11093 20640 11157 20644
rect 17822 20700 17886 20704
rect 17822 20644 17826 20700
rect 17826 20644 17882 20700
rect 17882 20644 17886 20700
rect 17822 20640 17886 20644
rect 17902 20700 17966 20704
rect 17902 20644 17906 20700
rect 17906 20644 17962 20700
rect 17962 20644 17966 20700
rect 17902 20640 17966 20644
rect 17982 20700 18046 20704
rect 17982 20644 17986 20700
rect 17986 20644 18042 20700
rect 18042 20644 18046 20700
rect 17982 20640 18046 20644
rect 18062 20700 18126 20704
rect 18062 20644 18066 20700
rect 18066 20644 18122 20700
rect 18122 20644 18126 20700
rect 18062 20640 18126 20644
rect 24791 20700 24855 20704
rect 24791 20644 24795 20700
rect 24795 20644 24851 20700
rect 24851 20644 24855 20700
rect 24791 20640 24855 20644
rect 24871 20700 24935 20704
rect 24871 20644 24875 20700
rect 24875 20644 24931 20700
rect 24931 20644 24935 20700
rect 24871 20640 24935 20644
rect 24951 20700 25015 20704
rect 24951 20644 24955 20700
rect 24955 20644 25011 20700
rect 25011 20644 25015 20700
rect 24951 20640 25015 20644
rect 25031 20700 25095 20704
rect 25031 20644 25035 20700
rect 25035 20644 25091 20700
rect 25091 20644 25095 20700
rect 25031 20640 25095 20644
rect 7368 20156 7432 20160
rect 7368 20100 7372 20156
rect 7372 20100 7428 20156
rect 7428 20100 7432 20156
rect 7368 20096 7432 20100
rect 7448 20156 7512 20160
rect 7448 20100 7452 20156
rect 7452 20100 7508 20156
rect 7508 20100 7512 20156
rect 7448 20096 7512 20100
rect 7528 20156 7592 20160
rect 7528 20100 7532 20156
rect 7532 20100 7588 20156
rect 7588 20100 7592 20156
rect 7528 20096 7592 20100
rect 7608 20156 7672 20160
rect 7608 20100 7612 20156
rect 7612 20100 7668 20156
rect 7668 20100 7672 20156
rect 7608 20096 7672 20100
rect 14337 20156 14401 20160
rect 14337 20100 14341 20156
rect 14341 20100 14397 20156
rect 14397 20100 14401 20156
rect 14337 20096 14401 20100
rect 14417 20156 14481 20160
rect 14417 20100 14421 20156
rect 14421 20100 14477 20156
rect 14477 20100 14481 20156
rect 14417 20096 14481 20100
rect 14497 20156 14561 20160
rect 14497 20100 14501 20156
rect 14501 20100 14557 20156
rect 14557 20100 14561 20156
rect 14497 20096 14561 20100
rect 14577 20156 14641 20160
rect 14577 20100 14581 20156
rect 14581 20100 14637 20156
rect 14637 20100 14641 20156
rect 14577 20096 14641 20100
rect 21306 20156 21370 20160
rect 21306 20100 21310 20156
rect 21310 20100 21366 20156
rect 21366 20100 21370 20156
rect 21306 20096 21370 20100
rect 21386 20156 21450 20160
rect 21386 20100 21390 20156
rect 21390 20100 21446 20156
rect 21446 20100 21450 20156
rect 21386 20096 21450 20100
rect 21466 20156 21530 20160
rect 21466 20100 21470 20156
rect 21470 20100 21526 20156
rect 21526 20100 21530 20156
rect 21466 20096 21530 20100
rect 21546 20156 21610 20160
rect 21546 20100 21550 20156
rect 21550 20100 21606 20156
rect 21606 20100 21610 20156
rect 21546 20096 21610 20100
rect 28275 20156 28339 20160
rect 28275 20100 28279 20156
rect 28279 20100 28335 20156
rect 28335 20100 28339 20156
rect 28275 20096 28339 20100
rect 28355 20156 28419 20160
rect 28355 20100 28359 20156
rect 28359 20100 28415 20156
rect 28415 20100 28419 20156
rect 28355 20096 28419 20100
rect 28435 20156 28499 20160
rect 28435 20100 28439 20156
rect 28439 20100 28495 20156
rect 28495 20100 28499 20156
rect 28435 20096 28499 20100
rect 28515 20156 28579 20160
rect 28515 20100 28519 20156
rect 28519 20100 28575 20156
rect 28575 20100 28579 20156
rect 28515 20096 28579 20100
rect 3884 19612 3948 19616
rect 3884 19556 3888 19612
rect 3888 19556 3944 19612
rect 3944 19556 3948 19612
rect 3884 19552 3948 19556
rect 3964 19612 4028 19616
rect 3964 19556 3968 19612
rect 3968 19556 4024 19612
rect 4024 19556 4028 19612
rect 3964 19552 4028 19556
rect 4044 19612 4108 19616
rect 4044 19556 4048 19612
rect 4048 19556 4104 19612
rect 4104 19556 4108 19612
rect 4044 19552 4108 19556
rect 4124 19612 4188 19616
rect 4124 19556 4128 19612
rect 4128 19556 4184 19612
rect 4184 19556 4188 19612
rect 4124 19552 4188 19556
rect 10853 19612 10917 19616
rect 10853 19556 10857 19612
rect 10857 19556 10913 19612
rect 10913 19556 10917 19612
rect 10853 19552 10917 19556
rect 10933 19612 10997 19616
rect 10933 19556 10937 19612
rect 10937 19556 10993 19612
rect 10993 19556 10997 19612
rect 10933 19552 10997 19556
rect 11013 19612 11077 19616
rect 11013 19556 11017 19612
rect 11017 19556 11073 19612
rect 11073 19556 11077 19612
rect 11013 19552 11077 19556
rect 11093 19612 11157 19616
rect 11093 19556 11097 19612
rect 11097 19556 11153 19612
rect 11153 19556 11157 19612
rect 11093 19552 11157 19556
rect 17822 19612 17886 19616
rect 17822 19556 17826 19612
rect 17826 19556 17882 19612
rect 17882 19556 17886 19612
rect 17822 19552 17886 19556
rect 17902 19612 17966 19616
rect 17902 19556 17906 19612
rect 17906 19556 17962 19612
rect 17962 19556 17966 19612
rect 17902 19552 17966 19556
rect 17982 19612 18046 19616
rect 17982 19556 17986 19612
rect 17986 19556 18042 19612
rect 18042 19556 18046 19612
rect 17982 19552 18046 19556
rect 18062 19612 18126 19616
rect 18062 19556 18066 19612
rect 18066 19556 18122 19612
rect 18122 19556 18126 19612
rect 18062 19552 18126 19556
rect 24791 19612 24855 19616
rect 24791 19556 24795 19612
rect 24795 19556 24851 19612
rect 24851 19556 24855 19612
rect 24791 19552 24855 19556
rect 24871 19612 24935 19616
rect 24871 19556 24875 19612
rect 24875 19556 24931 19612
rect 24931 19556 24935 19612
rect 24871 19552 24935 19556
rect 24951 19612 25015 19616
rect 24951 19556 24955 19612
rect 24955 19556 25011 19612
rect 25011 19556 25015 19612
rect 24951 19552 25015 19556
rect 25031 19612 25095 19616
rect 25031 19556 25035 19612
rect 25035 19556 25091 19612
rect 25091 19556 25095 19612
rect 25031 19552 25095 19556
rect 7368 19068 7432 19072
rect 7368 19012 7372 19068
rect 7372 19012 7428 19068
rect 7428 19012 7432 19068
rect 7368 19008 7432 19012
rect 7448 19068 7512 19072
rect 7448 19012 7452 19068
rect 7452 19012 7508 19068
rect 7508 19012 7512 19068
rect 7448 19008 7512 19012
rect 7528 19068 7592 19072
rect 7528 19012 7532 19068
rect 7532 19012 7588 19068
rect 7588 19012 7592 19068
rect 7528 19008 7592 19012
rect 7608 19068 7672 19072
rect 7608 19012 7612 19068
rect 7612 19012 7668 19068
rect 7668 19012 7672 19068
rect 7608 19008 7672 19012
rect 14337 19068 14401 19072
rect 14337 19012 14341 19068
rect 14341 19012 14397 19068
rect 14397 19012 14401 19068
rect 14337 19008 14401 19012
rect 14417 19068 14481 19072
rect 14417 19012 14421 19068
rect 14421 19012 14477 19068
rect 14477 19012 14481 19068
rect 14417 19008 14481 19012
rect 14497 19068 14561 19072
rect 14497 19012 14501 19068
rect 14501 19012 14557 19068
rect 14557 19012 14561 19068
rect 14497 19008 14561 19012
rect 14577 19068 14641 19072
rect 14577 19012 14581 19068
rect 14581 19012 14637 19068
rect 14637 19012 14641 19068
rect 14577 19008 14641 19012
rect 21306 19068 21370 19072
rect 21306 19012 21310 19068
rect 21310 19012 21366 19068
rect 21366 19012 21370 19068
rect 21306 19008 21370 19012
rect 21386 19068 21450 19072
rect 21386 19012 21390 19068
rect 21390 19012 21446 19068
rect 21446 19012 21450 19068
rect 21386 19008 21450 19012
rect 21466 19068 21530 19072
rect 21466 19012 21470 19068
rect 21470 19012 21526 19068
rect 21526 19012 21530 19068
rect 21466 19008 21530 19012
rect 21546 19068 21610 19072
rect 21546 19012 21550 19068
rect 21550 19012 21606 19068
rect 21606 19012 21610 19068
rect 21546 19008 21610 19012
rect 28275 19068 28339 19072
rect 28275 19012 28279 19068
rect 28279 19012 28335 19068
rect 28335 19012 28339 19068
rect 28275 19008 28339 19012
rect 28355 19068 28419 19072
rect 28355 19012 28359 19068
rect 28359 19012 28415 19068
rect 28415 19012 28419 19068
rect 28355 19008 28419 19012
rect 28435 19068 28499 19072
rect 28435 19012 28439 19068
rect 28439 19012 28495 19068
rect 28495 19012 28499 19068
rect 28435 19008 28499 19012
rect 28515 19068 28579 19072
rect 28515 19012 28519 19068
rect 28519 19012 28575 19068
rect 28575 19012 28579 19068
rect 28515 19008 28579 19012
rect 3884 18524 3948 18528
rect 3884 18468 3888 18524
rect 3888 18468 3944 18524
rect 3944 18468 3948 18524
rect 3884 18464 3948 18468
rect 3964 18524 4028 18528
rect 3964 18468 3968 18524
rect 3968 18468 4024 18524
rect 4024 18468 4028 18524
rect 3964 18464 4028 18468
rect 4044 18524 4108 18528
rect 4044 18468 4048 18524
rect 4048 18468 4104 18524
rect 4104 18468 4108 18524
rect 4044 18464 4108 18468
rect 4124 18524 4188 18528
rect 4124 18468 4128 18524
rect 4128 18468 4184 18524
rect 4184 18468 4188 18524
rect 4124 18464 4188 18468
rect 10853 18524 10917 18528
rect 10853 18468 10857 18524
rect 10857 18468 10913 18524
rect 10913 18468 10917 18524
rect 10853 18464 10917 18468
rect 10933 18524 10997 18528
rect 10933 18468 10937 18524
rect 10937 18468 10993 18524
rect 10993 18468 10997 18524
rect 10933 18464 10997 18468
rect 11013 18524 11077 18528
rect 11013 18468 11017 18524
rect 11017 18468 11073 18524
rect 11073 18468 11077 18524
rect 11013 18464 11077 18468
rect 11093 18524 11157 18528
rect 11093 18468 11097 18524
rect 11097 18468 11153 18524
rect 11153 18468 11157 18524
rect 11093 18464 11157 18468
rect 17822 18524 17886 18528
rect 17822 18468 17826 18524
rect 17826 18468 17882 18524
rect 17882 18468 17886 18524
rect 17822 18464 17886 18468
rect 17902 18524 17966 18528
rect 17902 18468 17906 18524
rect 17906 18468 17962 18524
rect 17962 18468 17966 18524
rect 17902 18464 17966 18468
rect 17982 18524 18046 18528
rect 17982 18468 17986 18524
rect 17986 18468 18042 18524
rect 18042 18468 18046 18524
rect 17982 18464 18046 18468
rect 18062 18524 18126 18528
rect 18062 18468 18066 18524
rect 18066 18468 18122 18524
rect 18122 18468 18126 18524
rect 18062 18464 18126 18468
rect 24791 18524 24855 18528
rect 24791 18468 24795 18524
rect 24795 18468 24851 18524
rect 24851 18468 24855 18524
rect 24791 18464 24855 18468
rect 24871 18524 24935 18528
rect 24871 18468 24875 18524
rect 24875 18468 24931 18524
rect 24931 18468 24935 18524
rect 24871 18464 24935 18468
rect 24951 18524 25015 18528
rect 24951 18468 24955 18524
rect 24955 18468 25011 18524
rect 25011 18468 25015 18524
rect 24951 18464 25015 18468
rect 25031 18524 25095 18528
rect 25031 18468 25035 18524
rect 25035 18468 25091 18524
rect 25091 18468 25095 18524
rect 25031 18464 25095 18468
rect 7368 17980 7432 17984
rect 7368 17924 7372 17980
rect 7372 17924 7428 17980
rect 7428 17924 7432 17980
rect 7368 17920 7432 17924
rect 7448 17980 7512 17984
rect 7448 17924 7452 17980
rect 7452 17924 7508 17980
rect 7508 17924 7512 17980
rect 7448 17920 7512 17924
rect 7528 17980 7592 17984
rect 7528 17924 7532 17980
rect 7532 17924 7588 17980
rect 7588 17924 7592 17980
rect 7528 17920 7592 17924
rect 7608 17980 7672 17984
rect 7608 17924 7612 17980
rect 7612 17924 7668 17980
rect 7668 17924 7672 17980
rect 7608 17920 7672 17924
rect 14337 17980 14401 17984
rect 14337 17924 14341 17980
rect 14341 17924 14397 17980
rect 14397 17924 14401 17980
rect 14337 17920 14401 17924
rect 14417 17980 14481 17984
rect 14417 17924 14421 17980
rect 14421 17924 14477 17980
rect 14477 17924 14481 17980
rect 14417 17920 14481 17924
rect 14497 17980 14561 17984
rect 14497 17924 14501 17980
rect 14501 17924 14557 17980
rect 14557 17924 14561 17980
rect 14497 17920 14561 17924
rect 14577 17980 14641 17984
rect 14577 17924 14581 17980
rect 14581 17924 14637 17980
rect 14637 17924 14641 17980
rect 14577 17920 14641 17924
rect 21306 17980 21370 17984
rect 21306 17924 21310 17980
rect 21310 17924 21366 17980
rect 21366 17924 21370 17980
rect 21306 17920 21370 17924
rect 21386 17980 21450 17984
rect 21386 17924 21390 17980
rect 21390 17924 21446 17980
rect 21446 17924 21450 17980
rect 21386 17920 21450 17924
rect 21466 17980 21530 17984
rect 21466 17924 21470 17980
rect 21470 17924 21526 17980
rect 21526 17924 21530 17980
rect 21466 17920 21530 17924
rect 21546 17980 21610 17984
rect 21546 17924 21550 17980
rect 21550 17924 21606 17980
rect 21606 17924 21610 17980
rect 21546 17920 21610 17924
rect 28275 17980 28339 17984
rect 28275 17924 28279 17980
rect 28279 17924 28335 17980
rect 28335 17924 28339 17980
rect 28275 17920 28339 17924
rect 28355 17980 28419 17984
rect 28355 17924 28359 17980
rect 28359 17924 28415 17980
rect 28415 17924 28419 17980
rect 28355 17920 28419 17924
rect 28435 17980 28499 17984
rect 28435 17924 28439 17980
rect 28439 17924 28495 17980
rect 28495 17924 28499 17980
rect 28435 17920 28499 17924
rect 28515 17980 28579 17984
rect 28515 17924 28519 17980
rect 28519 17924 28575 17980
rect 28575 17924 28579 17980
rect 28515 17920 28579 17924
rect 3884 17436 3948 17440
rect 3884 17380 3888 17436
rect 3888 17380 3944 17436
rect 3944 17380 3948 17436
rect 3884 17376 3948 17380
rect 3964 17436 4028 17440
rect 3964 17380 3968 17436
rect 3968 17380 4024 17436
rect 4024 17380 4028 17436
rect 3964 17376 4028 17380
rect 4044 17436 4108 17440
rect 4044 17380 4048 17436
rect 4048 17380 4104 17436
rect 4104 17380 4108 17436
rect 4044 17376 4108 17380
rect 4124 17436 4188 17440
rect 4124 17380 4128 17436
rect 4128 17380 4184 17436
rect 4184 17380 4188 17436
rect 4124 17376 4188 17380
rect 10853 17436 10917 17440
rect 10853 17380 10857 17436
rect 10857 17380 10913 17436
rect 10913 17380 10917 17436
rect 10853 17376 10917 17380
rect 10933 17436 10997 17440
rect 10933 17380 10937 17436
rect 10937 17380 10993 17436
rect 10993 17380 10997 17436
rect 10933 17376 10997 17380
rect 11013 17436 11077 17440
rect 11013 17380 11017 17436
rect 11017 17380 11073 17436
rect 11073 17380 11077 17436
rect 11013 17376 11077 17380
rect 11093 17436 11157 17440
rect 11093 17380 11097 17436
rect 11097 17380 11153 17436
rect 11153 17380 11157 17436
rect 11093 17376 11157 17380
rect 17822 17436 17886 17440
rect 17822 17380 17826 17436
rect 17826 17380 17882 17436
rect 17882 17380 17886 17436
rect 17822 17376 17886 17380
rect 17902 17436 17966 17440
rect 17902 17380 17906 17436
rect 17906 17380 17962 17436
rect 17962 17380 17966 17436
rect 17902 17376 17966 17380
rect 17982 17436 18046 17440
rect 17982 17380 17986 17436
rect 17986 17380 18042 17436
rect 18042 17380 18046 17436
rect 17982 17376 18046 17380
rect 18062 17436 18126 17440
rect 18062 17380 18066 17436
rect 18066 17380 18122 17436
rect 18122 17380 18126 17436
rect 18062 17376 18126 17380
rect 24791 17436 24855 17440
rect 24791 17380 24795 17436
rect 24795 17380 24851 17436
rect 24851 17380 24855 17436
rect 24791 17376 24855 17380
rect 24871 17436 24935 17440
rect 24871 17380 24875 17436
rect 24875 17380 24931 17436
rect 24931 17380 24935 17436
rect 24871 17376 24935 17380
rect 24951 17436 25015 17440
rect 24951 17380 24955 17436
rect 24955 17380 25011 17436
rect 25011 17380 25015 17436
rect 24951 17376 25015 17380
rect 25031 17436 25095 17440
rect 25031 17380 25035 17436
rect 25035 17380 25091 17436
rect 25091 17380 25095 17436
rect 25031 17376 25095 17380
rect 7368 16892 7432 16896
rect 7368 16836 7372 16892
rect 7372 16836 7428 16892
rect 7428 16836 7432 16892
rect 7368 16832 7432 16836
rect 7448 16892 7512 16896
rect 7448 16836 7452 16892
rect 7452 16836 7508 16892
rect 7508 16836 7512 16892
rect 7448 16832 7512 16836
rect 7528 16892 7592 16896
rect 7528 16836 7532 16892
rect 7532 16836 7588 16892
rect 7588 16836 7592 16892
rect 7528 16832 7592 16836
rect 7608 16892 7672 16896
rect 7608 16836 7612 16892
rect 7612 16836 7668 16892
rect 7668 16836 7672 16892
rect 7608 16832 7672 16836
rect 14337 16892 14401 16896
rect 14337 16836 14341 16892
rect 14341 16836 14397 16892
rect 14397 16836 14401 16892
rect 14337 16832 14401 16836
rect 14417 16892 14481 16896
rect 14417 16836 14421 16892
rect 14421 16836 14477 16892
rect 14477 16836 14481 16892
rect 14417 16832 14481 16836
rect 14497 16892 14561 16896
rect 14497 16836 14501 16892
rect 14501 16836 14557 16892
rect 14557 16836 14561 16892
rect 14497 16832 14561 16836
rect 14577 16892 14641 16896
rect 14577 16836 14581 16892
rect 14581 16836 14637 16892
rect 14637 16836 14641 16892
rect 14577 16832 14641 16836
rect 21306 16892 21370 16896
rect 21306 16836 21310 16892
rect 21310 16836 21366 16892
rect 21366 16836 21370 16892
rect 21306 16832 21370 16836
rect 21386 16892 21450 16896
rect 21386 16836 21390 16892
rect 21390 16836 21446 16892
rect 21446 16836 21450 16892
rect 21386 16832 21450 16836
rect 21466 16892 21530 16896
rect 21466 16836 21470 16892
rect 21470 16836 21526 16892
rect 21526 16836 21530 16892
rect 21466 16832 21530 16836
rect 21546 16892 21610 16896
rect 21546 16836 21550 16892
rect 21550 16836 21606 16892
rect 21606 16836 21610 16892
rect 21546 16832 21610 16836
rect 28275 16892 28339 16896
rect 28275 16836 28279 16892
rect 28279 16836 28335 16892
rect 28335 16836 28339 16892
rect 28275 16832 28339 16836
rect 28355 16892 28419 16896
rect 28355 16836 28359 16892
rect 28359 16836 28415 16892
rect 28415 16836 28419 16892
rect 28355 16832 28419 16836
rect 28435 16892 28499 16896
rect 28435 16836 28439 16892
rect 28439 16836 28495 16892
rect 28495 16836 28499 16892
rect 28435 16832 28499 16836
rect 28515 16892 28579 16896
rect 28515 16836 28519 16892
rect 28519 16836 28575 16892
rect 28575 16836 28579 16892
rect 28515 16832 28579 16836
rect 13492 16416 13556 16420
rect 13492 16360 13506 16416
rect 13506 16360 13556 16416
rect 13492 16356 13556 16360
rect 3884 16348 3948 16352
rect 3884 16292 3888 16348
rect 3888 16292 3944 16348
rect 3944 16292 3948 16348
rect 3884 16288 3948 16292
rect 3964 16348 4028 16352
rect 3964 16292 3968 16348
rect 3968 16292 4024 16348
rect 4024 16292 4028 16348
rect 3964 16288 4028 16292
rect 4044 16348 4108 16352
rect 4044 16292 4048 16348
rect 4048 16292 4104 16348
rect 4104 16292 4108 16348
rect 4044 16288 4108 16292
rect 4124 16348 4188 16352
rect 4124 16292 4128 16348
rect 4128 16292 4184 16348
rect 4184 16292 4188 16348
rect 4124 16288 4188 16292
rect 10853 16348 10917 16352
rect 10853 16292 10857 16348
rect 10857 16292 10913 16348
rect 10913 16292 10917 16348
rect 10853 16288 10917 16292
rect 10933 16348 10997 16352
rect 10933 16292 10937 16348
rect 10937 16292 10993 16348
rect 10993 16292 10997 16348
rect 10933 16288 10997 16292
rect 11013 16348 11077 16352
rect 11013 16292 11017 16348
rect 11017 16292 11073 16348
rect 11073 16292 11077 16348
rect 11013 16288 11077 16292
rect 11093 16348 11157 16352
rect 11093 16292 11097 16348
rect 11097 16292 11153 16348
rect 11153 16292 11157 16348
rect 11093 16288 11157 16292
rect 17822 16348 17886 16352
rect 17822 16292 17826 16348
rect 17826 16292 17882 16348
rect 17882 16292 17886 16348
rect 17822 16288 17886 16292
rect 17902 16348 17966 16352
rect 17902 16292 17906 16348
rect 17906 16292 17962 16348
rect 17962 16292 17966 16348
rect 17902 16288 17966 16292
rect 17982 16348 18046 16352
rect 17982 16292 17986 16348
rect 17986 16292 18042 16348
rect 18042 16292 18046 16348
rect 17982 16288 18046 16292
rect 18062 16348 18126 16352
rect 18062 16292 18066 16348
rect 18066 16292 18122 16348
rect 18122 16292 18126 16348
rect 18062 16288 18126 16292
rect 24791 16348 24855 16352
rect 24791 16292 24795 16348
rect 24795 16292 24851 16348
rect 24851 16292 24855 16348
rect 24791 16288 24855 16292
rect 24871 16348 24935 16352
rect 24871 16292 24875 16348
rect 24875 16292 24931 16348
rect 24931 16292 24935 16348
rect 24871 16288 24935 16292
rect 24951 16348 25015 16352
rect 24951 16292 24955 16348
rect 24955 16292 25011 16348
rect 25011 16292 25015 16348
rect 24951 16288 25015 16292
rect 25031 16348 25095 16352
rect 25031 16292 25035 16348
rect 25035 16292 25091 16348
rect 25091 16292 25095 16348
rect 25031 16288 25095 16292
rect 7368 15804 7432 15808
rect 7368 15748 7372 15804
rect 7372 15748 7428 15804
rect 7428 15748 7432 15804
rect 7368 15744 7432 15748
rect 7448 15804 7512 15808
rect 7448 15748 7452 15804
rect 7452 15748 7508 15804
rect 7508 15748 7512 15804
rect 7448 15744 7512 15748
rect 7528 15804 7592 15808
rect 7528 15748 7532 15804
rect 7532 15748 7588 15804
rect 7588 15748 7592 15804
rect 7528 15744 7592 15748
rect 7608 15804 7672 15808
rect 7608 15748 7612 15804
rect 7612 15748 7668 15804
rect 7668 15748 7672 15804
rect 7608 15744 7672 15748
rect 14337 15804 14401 15808
rect 14337 15748 14341 15804
rect 14341 15748 14397 15804
rect 14397 15748 14401 15804
rect 14337 15744 14401 15748
rect 14417 15804 14481 15808
rect 14417 15748 14421 15804
rect 14421 15748 14477 15804
rect 14477 15748 14481 15804
rect 14417 15744 14481 15748
rect 14497 15804 14561 15808
rect 14497 15748 14501 15804
rect 14501 15748 14557 15804
rect 14557 15748 14561 15804
rect 14497 15744 14561 15748
rect 14577 15804 14641 15808
rect 14577 15748 14581 15804
rect 14581 15748 14637 15804
rect 14637 15748 14641 15804
rect 14577 15744 14641 15748
rect 21306 15804 21370 15808
rect 21306 15748 21310 15804
rect 21310 15748 21366 15804
rect 21366 15748 21370 15804
rect 21306 15744 21370 15748
rect 21386 15804 21450 15808
rect 21386 15748 21390 15804
rect 21390 15748 21446 15804
rect 21446 15748 21450 15804
rect 21386 15744 21450 15748
rect 21466 15804 21530 15808
rect 21466 15748 21470 15804
rect 21470 15748 21526 15804
rect 21526 15748 21530 15804
rect 21466 15744 21530 15748
rect 21546 15804 21610 15808
rect 21546 15748 21550 15804
rect 21550 15748 21606 15804
rect 21606 15748 21610 15804
rect 21546 15744 21610 15748
rect 28275 15804 28339 15808
rect 28275 15748 28279 15804
rect 28279 15748 28335 15804
rect 28335 15748 28339 15804
rect 28275 15744 28339 15748
rect 28355 15804 28419 15808
rect 28355 15748 28359 15804
rect 28359 15748 28415 15804
rect 28415 15748 28419 15804
rect 28355 15744 28419 15748
rect 28435 15804 28499 15808
rect 28435 15748 28439 15804
rect 28439 15748 28495 15804
rect 28495 15748 28499 15804
rect 28435 15744 28499 15748
rect 28515 15804 28579 15808
rect 28515 15748 28519 15804
rect 28519 15748 28575 15804
rect 28575 15748 28579 15804
rect 28515 15744 28579 15748
rect 3884 15260 3948 15264
rect 3884 15204 3888 15260
rect 3888 15204 3944 15260
rect 3944 15204 3948 15260
rect 3884 15200 3948 15204
rect 3964 15260 4028 15264
rect 3964 15204 3968 15260
rect 3968 15204 4024 15260
rect 4024 15204 4028 15260
rect 3964 15200 4028 15204
rect 4044 15260 4108 15264
rect 4044 15204 4048 15260
rect 4048 15204 4104 15260
rect 4104 15204 4108 15260
rect 4044 15200 4108 15204
rect 4124 15260 4188 15264
rect 4124 15204 4128 15260
rect 4128 15204 4184 15260
rect 4184 15204 4188 15260
rect 4124 15200 4188 15204
rect 10853 15260 10917 15264
rect 10853 15204 10857 15260
rect 10857 15204 10913 15260
rect 10913 15204 10917 15260
rect 10853 15200 10917 15204
rect 10933 15260 10997 15264
rect 10933 15204 10937 15260
rect 10937 15204 10993 15260
rect 10993 15204 10997 15260
rect 10933 15200 10997 15204
rect 11013 15260 11077 15264
rect 11013 15204 11017 15260
rect 11017 15204 11073 15260
rect 11073 15204 11077 15260
rect 11013 15200 11077 15204
rect 11093 15260 11157 15264
rect 11093 15204 11097 15260
rect 11097 15204 11153 15260
rect 11153 15204 11157 15260
rect 11093 15200 11157 15204
rect 17822 15260 17886 15264
rect 17822 15204 17826 15260
rect 17826 15204 17882 15260
rect 17882 15204 17886 15260
rect 17822 15200 17886 15204
rect 17902 15260 17966 15264
rect 17902 15204 17906 15260
rect 17906 15204 17962 15260
rect 17962 15204 17966 15260
rect 17902 15200 17966 15204
rect 17982 15260 18046 15264
rect 17982 15204 17986 15260
rect 17986 15204 18042 15260
rect 18042 15204 18046 15260
rect 17982 15200 18046 15204
rect 18062 15260 18126 15264
rect 18062 15204 18066 15260
rect 18066 15204 18122 15260
rect 18122 15204 18126 15260
rect 18062 15200 18126 15204
rect 24791 15260 24855 15264
rect 24791 15204 24795 15260
rect 24795 15204 24851 15260
rect 24851 15204 24855 15260
rect 24791 15200 24855 15204
rect 24871 15260 24935 15264
rect 24871 15204 24875 15260
rect 24875 15204 24931 15260
rect 24931 15204 24935 15260
rect 24871 15200 24935 15204
rect 24951 15260 25015 15264
rect 24951 15204 24955 15260
rect 24955 15204 25011 15260
rect 25011 15204 25015 15260
rect 24951 15200 25015 15204
rect 25031 15260 25095 15264
rect 25031 15204 25035 15260
rect 25035 15204 25091 15260
rect 25091 15204 25095 15260
rect 25031 15200 25095 15204
rect 7368 14716 7432 14720
rect 7368 14660 7372 14716
rect 7372 14660 7428 14716
rect 7428 14660 7432 14716
rect 7368 14656 7432 14660
rect 7448 14716 7512 14720
rect 7448 14660 7452 14716
rect 7452 14660 7508 14716
rect 7508 14660 7512 14716
rect 7448 14656 7512 14660
rect 7528 14716 7592 14720
rect 7528 14660 7532 14716
rect 7532 14660 7588 14716
rect 7588 14660 7592 14716
rect 7528 14656 7592 14660
rect 7608 14716 7672 14720
rect 7608 14660 7612 14716
rect 7612 14660 7668 14716
rect 7668 14660 7672 14716
rect 7608 14656 7672 14660
rect 14337 14716 14401 14720
rect 14337 14660 14341 14716
rect 14341 14660 14397 14716
rect 14397 14660 14401 14716
rect 14337 14656 14401 14660
rect 14417 14716 14481 14720
rect 14417 14660 14421 14716
rect 14421 14660 14477 14716
rect 14477 14660 14481 14716
rect 14417 14656 14481 14660
rect 14497 14716 14561 14720
rect 14497 14660 14501 14716
rect 14501 14660 14557 14716
rect 14557 14660 14561 14716
rect 14497 14656 14561 14660
rect 14577 14716 14641 14720
rect 14577 14660 14581 14716
rect 14581 14660 14637 14716
rect 14637 14660 14641 14716
rect 14577 14656 14641 14660
rect 21306 14716 21370 14720
rect 21306 14660 21310 14716
rect 21310 14660 21366 14716
rect 21366 14660 21370 14716
rect 21306 14656 21370 14660
rect 21386 14716 21450 14720
rect 21386 14660 21390 14716
rect 21390 14660 21446 14716
rect 21446 14660 21450 14716
rect 21386 14656 21450 14660
rect 21466 14716 21530 14720
rect 21466 14660 21470 14716
rect 21470 14660 21526 14716
rect 21526 14660 21530 14716
rect 21466 14656 21530 14660
rect 21546 14716 21610 14720
rect 21546 14660 21550 14716
rect 21550 14660 21606 14716
rect 21606 14660 21610 14716
rect 21546 14656 21610 14660
rect 28275 14716 28339 14720
rect 28275 14660 28279 14716
rect 28279 14660 28335 14716
rect 28335 14660 28339 14716
rect 28275 14656 28339 14660
rect 28355 14716 28419 14720
rect 28355 14660 28359 14716
rect 28359 14660 28415 14716
rect 28415 14660 28419 14716
rect 28355 14656 28419 14660
rect 28435 14716 28499 14720
rect 28435 14660 28439 14716
rect 28439 14660 28495 14716
rect 28495 14660 28499 14716
rect 28435 14656 28499 14660
rect 28515 14716 28579 14720
rect 28515 14660 28519 14716
rect 28519 14660 28575 14716
rect 28575 14660 28579 14716
rect 28515 14656 28579 14660
rect 3884 14172 3948 14176
rect 3884 14116 3888 14172
rect 3888 14116 3944 14172
rect 3944 14116 3948 14172
rect 3884 14112 3948 14116
rect 3964 14172 4028 14176
rect 3964 14116 3968 14172
rect 3968 14116 4024 14172
rect 4024 14116 4028 14172
rect 3964 14112 4028 14116
rect 4044 14172 4108 14176
rect 4044 14116 4048 14172
rect 4048 14116 4104 14172
rect 4104 14116 4108 14172
rect 4044 14112 4108 14116
rect 4124 14172 4188 14176
rect 4124 14116 4128 14172
rect 4128 14116 4184 14172
rect 4184 14116 4188 14172
rect 4124 14112 4188 14116
rect 10853 14172 10917 14176
rect 10853 14116 10857 14172
rect 10857 14116 10913 14172
rect 10913 14116 10917 14172
rect 10853 14112 10917 14116
rect 10933 14172 10997 14176
rect 10933 14116 10937 14172
rect 10937 14116 10993 14172
rect 10993 14116 10997 14172
rect 10933 14112 10997 14116
rect 11013 14172 11077 14176
rect 11013 14116 11017 14172
rect 11017 14116 11073 14172
rect 11073 14116 11077 14172
rect 11013 14112 11077 14116
rect 11093 14172 11157 14176
rect 11093 14116 11097 14172
rect 11097 14116 11153 14172
rect 11153 14116 11157 14172
rect 11093 14112 11157 14116
rect 17822 14172 17886 14176
rect 17822 14116 17826 14172
rect 17826 14116 17882 14172
rect 17882 14116 17886 14172
rect 17822 14112 17886 14116
rect 17902 14172 17966 14176
rect 17902 14116 17906 14172
rect 17906 14116 17962 14172
rect 17962 14116 17966 14172
rect 17902 14112 17966 14116
rect 17982 14172 18046 14176
rect 17982 14116 17986 14172
rect 17986 14116 18042 14172
rect 18042 14116 18046 14172
rect 17982 14112 18046 14116
rect 18062 14172 18126 14176
rect 18062 14116 18066 14172
rect 18066 14116 18122 14172
rect 18122 14116 18126 14172
rect 18062 14112 18126 14116
rect 24791 14172 24855 14176
rect 24791 14116 24795 14172
rect 24795 14116 24851 14172
rect 24851 14116 24855 14172
rect 24791 14112 24855 14116
rect 24871 14172 24935 14176
rect 24871 14116 24875 14172
rect 24875 14116 24931 14172
rect 24931 14116 24935 14172
rect 24871 14112 24935 14116
rect 24951 14172 25015 14176
rect 24951 14116 24955 14172
rect 24955 14116 25011 14172
rect 25011 14116 25015 14172
rect 24951 14112 25015 14116
rect 25031 14172 25095 14176
rect 25031 14116 25035 14172
rect 25035 14116 25091 14172
rect 25091 14116 25095 14172
rect 25031 14112 25095 14116
rect 7368 13628 7432 13632
rect 7368 13572 7372 13628
rect 7372 13572 7428 13628
rect 7428 13572 7432 13628
rect 7368 13568 7432 13572
rect 7448 13628 7512 13632
rect 7448 13572 7452 13628
rect 7452 13572 7508 13628
rect 7508 13572 7512 13628
rect 7448 13568 7512 13572
rect 7528 13628 7592 13632
rect 7528 13572 7532 13628
rect 7532 13572 7588 13628
rect 7588 13572 7592 13628
rect 7528 13568 7592 13572
rect 7608 13628 7672 13632
rect 7608 13572 7612 13628
rect 7612 13572 7668 13628
rect 7668 13572 7672 13628
rect 7608 13568 7672 13572
rect 14337 13628 14401 13632
rect 14337 13572 14341 13628
rect 14341 13572 14397 13628
rect 14397 13572 14401 13628
rect 14337 13568 14401 13572
rect 14417 13628 14481 13632
rect 14417 13572 14421 13628
rect 14421 13572 14477 13628
rect 14477 13572 14481 13628
rect 14417 13568 14481 13572
rect 14497 13628 14561 13632
rect 14497 13572 14501 13628
rect 14501 13572 14557 13628
rect 14557 13572 14561 13628
rect 14497 13568 14561 13572
rect 14577 13628 14641 13632
rect 14577 13572 14581 13628
rect 14581 13572 14637 13628
rect 14637 13572 14641 13628
rect 14577 13568 14641 13572
rect 21306 13628 21370 13632
rect 21306 13572 21310 13628
rect 21310 13572 21366 13628
rect 21366 13572 21370 13628
rect 21306 13568 21370 13572
rect 21386 13628 21450 13632
rect 21386 13572 21390 13628
rect 21390 13572 21446 13628
rect 21446 13572 21450 13628
rect 21386 13568 21450 13572
rect 21466 13628 21530 13632
rect 21466 13572 21470 13628
rect 21470 13572 21526 13628
rect 21526 13572 21530 13628
rect 21466 13568 21530 13572
rect 21546 13628 21610 13632
rect 21546 13572 21550 13628
rect 21550 13572 21606 13628
rect 21606 13572 21610 13628
rect 21546 13568 21610 13572
rect 28275 13628 28339 13632
rect 28275 13572 28279 13628
rect 28279 13572 28335 13628
rect 28335 13572 28339 13628
rect 28275 13568 28339 13572
rect 28355 13628 28419 13632
rect 28355 13572 28359 13628
rect 28359 13572 28415 13628
rect 28415 13572 28419 13628
rect 28355 13568 28419 13572
rect 28435 13628 28499 13632
rect 28435 13572 28439 13628
rect 28439 13572 28495 13628
rect 28495 13572 28499 13628
rect 28435 13568 28499 13572
rect 28515 13628 28579 13632
rect 28515 13572 28519 13628
rect 28519 13572 28575 13628
rect 28575 13572 28579 13628
rect 28515 13568 28579 13572
rect 3884 13084 3948 13088
rect 3884 13028 3888 13084
rect 3888 13028 3944 13084
rect 3944 13028 3948 13084
rect 3884 13024 3948 13028
rect 3964 13084 4028 13088
rect 3964 13028 3968 13084
rect 3968 13028 4024 13084
rect 4024 13028 4028 13084
rect 3964 13024 4028 13028
rect 4044 13084 4108 13088
rect 4044 13028 4048 13084
rect 4048 13028 4104 13084
rect 4104 13028 4108 13084
rect 4044 13024 4108 13028
rect 4124 13084 4188 13088
rect 4124 13028 4128 13084
rect 4128 13028 4184 13084
rect 4184 13028 4188 13084
rect 4124 13024 4188 13028
rect 10853 13084 10917 13088
rect 10853 13028 10857 13084
rect 10857 13028 10913 13084
rect 10913 13028 10917 13084
rect 10853 13024 10917 13028
rect 10933 13084 10997 13088
rect 10933 13028 10937 13084
rect 10937 13028 10993 13084
rect 10993 13028 10997 13084
rect 10933 13024 10997 13028
rect 11013 13084 11077 13088
rect 11013 13028 11017 13084
rect 11017 13028 11073 13084
rect 11073 13028 11077 13084
rect 11013 13024 11077 13028
rect 11093 13084 11157 13088
rect 11093 13028 11097 13084
rect 11097 13028 11153 13084
rect 11153 13028 11157 13084
rect 11093 13024 11157 13028
rect 17822 13084 17886 13088
rect 17822 13028 17826 13084
rect 17826 13028 17882 13084
rect 17882 13028 17886 13084
rect 17822 13024 17886 13028
rect 17902 13084 17966 13088
rect 17902 13028 17906 13084
rect 17906 13028 17962 13084
rect 17962 13028 17966 13084
rect 17902 13024 17966 13028
rect 17982 13084 18046 13088
rect 17982 13028 17986 13084
rect 17986 13028 18042 13084
rect 18042 13028 18046 13084
rect 17982 13024 18046 13028
rect 18062 13084 18126 13088
rect 18062 13028 18066 13084
rect 18066 13028 18122 13084
rect 18122 13028 18126 13084
rect 18062 13024 18126 13028
rect 24791 13084 24855 13088
rect 24791 13028 24795 13084
rect 24795 13028 24851 13084
rect 24851 13028 24855 13084
rect 24791 13024 24855 13028
rect 24871 13084 24935 13088
rect 24871 13028 24875 13084
rect 24875 13028 24931 13084
rect 24931 13028 24935 13084
rect 24871 13024 24935 13028
rect 24951 13084 25015 13088
rect 24951 13028 24955 13084
rect 24955 13028 25011 13084
rect 25011 13028 25015 13084
rect 24951 13024 25015 13028
rect 25031 13084 25095 13088
rect 25031 13028 25035 13084
rect 25035 13028 25091 13084
rect 25091 13028 25095 13084
rect 25031 13024 25095 13028
rect 7368 12540 7432 12544
rect 7368 12484 7372 12540
rect 7372 12484 7428 12540
rect 7428 12484 7432 12540
rect 7368 12480 7432 12484
rect 7448 12540 7512 12544
rect 7448 12484 7452 12540
rect 7452 12484 7508 12540
rect 7508 12484 7512 12540
rect 7448 12480 7512 12484
rect 7528 12540 7592 12544
rect 7528 12484 7532 12540
rect 7532 12484 7588 12540
rect 7588 12484 7592 12540
rect 7528 12480 7592 12484
rect 7608 12540 7672 12544
rect 7608 12484 7612 12540
rect 7612 12484 7668 12540
rect 7668 12484 7672 12540
rect 7608 12480 7672 12484
rect 14337 12540 14401 12544
rect 14337 12484 14341 12540
rect 14341 12484 14397 12540
rect 14397 12484 14401 12540
rect 14337 12480 14401 12484
rect 14417 12540 14481 12544
rect 14417 12484 14421 12540
rect 14421 12484 14477 12540
rect 14477 12484 14481 12540
rect 14417 12480 14481 12484
rect 14497 12540 14561 12544
rect 14497 12484 14501 12540
rect 14501 12484 14557 12540
rect 14557 12484 14561 12540
rect 14497 12480 14561 12484
rect 14577 12540 14641 12544
rect 14577 12484 14581 12540
rect 14581 12484 14637 12540
rect 14637 12484 14641 12540
rect 14577 12480 14641 12484
rect 21306 12540 21370 12544
rect 21306 12484 21310 12540
rect 21310 12484 21366 12540
rect 21366 12484 21370 12540
rect 21306 12480 21370 12484
rect 21386 12540 21450 12544
rect 21386 12484 21390 12540
rect 21390 12484 21446 12540
rect 21446 12484 21450 12540
rect 21386 12480 21450 12484
rect 21466 12540 21530 12544
rect 21466 12484 21470 12540
rect 21470 12484 21526 12540
rect 21526 12484 21530 12540
rect 21466 12480 21530 12484
rect 21546 12540 21610 12544
rect 21546 12484 21550 12540
rect 21550 12484 21606 12540
rect 21606 12484 21610 12540
rect 21546 12480 21610 12484
rect 28275 12540 28339 12544
rect 28275 12484 28279 12540
rect 28279 12484 28335 12540
rect 28335 12484 28339 12540
rect 28275 12480 28339 12484
rect 28355 12540 28419 12544
rect 28355 12484 28359 12540
rect 28359 12484 28415 12540
rect 28415 12484 28419 12540
rect 28355 12480 28419 12484
rect 28435 12540 28499 12544
rect 28435 12484 28439 12540
rect 28439 12484 28495 12540
rect 28495 12484 28499 12540
rect 28435 12480 28499 12484
rect 28515 12540 28579 12544
rect 28515 12484 28519 12540
rect 28519 12484 28575 12540
rect 28575 12484 28579 12540
rect 28515 12480 28579 12484
rect 3884 11996 3948 12000
rect 3884 11940 3888 11996
rect 3888 11940 3944 11996
rect 3944 11940 3948 11996
rect 3884 11936 3948 11940
rect 3964 11996 4028 12000
rect 3964 11940 3968 11996
rect 3968 11940 4024 11996
rect 4024 11940 4028 11996
rect 3964 11936 4028 11940
rect 4044 11996 4108 12000
rect 4044 11940 4048 11996
rect 4048 11940 4104 11996
rect 4104 11940 4108 11996
rect 4044 11936 4108 11940
rect 4124 11996 4188 12000
rect 4124 11940 4128 11996
rect 4128 11940 4184 11996
rect 4184 11940 4188 11996
rect 4124 11936 4188 11940
rect 10853 11996 10917 12000
rect 10853 11940 10857 11996
rect 10857 11940 10913 11996
rect 10913 11940 10917 11996
rect 10853 11936 10917 11940
rect 10933 11996 10997 12000
rect 10933 11940 10937 11996
rect 10937 11940 10993 11996
rect 10993 11940 10997 11996
rect 10933 11936 10997 11940
rect 11013 11996 11077 12000
rect 11013 11940 11017 11996
rect 11017 11940 11073 11996
rect 11073 11940 11077 11996
rect 11013 11936 11077 11940
rect 11093 11996 11157 12000
rect 11093 11940 11097 11996
rect 11097 11940 11153 11996
rect 11153 11940 11157 11996
rect 11093 11936 11157 11940
rect 17822 11996 17886 12000
rect 17822 11940 17826 11996
rect 17826 11940 17882 11996
rect 17882 11940 17886 11996
rect 17822 11936 17886 11940
rect 17902 11996 17966 12000
rect 17902 11940 17906 11996
rect 17906 11940 17962 11996
rect 17962 11940 17966 11996
rect 17902 11936 17966 11940
rect 17982 11996 18046 12000
rect 17982 11940 17986 11996
rect 17986 11940 18042 11996
rect 18042 11940 18046 11996
rect 17982 11936 18046 11940
rect 18062 11996 18126 12000
rect 18062 11940 18066 11996
rect 18066 11940 18122 11996
rect 18122 11940 18126 11996
rect 18062 11936 18126 11940
rect 24791 11996 24855 12000
rect 24791 11940 24795 11996
rect 24795 11940 24851 11996
rect 24851 11940 24855 11996
rect 24791 11936 24855 11940
rect 24871 11996 24935 12000
rect 24871 11940 24875 11996
rect 24875 11940 24931 11996
rect 24931 11940 24935 11996
rect 24871 11936 24935 11940
rect 24951 11996 25015 12000
rect 24951 11940 24955 11996
rect 24955 11940 25011 11996
rect 25011 11940 25015 11996
rect 24951 11936 25015 11940
rect 25031 11996 25095 12000
rect 25031 11940 25035 11996
rect 25035 11940 25091 11996
rect 25091 11940 25095 11996
rect 25031 11936 25095 11940
rect 7368 11452 7432 11456
rect 7368 11396 7372 11452
rect 7372 11396 7428 11452
rect 7428 11396 7432 11452
rect 7368 11392 7432 11396
rect 7448 11452 7512 11456
rect 7448 11396 7452 11452
rect 7452 11396 7508 11452
rect 7508 11396 7512 11452
rect 7448 11392 7512 11396
rect 7528 11452 7592 11456
rect 7528 11396 7532 11452
rect 7532 11396 7588 11452
rect 7588 11396 7592 11452
rect 7528 11392 7592 11396
rect 7608 11452 7672 11456
rect 7608 11396 7612 11452
rect 7612 11396 7668 11452
rect 7668 11396 7672 11452
rect 7608 11392 7672 11396
rect 14337 11452 14401 11456
rect 14337 11396 14341 11452
rect 14341 11396 14397 11452
rect 14397 11396 14401 11452
rect 14337 11392 14401 11396
rect 14417 11452 14481 11456
rect 14417 11396 14421 11452
rect 14421 11396 14477 11452
rect 14477 11396 14481 11452
rect 14417 11392 14481 11396
rect 14497 11452 14561 11456
rect 14497 11396 14501 11452
rect 14501 11396 14557 11452
rect 14557 11396 14561 11452
rect 14497 11392 14561 11396
rect 14577 11452 14641 11456
rect 14577 11396 14581 11452
rect 14581 11396 14637 11452
rect 14637 11396 14641 11452
rect 14577 11392 14641 11396
rect 21306 11452 21370 11456
rect 21306 11396 21310 11452
rect 21310 11396 21366 11452
rect 21366 11396 21370 11452
rect 21306 11392 21370 11396
rect 21386 11452 21450 11456
rect 21386 11396 21390 11452
rect 21390 11396 21446 11452
rect 21446 11396 21450 11452
rect 21386 11392 21450 11396
rect 21466 11452 21530 11456
rect 21466 11396 21470 11452
rect 21470 11396 21526 11452
rect 21526 11396 21530 11452
rect 21466 11392 21530 11396
rect 21546 11452 21610 11456
rect 21546 11396 21550 11452
rect 21550 11396 21606 11452
rect 21606 11396 21610 11452
rect 21546 11392 21610 11396
rect 28275 11452 28339 11456
rect 28275 11396 28279 11452
rect 28279 11396 28335 11452
rect 28335 11396 28339 11452
rect 28275 11392 28339 11396
rect 28355 11452 28419 11456
rect 28355 11396 28359 11452
rect 28359 11396 28415 11452
rect 28415 11396 28419 11452
rect 28355 11392 28419 11396
rect 28435 11452 28499 11456
rect 28435 11396 28439 11452
rect 28439 11396 28495 11452
rect 28495 11396 28499 11452
rect 28435 11392 28499 11396
rect 28515 11452 28579 11456
rect 28515 11396 28519 11452
rect 28519 11396 28575 11452
rect 28575 11396 28579 11452
rect 28515 11392 28579 11396
rect 3884 10908 3948 10912
rect 3884 10852 3888 10908
rect 3888 10852 3944 10908
rect 3944 10852 3948 10908
rect 3884 10848 3948 10852
rect 3964 10908 4028 10912
rect 3964 10852 3968 10908
rect 3968 10852 4024 10908
rect 4024 10852 4028 10908
rect 3964 10848 4028 10852
rect 4044 10908 4108 10912
rect 4044 10852 4048 10908
rect 4048 10852 4104 10908
rect 4104 10852 4108 10908
rect 4044 10848 4108 10852
rect 4124 10908 4188 10912
rect 4124 10852 4128 10908
rect 4128 10852 4184 10908
rect 4184 10852 4188 10908
rect 4124 10848 4188 10852
rect 10853 10908 10917 10912
rect 10853 10852 10857 10908
rect 10857 10852 10913 10908
rect 10913 10852 10917 10908
rect 10853 10848 10917 10852
rect 10933 10908 10997 10912
rect 10933 10852 10937 10908
rect 10937 10852 10993 10908
rect 10993 10852 10997 10908
rect 10933 10848 10997 10852
rect 11013 10908 11077 10912
rect 11013 10852 11017 10908
rect 11017 10852 11073 10908
rect 11073 10852 11077 10908
rect 11013 10848 11077 10852
rect 11093 10908 11157 10912
rect 11093 10852 11097 10908
rect 11097 10852 11153 10908
rect 11153 10852 11157 10908
rect 11093 10848 11157 10852
rect 17822 10908 17886 10912
rect 17822 10852 17826 10908
rect 17826 10852 17882 10908
rect 17882 10852 17886 10908
rect 17822 10848 17886 10852
rect 17902 10908 17966 10912
rect 17902 10852 17906 10908
rect 17906 10852 17962 10908
rect 17962 10852 17966 10908
rect 17902 10848 17966 10852
rect 17982 10908 18046 10912
rect 17982 10852 17986 10908
rect 17986 10852 18042 10908
rect 18042 10852 18046 10908
rect 17982 10848 18046 10852
rect 18062 10908 18126 10912
rect 18062 10852 18066 10908
rect 18066 10852 18122 10908
rect 18122 10852 18126 10908
rect 18062 10848 18126 10852
rect 24791 10908 24855 10912
rect 24791 10852 24795 10908
rect 24795 10852 24851 10908
rect 24851 10852 24855 10908
rect 24791 10848 24855 10852
rect 24871 10908 24935 10912
rect 24871 10852 24875 10908
rect 24875 10852 24931 10908
rect 24931 10852 24935 10908
rect 24871 10848 24935 10852
rect 24951 10908 25015 10912
rect 24951 10852 24955 10908
rect 24955 10852 25011 10908
rect 25011 10852 25015 10908
rect 24951 10848 25015 10852
rect 25031 10908 25095 10912
rect 25031 10852 25035 10908
rect 25035 10852 25091 10908
rect 25091 10852 25095 10908
rect 25031 10848 25095 10852
rect 7368 10364 7432 10368
rect 7368 10308 7372 10364
rect 7372 10308 7428 10364
rect 7428 10308 7432 10364
rect 7368 10304 7432 10308
rect 7448 10364 7512 10368
rect 7448 10308 7452 10364
rect 7452 10308 7508 10364
rect 7508 10308 7512 10364
rect 7448 10304 7512 10308
rect 7528 10364 7592 10368
rect 7528 10308 7532 10364
rect 7532 10308 7588 10364
rect 7588 10308 7592 10364
rect 7528 10304 7592 10308
rect 7608 10364 7672 10368
rect 7608 10308 7612 10364
rect 7612 10308 7668 10364
rect 7668 10308 7672 10364
rect 7608 10304 7672 10308
rect 14337 10364 14401 10368
rect 14337 10308 14341 10364
rect 14341 10308 14397 10364
rect 14397 10308 14401 10364
rect 14337 10304 14401 10308
rect 14417 10364 14481 10368
rect 14417 10308 14421 10364
rect 14421 10308 14477 10364
rect 14477 10308 14481 10364
rect 14417 10304 14481 10308
rect 14497 10364 14561 10368
rect 14497 10308 14501 10364
rect 14501 10308 14557 10364
rect 14557 10308 14561 10364
rect 14497 10304 14561 10308
rect 14577 10364 14641 10368
rect 14577 10308 14581 10364
rect 14581 10308 14637 10364
rect 14637 10308 14641 10364
rect 14577 10304 14641 10308
rect 21306 10364 21370 10368
rect 21306 10308 21310 10364
rect 21310 10308 21366 10364
rect 21366 10308 21370 10364
rect 21306 10304 21370 10308
rect 21386 10364 21450 10368
rect 21386 10308 21390 10364
rect 21390 10308 21446 10364
rect 21446 10308 21450 10364
rect 21386 10304 21450 10308
rect 21466 10364 21530 10368
rect 21466 10308 21470 10364
rect 21470 10308 21526 10364
rect 21526 10308 21530 10364
rect 21466 10304 21530 10308
rect 21546 10364 21610 10368
rect 21546 10308 21550 10364
rect 21550 10308 21606 10364
rect 21606 10308 21610 10364
rect 21546 10304 21610 10308
rect 28275 10364 28339 10368
rect 28275 10308 28279 10364
rect 28279 10308 28335 10364
rect 28335 10308 28339 10364
rect 28275 10304 28339 10308
rect 28355 10364 28419 10368
rect 28355 10308 28359 10364
rect 28359 10308 28415 10364
rect 28415 10308 28419 10364
rect 28355 10304 28419 10308
rect 28435 10364 28499 10368
rect 28435 10308 28439 10364
rect 28439 10308 28495 10364
rect 28495 10308 28499 10364
rect 28435 10304 28499 10308
rect 28515 10364 28579 10368
rect 28515 10308 28519 10364
rect 28519 10308 28575 10364
rect 28575 10308 28579 10364
rect 28515 10304 28579 10308
rect 3884 9820 3948 9824
rect 3884 9764 3888 9820
rect 3888 9764 3944 9820
rect 3944 9764 3948 9820
rect 3884 9760 3948 9764
rect 3964 9820 4028 9824
rect 3964 9764 3968 9820
rect 3968 9764 4024 9820
rect 4024 9764 4028 9820
rect 3964 9760 4028 9764
rect 4044 9820 4108 9824
rect 4044 9764 4048 9820
rect 4048 9764 4104 9820
rect 4104 9764 4108 9820
rect 4044 9760 4108 9764
rect 4124 9820 4188 9824
rect 4124 9764 4128 9820
rect 4128 9764 4184 9820
rect 4184 9764 4188 9820
rect 4124 9760 4188 9764
rect 10853 9820 10917 9824
rect 10853 9764 10857 9820
rect 10857 9764 10913 9820
rect 10913 9764 10917 9820
rect 10853 9760 10917 9764
rect 10933 9820 10997 9824
rect 10933 9764 10937 9820
rect 10937 9764 10993 9820
rect 10993 9764 10997 9820
rect 10933 9760 10997 9764
rect 11013 9820 11077 9824
rect 11013 9764 11017 9820
rect 11017 9764 11073 9820
rect 11073 9764 11077 9820
rect 11013 9760 11077 9764
rect 11093 9820 11157 9824
rect 11093 9764 11097 9820
rect 11097 9764 11153 9820
rect 11153 9764 11157 9820
rect 11093 9760 11157 9764
rect 17822 9820 17886 9824
rect 17822 9764 17826 9820
rect 17826 9764 17882 9820
rect 17882 9764 17886 9820
rect 17822 9760 17886 9764
rect 17902 9820 17966 9824
rect 17902 9764 17906 9820
rect 17906 9764 17962 9820
rect 17962 9764 17966 9820
rect 17902 9760 17966 9764
rect 17982 9820 18046 9824
rect 17982 9764 17986 9820
rect 17986 9764 18042 9820
rect 18042 9764 18046 9820
rect 17982 9760 18046 9764
rect 18062 9820 18126 9824
rect 18062 9764 18066 9820
rect 18066 9764 18122 9820
rect 18122 9764 18126 9820
rect 18062 9760 18126 9764
rect 24791 9820 24855 9824
rect 24791 9764 24795 9820
rect 24795 9764 24851 9820
rect 24851 9764 24855 9820
rect 24791 9760 24855 9764
rect 24871 9820 24935 9824
rect 24871 9764 24875 9820
rect 24875 9764 24931 9820
rect 24931 9764 24935 9820
rect 24871 9760 24935 9764
rect 24951 9820 25015 9824
rect 24951 9764 24955 9820
rect 24955 9764 25011 9820
rect 25011 9764 25015 9820
rect 24951 9760 25015 9764
rect 25031 9820 25095 9824
rect 25031 9764 25035 9820
rect 25035 9764 25091 9820
rect 25091 9764 25095 9820
rect 25031 9760 25095 9764
rect 7368 9276 7432 9280
rect 7368 9220 7372 9276
rect 7372 9220 7428 9276
rect 7428 9220 7432 9276
rect 7368 9216 7432 9220
rect 7448 9276 7512 9280
rect 7448 9220 7452 9276
rect 7452 9220 7508 9276
rect 7508 9220 7512 9276
rect 7448 9216 7512 9220
rect 7528 9276 7592 9280
rect 7528 9220 7532 9276
rect 7532 9220 7588 9276
rect 7588 9220 7592 9276
rect 7528 9216 7592 9220
rect 7608 9276 7672 9280
rect 7608 9220 7612 9276
rect 7612 9220 7668 9276
rect 7668 9220 7672 9276
rect 7608 9216 7672 9220
rect 14337 9276 14401 9280
rect 14337 9220 14341 9276
rect 14341 9220 14397 9276
rect 14397 9220 14401 9276
rect 14337 9216 14401 9220
rect 14417 9276 14481 9280
rect 14417 9220 14421 9276
rect 14421 9220 14477 9276
rect 14477 9220 14481 9276
rect 14417 9216 14481 9220
rect 14497 9276 14561 9280
rect 14497 9220 14501 9276
rect 14501 9220 14557 9276
rect 14557 9220 14561 9276
rect 14497 9216 14561 9220
rect 14577 9276 14641 9280
rect 14577 9220 14581 9276
rect 14581 9220 14637 9276
rect 14637 9220 14641 9276
rect 14577 9216 14641 9220
rect 21306 9276 21370 9280
rect 21306 9220 21310 9276
rect 21310 9220 21366 9276
rect 21366 9220 21370 9276
rect 21306 9216 21370 9220
rect 21386 9276 21450 9280
rect 21386 9220 21390 9276
rect 21390 9220 21446 9276
rect 21446 9220 21450 9276
rect 21386 9216 21450 9220
rect 21466 9276 21530 9280
rect 21466 9220 21470 9276
rect 21470 9220 21526 9276
rect 21526 9220 21530 9276
rect 21466 9216 21530 9220
rect 21546 9276 21610 9280
rect 21546 9220 21550 9276
rect 21550 9220 21606 9276
rect 21606 9220 21610 9276
rect 21546 9216 21610 9220
rect 28275 9276 28339 9280
rect 28275 9220 28279 9276
rect 28279 9220 28335 9276
rect 28335 9220 28339 9276
rect 28275 9216 28339 9220
rect 28355 9276 28419 9280
rect 28355 9220 28359 9276
rect 28359 9220 28415 9276
rect 28415 9220 28419 9276
rect 28355 9216 28419 9220
rect 28435 9276 28499 9280
rect 28435 9220 28439 9276
rect 28439 9220 28495 9276
rect 28495 9220 28499 9276
rect 28435 9216 28499 9220
rect 28515 9276 28579 9280
rect 28515 9220 28519 9276
rect 28519 9220 28575 9276
rect 28575 9220 28579 9276
rect 28515 9216 28579 9220
rect 3884 8732 3948 8736
rect 3884 8676 3888 8732
rect 3888 8676 3944 8732
rect 3944 8676 3948 8732
rect 3884 8672 3948 8676
rect 3964 8732 4028 8736
rect 3964 8676 3968 8732
rect 3968 8676 4024 8732
rect 4024 8676 4028 8732
rect 3964 8672 4028 8676
rect 4044 8732 4108 8736
rect 4044 8676 4048 8732
rect 4048 8676 4104 8732
rect 4104 8676 4108 8732
rect 4044 8672 4108 8676
rect 4124 8732 4188 8736
rect 4124 8676 4128 8732
rect 4128 8676 4184 8732
rect 4184 8676 4188 8732
rect 4124 8672 4188 8676
rect 10853 8732 10917 8736
rect 10853 8676 10857 8732
rect 10857 8676 10913 8732
rect 10913 8676 10917 8732
rect 10853 8672 10917 8676
rect 10933 8732 10997 8736
rect 10933 8676 10937 8732
rect 10937 8676 10993 8732
rect 10993 8676 10997 8732
rect 10933 8672 10997 8676
rect 11013 8732 11077 8736
rect 11013 8676 11017 8732
rect 11017 8676 11073 8732
rect 11073 8676 11077 8732
rect 11013 8672 11077 8676
rect 11093 8732 11157 8736
rect 11093 8676 11097 8732
rect 11097 8676 11153 8732
rect 11153 8676 11157 8732
rect 11093 8672 11157 8676
rect 17822 8732 17886 8736
rect 17822 8676 17826 8732
rect 17826 8676 17882 8732
rect 17882 8676 17886 8732
rect 17822 8672 17886 8676
rect 17902 8732 17966 8736
rect 17902 8676 17906 8732
rect 17906 8676 17962 8732
rect 17962 8676 17966 8732
rect 17902 8672 17966 8676
rect 17982 8732 18046 8736
rect 17982 8676 17986 8732
rect 17986 8676 18042 8732
rect 18042 8676 18046 8732
rect 17982 8672 18046 8676
rect 18062 8732 18126 8736
rect 18062 8676 18066 8732
rect 18066 8676 18122 8732
rect 18122 8676 18126 8732
rect 18062 8672 18126 8676
rect 24791 8732 24855 8736
rect 24791 8676 24795 8732
rect 24795 8676 24851 8732
rect 24851 8676 24855 8732
rect 24791 8672 24855 8676
rect 24871 8732 24935 8736
rect 24871 8676 24875 8732
rect 24875 8676 24931 8732
rect 24931 8676 24935 8732
rect 24871 8672 24935 8676
rect 24951 8732 25015 8736
rect 24951 8676 24955 8732
rect 24955 8676 25011 8732
rect 25011 8676 25015 8732
rect 24951 8672 25015 8676
rect 25031 8732 25095 8736
rect 25031 8676 25035 8732
rect 25035 8676 25091 8732
rect 25091 8676 25095 8732
rect 25031 8672 25095 8676
rect 7368 8188 7432 8192
rect 7368 8132 7372 8188
rect 7372 8132 7428 8188
rect 7428 8132 7432 8188
rect 7368 8128 7432 8132
rect 7448 8188 7512 8192
rect 7448 8132 7452 8188
rect 7452 8132 7508 8188
rect 7508 8132 7512 8188
rect 7448 8128 7512 8132
rect 7528 8188 7592 8192
rect 7528 8132 7532 8188
rect 7532 8132 7588 8188
rect 7588 8132 7592 8188
rect 7528 8128 7592 8132
rect 7608 8188 7672 8192
rect 7608 8132 7612 8188
rect 7612 8132 7668 8188
rect 7668 8132 7672 8188
rect 7608 8128 7672 8132
rect 14337 8188 14401 8192
rect 14337 8132 14341 8188
rect 14341 8132 14397 8188
rect 14397 8132 14401 8188
rect 14337 8128 14401 8132
rect 14417 8188 14481 8192
rect 14417 8132 14421 8188
rect 14421 8132 14477 8188
rect 14477 8132 14481 8188
rect 14417 8128 14481 8132
rect 14497 8188 14561 8192
rect 14497 8132 14501 8188
rect 14501 8132 14557 8188
rect 14557 8132 14561 8188
rect 14497 8128 14561 8132
rect 14577 8188 14641 8192
rect 14577 8132 14581 8188
rect 14581 8132 14637 8188
rect 14637 8132 14641 8188
rect 14577 8128 14641 8132
rect 21306 8188 21370 8192
rect 21306 8132 21310 8188
rect 21310 8132 21366 8188
rect 21366 8132 21370 8188
rect 21306 8128 21370 8132
rect 21386 8188 21450 8192
rect 21386 8132 21390 8188
rect 21390 8132 21446 8188
rect 21446 8132 21450 8188
rect 21386 8128 21450 8132
rect 21466 8188 21530 8192
rect 21466 8132 21470 8188
rect 21470 8132 21526 8188
rect 21526 8132 21530 8188
rect 21466 8128 21530 8132
rect 21546 8188 21610 8192
rect 21546 8132 21550 8188
rect 21550 8132 21606 8188
rect 21606 8132 21610 8188
rect 21546 8128 21610 8132
rect 28275 8188 28339 8192
rect 28275 8132 28279 8188
rect 28279 8132 28335 8188
rect 28335 8132 28339 8188
rect 28275 8128 28339 8132
rect 28355 8188 28419 8192
rect 28355 8132 28359 8188
rect 28359 8132 28415 8188
rect 28415 8132 28419 8188
rect 28355 8128 28419 8132
rect 28435 8188 28499 8192
rect 28435 8132 28439 8188
rect 28439 8132 28495 8188
rect 28495 8132 28499 8188
rect 28435 8128 28499 8132
rect 28515 8188 28579 8192
rect 28515 8132 28519 8188
rect 28519 8132 28575 8188
rect 28575 8132 28579 8188
rect 28515 8128 28579 8132
rect 3884 7644 3948 7648
rect 3884 7588 3888 7644
rect 3888 7588 3944 7644
rect 3944 7588 3948 7644
rect 3884 7584 3948 7588
rect 3964 7644 4028 7648
rect 3964 7588 3968 7644
rect 3968 7588 4024 7644
rect 4024 7588 4028 7644
rect 3964 7584 4028 7588
rect 4044 7644 4108 7648
rect 4044 7588 4048 7644
rect 4048 7588 4104 7644
rect 4104 7588 4108 7644
rect 4044 7584 4108 7588
rect 4124 7644 4188 7648
rect 4124 7588 4128 7644
rect 4128 7588 4184 7644
rect 4184 7588 4188 7644
rect 4124 7584 4188 7588
rect 10853 7644 10917 7648
rect 10853 7588 10857 7644
rect 10857 7588 10913 7644
rect 10913 7588 10917 7644
rect 10853 7584 10917 7588
rect 10933 7644 10997 7648
rect 10933 7588 10937 7644
rect 10937 7588 10993 7644
rect 10993 7588 10997 7644
rect 10933 7584 10997 7588
rect 11013 7644 11077 7648
rect 11013 7588 11017 7644
rect 11017 7588 11073 7644
rect 11073 7588 11077 7644
rect 11013 7584 11077 7588
rect 11093 7644 11157 7648
rect 11093 7588 11097 7644
rect 11097 7588 11153 7644
rect 11153 7588 11157 7644
rect 11093 7584 11157 7588
rect 17822 7644 17886 7648
rect 17822 7588 17826 7644
rect 17826 7588 17882 7644
rect 17882 7588 17886 7644
rect 17822 7584 17886 7588
rect 17902 7644 17966 7648
rect 17902 7588 17906 7644
rect 17906 7588 17962 7644
rect 17962 7588 17966 7644
rect 17902 7584 17966 7588
rect 17982 7644 18046 7648
rect 17982 7588 17986 7644
rect 17986 7588 18042 7644
rect 18042 7588 18046 7644
rect 17982 7584 18046 7588
rect 18062 7644 18126 7648
rect 18062 7588 18066 7644
rect 18066 7588 18122 7644
rect 18122 7588 18126 7644
rect 18062 7584 18126 7588
rect 24791 7644 24855 7648
rect 24791 7588 24795 7644
rect 24795 7588 24851 7644
rect 24851 7588 24855 7644
rect 24791 7584 24855 7588
rect 24871 7644 24935 7648
rect 24871 7588 24875 7644
rect 24875 7588 24931 7644
rect 24931 7588 24935 7644
rect 24871 7584 24935 7588
rect 24951 7644 25015 7648
rect 24951 7588 24955 7644
rect 24955 7588 25011 7644
rect 25011 7588 25015 7644
rect 24951 7584 25015 7588
rect 25031 7644 25095 7648
rect 25031 7588 25035 7644
rect 25035 7588 25091 7644
rect 25091 7588 25095 7644
rect 25031 7584 25095 7588
rect 7368 7100 7432 7104
rect 7368 7044 7372 7100
rect 7372 7044 7428 7100
rect 7428 7044 7432 7100
rect 7368 7040 7432 7044
rect 7448 7100 7512 7104
rect 7448 7044 7452 7100
rect 7452 7044 7508 7100
rect 7508 7044 7512 7100
rect 7448 7040 7512 7044
rect 7528 7100 7592 7104
rect 7528 7044 7532 7100
rect 7532 7044 7588 7100
rect 7588 7044 7592 7100
rect 7528 7040 7592 7044
rect 7608 7100 7672 7104
rect 7608 7044 7612 7100
rect 7612 7044 7668 7100
rect 7668 7044 7672 7100
rect 7608 7040 7672 7044
rect 14337 7100 14401 7104
rect 14337 7044 14341 7100
rect 14341 7044 14397 7100
rect 14397 7044 14401 7100
rect 14337 7040 14401 7044
rect 14417 7100 14481 7104
rect 14417 7044 14421 7100
rect 14421 7044 14477 7100
rect 14477 7044 14481 7100
rect 14417 7040 14481 7044
rect 14497 7100 14561 7104
rect 14497 7044 14501 7100
rect 14501 7044 14557 7100
rect 14557 7044 14561 7100
rect 14497 7040 14561 7044
rect 14577 7100 14641 7104
rect 14577 7044 14581 7100
rect 14581 7044 14637 7100
rect 14637 7044 14641 7100
rect 14577 7040 14641 7044
rect 21306 7100 21370 7104
rect 21306 7044 21310 7100
rect 21310 7044 21366 7100
rect 21366 7044 21370 7100
rect 21306 7040 21370 7044
rect 21386 7100 21450 7104
rect 21386 7044 21390 7100
rect 21390 7044 21446 7100
rect 21446 7044 21450 7100
rect 21386 7040 21450 7044
rect 21466 7100 21530 7104
rect 21466 7044 21470 7100
rect 21470 7044 21526 7100
rect 21526 7044 21530 7100
rect 21466 7040 21530 7044
rect 21546 7100 21610 7104
rect 21546 7044 21550 7100
rect 21550 7044 21606 7100
rect 21606 7044 21610 7100
rect 21546 7040 21610 7044
rect 28275 7100 28339 7104
rect 28275 7044 28279 7100
rect 28279 7044 28335 7100
rect 28335 7044 28339 7100
rect 28275 7040 28339 7044
rect 28355 7100 28419 7104
rect 28355 7044 28359 7100
rect 28359 7044 28415 7100
rect 28415 7044 28419 7100
rect 28355 7040 28419 7044
rect 28435 7100 28499 7104
rect 28435 7044 28439 7100
rect 28439 7044 28495 7100
rect 28495 7044 28499 7100
rect 28435 7040 28499 7044
rect 28515 7100 28579 7104
rect 28515 7044 28519 7100
rect 28519 7044 28575 7100
rect 28575 7044 28579 7100
rect 28515 7040 28579 7044
rect 3884 6556 3948 6560
rect 3884 6500 3888 6556
rect 3888 6500 3944 6556
rect 3944 6500 3948 6556
rect 3884 6496 3948 6500
rect 3964 6556 4028 6560
rect 3964 6500 3968 6556
rect 3968 6500 4024 6556
rect 4024 6500 4028 6556
rect 3964 6496 4028 6500
rect 4044 6556 4108 6560
rect 4044 6500 4048 6556
rect 4048 6500 4104 6556
rect 4104 6500 4108 6556
rect 4044 6496 4108 6500
rect 4124 6556 4188 6560
rect 4124 6500 4128 6556
rect 4128 6500 4184 6556
rect 4184 6500 4188 6556
rect 4124 6496 4188 6500
rect 10853 6556 10917 6560
rect 10853 6500 10857 6556
rect 10857 6500 10913 6556
rect 10913 6500 10917 6556
rect 10853 6496 10917 6500
rect 10933 6556 10997 6560
rect 10933 6500 10937 6556
rect 10937 6500 10993 6556
rect 10993 6500 10997 6556
rect 10933 6496 10997 6500
rect 11013 6556 11077 6560
rect 11013 6500 11017 6556
rect 11017 6500 11073 6556
rect 11073 6500 11077 6556
rect 11013 6496 11077 6500
rect 11093 6556 11157 6560
rect 11093 6500 11097 6556
rect 11097 6500 11153 6556
rect 11153 6500 11157 6556
rect 11093 6496 11157 6500
rect 17822 6556 17886 6560
rect 17822 6500 17826 6556
rect 17826 6500 17882 6556
rect 17882 6500 17886 6556
rect 17822 6496 17886 6500
rect 17902 6556 17966 6560
rect 17902 6500 17906 6556
rect 17906 6500 17962 6556
rect 17962 6500 17966 6556
rect 17902 6496 17966 6500
rect 17982 6556 18046 6560
rect 17982 6500 17986 6556
rect 17986 6500 18042 6556
rect 18042 6500 18046 6556
rect 17982 6496 18046 6500
rect 18062 6556 18126 6560
rect 18062 6500 18066 6556
rect 18066 6500 18122 6556
rect 18122 6500 18126 6556
rect 18062 6496 18126 6500
rect 24791 6556 24855 6560
rect 24791 6500 24795 6556
rect 24795 6500 24851 6556
rect 24851 6500 24855 6556
rect 24791 6496 24855 6500
rect 24871 6556 24935 6560
rect 24871 6500 24875 6556
rect 24875 6500 24931 6556
rect 24931 6500 24935 6556
rect 24871 6496 24935 6500
rect 24951 6556 25015 6560
rect 24951 6500 24955 6556
rect 24955 6500 25011 6556
rect 25011 6500 25015 6556
rect 24951 6496 25015 6500
rect 25031 6556 25095 6560
rect 25031 6500 25035 6556
rect 25035 6500 25091 6556
rect 25091 6500 25095 6556
rect 25031 6496 25095 6500
rect 7368 6012 7432 6016
rect 7368 5956 7372 6012
rect 7372 5956 7428 6012
rect 7428 5956 7432 6012
rect 7368 5952 7432 5956
rect 7448 6012 7512 6016
rect 7448 5956 7452 6012
rect 7452 5956 7508 6012
rect 7508 5956 7512 6012
rect 7448 5952 7512 5956
rect 7528 6012 7592 6016
rect 7528 5956 7532 6012
rect 7532 5956 7588 6012
rect 7588 5956 7592 6012
rect 7528 5952 7592 5956
rect 7608 6012 7672 6016
rect 7608 5956 7612 6012
rect 7612 5956 7668 6012
rect 7668 5956 7672 6012
rect 7608 5952 7672 5956
rect 14337 6012 14401 6016
rect 14337 5956 14341 6012
rect 14341 5956 14397 6012
rect 14397 5956 14401 6012
rect 14337 5952 14401 5956
rect 14417 6012 14481 6016
rect 14417 5956 14421 6012
rect 14421 5956 14477 6012
rect 14477 5956 14481 6012
rect 14417 5952 14481 5956
rect 14497 6012 14561 6016
rect 14497 5956 14501 6012
rect 14501 5956 14557 6012
rect 14557 5956 14561 6012
rect 14497 5952 14561 5956
rect 14577 6012 14641 6016
rect 14577 5956 14581 6012
rect 14581 5956 14637 6012
rect 14637 5956 14641 6012
rect 14577 5952 14641 5956
rect 21306 6012 21370 6016
rect 21306 5956 21310 6012
rect 21310 5956 21366 6012
rect 21366 5956 21370 6012
rect 21306 5952 21370 5956
rect 21386 6012 21450 6016
rect 21386 5956 21390 6012
rect 21390 5956 21446 6012
rect 21446 5956 21450 6012
rect 21386 5952 21450 5956
rect 21466 6012 21530 6016
rect 21466 5956 21470 6012
rect 21470 5956 21526 6012
rect 21526 5956 21530 6012
rect 21466 5952 21530 5956
rect 21546 6012 21610 6016
rect 21546 5956 21550 6012
rect 21550 5956 21606 6012
rect 21606 5956 21610 6012
rect 21546 5952 21610 5956
rect 28275 6012 28339 6016
rect 28275 5956 28279 6012
rect 28279 5956 28335 6012
rect 28335 5956 28339 6012
rect 28275 5952 28339 5956
rect 28355 6012 28419 6016
rect 28355 5956 28359 6012
rect 28359 5956 28415 6012
rect 28415 5956 28419 6012
rect 28355 5952 28419 5956
rect 28435 6012 28499 6016
rect 28435 5956 28439 6012
rect 28439 5956 28495 6012
rect 28495 5956 28499 6012
rect 28435 5952 28499 5956
rect 28515 6012 28579 6016
rect 28515 5956 28519 6012
rect 28519 5956 28575 6012
rect 28575 5956 28579 6012
rect 28515 5952 28579 5956
rect 3884 5468 3948 5472
rect 3884 5412 3888 5468
rect 3888 5412 3944 5468
rect 3944 5412 3948 5468
rect 3884 5408 3948 5412
rect 3964 5468 4028 5472
rect 3964 5412 3968 5468
rect 3968 5412 4024 5468
rect 4024 5412 4028 5468
rect 3964 5408 4028 5412
rect 4044 5468 4108 5472
rect 4044 5412 4048 5468
rect 4048 5412 4104 5468
rect 4104 5412 4108 5468
rect 4044 5408 4108 5412
rect 4124 5468 4188 5472
rect 4124 5412 4128 5468
rect 4128 5412 4184 5468
rect 4184 5412 4188 5468
rect 4124 5408 4188 5412
rect 10853 5468 10917 5472
rect 10853 5412 10857 5468
rect 10857 5412 10913 5468
rect 10913 5412 10917 5468
rect 10853 5408 10917 5412
rect 10933 5468 10997 5472
rect 10933 5412 10937 5468
rect 10937 5412 10993 5468
rect 10993 5412 10997 5468
rect 10933 5408 10997 5412
rect 11013 5468 11077 5472
rect 11013 5412 11017 5468
rect 11017 5412 11073 5468
rect 11073 5412 11077 5468
rect 11013 5408 11077 5412
rect 11093 5468 11157 5472
rect 11093 5412 11097 5468
rect 11097 5412 11153 5468
rect 11153 5412 11157 5468
rect 11093 5408 11157 5412
rect 17822 5468 17886 5472
rect 17822 5412 17826 5468
rect 17826 5412 17882 5468
rect 17882 5412 17886 5468
rect 17822 5408 17886 5412
rect 17902 5468 17966 5472
rect 17902 5412 17906 5468
rect 17906 5412 17962 5468
rect 17962 5412 17966 5468
rect 17902 5408 17966 5412
rect 17982 5468 18046 5472
rect 17982 5412 17986 5468
rect 17986 5412 18042 5468
rect 18042 5412 18046 5468
rect 17982 5408 18046 5412
rect 18062 5468 18126 5472
rect 18062 5412 18066 5468
rect 18066 5412 18122 5468
rect 18122 5412 18126 5468
rect 18062 5408 18126 5412
rect 24791 5468 24855 5472
rect 24791 5412 24795 5468
rect 24795 5412 24851 5468
rect 24851 5412 24855 5468
rect 24791 5408 24855 5412
rect 24871 5468 24935 5472
rect 24871 5412 24875 5468
rect 24875 5412 24931 5468
rect 24931 5412 24935 5468
rect 24871 5408 24935 5412
rect 24951 5468 25015 5472
rect 24951 5412 24955 5468
rect 24955 5412 25011 5468
rect 25011 5412 25015 5468
rect 24951 5408 25015 5412
rect 25031 5468 25095 5472
rect 25031 5412 25035 5468
rect 25035 5412 25091 5468
rect 25091 5412 25095 5468
rect 25031 5408 25095 5412
rect 7368 4924 7432 4928
rect 7368 4868 7372 4924
rect 7372 4868 7428 4924
rect 7428 4868 7432 4924
rect 7368 4864 7432 4868
rect 7448 4924 7512 4928
rect 7448 4868 7452 4924
rect 7452 4868 7508 4924
rect 7508 4868 7512 4924
rect 7448 4864 7512 4868
rect 7528 4924 7592 4928
rect 7528 4868 7532 4924
rect 7532 4868 7588 4924
rect 7588 4868 7592 4924
rect 7528 4864 7592 4868
rect 7608 4924 7672 4928
rect 7608 4868 7612 4924
rect 7612 4868 7668 4924
rect 7668 4868 7672 4924
rect 7608 4864 7672 4868
rect 14337 4924 14401 4928
rect 14337 4868 14341 4924
rect 14341 4868 14397 4924
rect 14397 4868 14401 4924
rect 14337 4864 14401 4868
rect 14417 4924 14481 4928
rect 14417 4868 14421 4924
rect 14421 4868 14477 4924
rect 14477 4868 14481 4924
rect 14417 4864 14481 4868
rect 14497 4924 14561 4928
rect 14497 4868 14501 4924
rect 14501 4868 14557 4924
rect 14557 4868 14561 4924
rect 14497 4864 14561 4868
rect 14577 4924 14641 4928
rect 14577 4868 14581 4924
rect 14581 4868 14637 4924
rect 14637 4868 14641 4924
rect 14577 4864 14641 4868
rect 21306 4924 21370 4928
rect 21306 4868 21310 4924
rect 21310 4868 21366 4924
rect 21366 4868 21370 4924
rect 21306 4864 21370 4868
rect 21386 4924 21450 4928
rect 21386 4868 21390 4924
rect 21390 4868 21446 4924
rect 21446 4868 21450 4924
rect 21386 4864 21450 4868
rect 21466 4924 21530 4928
rect 21466 4868 21470 4924
rect 21470 4868 21526 4924
rect 21526 4868 21530 4924
rect 21466 4864 21530 4868
rect 21546 4924 21610 4928
rect 21546 4868 21550 4924
rect 21550 4868 21606 4924
rect 21606 4868 21610 4924
rect 21546 4864 21610 4868
rect 28275 4924 28339 4928
rect 28275 4868 28279 4924
rect 28279 4868 28335 4924
rect 28335 4868 28339 4924
rect 28275 4864 28339 4868
rect 28355 4924 28419 4928
rect 28355 4868 28359 4924
rect 28359 4868 28415 4924
rect 28415 4868 28419 4924
rect 28355 4864 28419 4868
rect 28435 4924 28499 4928
rect 28435 4868 28439 4924
rect 28439 4868 28495 4924
rect 28495 4868 28499 4924
rect 28435 4864 28499 4868
rect 28515 4924 28579 4928
rect 28515 4868 28519 4924
rect 28519 4868 28575 4924
rect 28575 4868 28579 4924
rect 28515 4864 28579 4868
rect 3884 4380 3948 4384
rect 3884 4324 3888 4380
rect 3888 4324 3944 4380
rect 3944 4324 3948 4380
rect 3884 4320 3948 4324
rect 3964 4380 4028 4384
rect 3964 4324 3968 4380
rect 3968 4324 4024 4380
rect 4024 4324 4028 4380
rect 3964 4320 4028 4324
rect 4044 4380 4108 4384
rect 4044 4324 4048 4380
rect 4048 4324 4104 4380
rect 4104 4324 4108 4380
rect 4044 4320 4108 4324
rect 4124 4380 4188 4384
rect 4124 4324 4128 4380
rect 4128 4324 4184 4380
rect 4184 4324 4188 4380
rect 4124 4320 4188 4324
rect 10853 4380 10917 4384
rect 10853 4324 10857 4380
rect 10857 4324 10913 4380
rect 10913 4324 10917 4380
rect 10853 4320 10917 4324
rect 10933 4380 10997 4384
rect 10933 4324 10937 4380
rect 10937 4324 10993 4380
rect 10993 4324 10997 4380
rect 10933 4320 10997 4324
rect 11013 4380 11077 4384
rect 11013 4324 11017 4380
rect 11017 4324 11073 4380
rect 11073 4324 11077 4380
rect 11013 4320 11077 4324
rect 11093 4380 11157 4384
rect 11093 4324 11097 4380
rect 11097 4324 11153 4380
rect 11153 4324 11157 4380
rect 11093 4320 11157 4324
rect 17822 4380 17886 4384
rect 17822 4324 17826 4380
rect 17826 4324 17882 4380
rect 17882 4324 17886 4380
rect 17822 4320 17886 4324
rect 17902 4380 17966 4384
rect 17902 4324 17906 4380
rect 17906 4324 17962 4380
rect 17962 4324 17966 4380
rect 17902 4320 17966 4324
rect 17982 4380 18046 4384
rect 17982 4324 17986 4380
rect 17986 4324 18042 4380
rect 18042 4324 18046 4380
rect 17982 4320 18046 4324
rect 18062 4380 18126 4384
rect 18062 4324 18066 4380
rect 18066 4324 18122 4380
rect 18122 4324 18126 4380
rect 18062 4320 18126 4324
rect 24791 4380 24855 4384
rect 24791 4324 24795 4380
rect 24795 4324 24851 4380
rect 24851 4324 24855 4380
rect 24791 4320 24855 4324
rect 24871 4380 24935 4384
rect 24871 4324 24875 4380
rect 24875 4324 24931 4380
rect 24931 4324 24935 4380
rect 24871 4320 24935 4324
rect 24951 4380 25015 4384
rect 24951 4324 24955 4380
rect 24955 4324 25011 4380
rect 25011 4324 25015 4380
rect 24951 4320 25015 4324
rect 25031 4380 25095 4384
rect 25031 4324 25035 4380
rect 25035 4324 25091 4380
rect 25091 4324 25095 4380
rect 25031 4320 25095 4324
rect 7368 3836 7432 3840
rect 7368 3780 7372 3836
rect 7372 3780 7428 3836
rect 7428 3780 7432 3836
rect 7368 3776 7432 3780
rect 7448 3836 7512 3840
rect 7448 3780 7452 3836
rect 7452 3780 7508 3836
rect 7508 3780 7512 3836
rect 7448 3776 7512 3780
rect 7528 3836 7592 3840
rect 7528 3780 7532 3836
rect 7532 3780 7588 3836
rect 7588 3780 7592 3836
rect 7528 3776 7592 3780
rect 7608 3836 7672 3840
rect 7608 3780 7612 3836
rect 7612 3780 7668 3836
rect 7668 3780 7672 3836
rect 7608 3776 7672 3780
rect 14337 3836 14401 3840
rect 14337 3780 14341 3836
rect 14341 3780 14397 3836
rect 14397 3780 14401 3836
rect 14337 3776 14401 3780
rect 14417 3836 14481 3840
rect 14417 3780 14421 3836
rect 14421 3780 14477 3836
rect 14477 3780 14481 3836
rect 14417 3776 14481 3780
rect 14497 3836 14561 3840
rect 14497 3780 14501 3836
rect 14501 3780 14557 3836
rect 14557 3780 14561 3836
rect 14497 3776 14561 3780
rect 14577 3836 14641 3840
rect 14577 3780 14581 3836
rect 14581 3780 14637 3836
rect 14637 3780 14641 3836
rect 14577 3776 14641 3780
rect 21306 3836 21370 3840
rect 21306 3780 21310 3836
rect 21310 3780 21366 3836
rect 21366 3780 21370 3836
rect 21306 3776 21370 3780
rect 21386 3836 21450 3840
rect 21386 3780 21390 3836
rect 21390 3780 21446 3836
rect 21446 3780 21450 3836
rect 21386 3776 21450 3780
rect 21466 3836 21530 3840
rect 21466 3780 21470 3836
rect 21470 3780 21526 3836
rect 21526 3780 21530 3836
rect 21466 3776 21530 3780
rect 21546 3836 21610 3840
rect 21546 3780 21550 3836
rect 21550 3780 21606 3836
rect 21606 3780 21610 3836
rect 21546 3776 21610 3780
rect 28275 3836 28339 3840
rect 28275 3780 28279 3836
rect 28279 3780 28335 3836
rect 28335 3780 28339 3836
rect 28275 3776 28339 3780
rect 28355 3836 28419 3840
rect 28355 3780 28359 3836
rect 28359 3780 28415 3836
rect 28415 3780 28419 3836
rect 28355 3776 28419 3780
rect 28435 3836 28499 3840
rect 28435 3780 28439 3836
rect 28439 3780 28495 3836
rect 28495 3780 28499 3836
rect 28435 3776 28499 3780
rect 28515 3836 28579 3840
rect 28515 3780 28519 3836
rect 28519 3780 28575 3836
rect 28575 3780 28579 3836
rect 28515 3776 28579 3780
rect 3884 3292 3948 3296
rect 3884 3236 3888 3292
rect 3888 3236 3944 3292
rect 3944 3236 3948 3292
rect 3884 3232 3948 3236
rect 3964 3292 4028 3296
rect 3964 3236 3968 3292
rect 3968 3236 4024 3292
rect 4024 3236 4028 3292
rect 3964 3232 4028 3236
rect 4044 3292 4108 3296
rect 4044 3236 4048 3292
rect 4048 3236 4104 3292
rect 4104 3236 4108 3292
rect 4044 3232 4108 3236
rect 4124 3292 4188 3296
rect 4124 3236 4128 3292
rect 4128 3236 4184 3292
rect 4184 3236 4188 3292
rect 4124 3232 4188 3236
rect 10853 3292 10917 3296
rect 10853 3236 10857 3292
rect 10857 3236 10913 3292
rect 10913 3236 10917 3292
rect 10853 3232 10917 3236
rect 10933 3292 10997 3296
rect 10933 3236 10937 3292
rect 10937 3236 10993 3292
rect 10993 3236 10997 3292
rect 10933 3232 10997 3236
rect 11013 3292 11077 3296
rect 11013 3236 11017 3292
rect 11017 3236 11073 3292
rect 11073 3236 11077 3292
rect 11013 3232 11077 3236
rect 11093 3292 11157 3296
rect 11093 3236 11097 3292
rect 11097 3236 11153 3292
rect 11153 3236 11157 3292
rect 11093 3232 11157 3236
rect 17822 3292 17886 3296
rect 17822 3236 17826 3292
rect 17826 3236 17882 3292
rect 17882 3236 17886 3292
rect 17822 3232 17886 3236
rect 17902 3292 17966 3296
rect 17902 3236 17906 3292
rect 17906 3236 17962 3292
rect 17962 3236 17966 3292
rect 17902 3232 17966 3236
rect 17982 3292 18046 3296
rect 17982 3236 17986 3292
rect 17986 3236 18042 3292
rect 18042 3236 18046 3292
rect 17982 3232 18046 3236
rect 18062 3292 18126 3296
rect 18062 3236 18066 3292
rect 18066 3236 18122 3292
rect 18122 3236 18126 3292
rect 18062 3232 18126 3236
rect 24791 3292 24855 3296
rect 24791 3236 24795 3292
rect 24795 3236 24851 3292
rect 24851 3236 24855 3292
rect 24791 3232 24855 3236
rect 24871 3292 24935 3296
rect 24871 3236 24875 3292
rect 24875 3236 24931 3292
rect 24931 3236 24935 3292
rect 24871 3232 24935 3236
rect 24951 3292 25015 3296
rect 24951 3236 24955 3292
rect 24955 3236 25011 3292
rect 25011 3236 25015 3292
rect 24951 3232 25015 3236
rect 25031 3292 25095 3296
rect 25031 3236 25035 3292
rect 25035 3236 25091 3292
rect 25091 3236 25095 3292
rect 25031 3232 25095 3236
rect 7368 2748 7432 2752
rect 7368 2692 7372 2748
rect 7372 2692 7428 2748
rect 7428 2692 7432 2748
rect 7368 2688 7432 2692
rect 7448 2748 7512 2752
rect 7448 2692 7452 2748
rect 7452 2692 7508 2748
rect 7508 2692 7512 2748
rect 7448 2688 7512 2692
rect 7528 2748 7592 2752
rect 7528 2692 7532 2748
rect 7532 2692 7588 2748
rect 7588 2692 7592 2748
rect 7528 2688 7592 2692
rect 7608 2748 7672 2752
rect 7608 2692 7612 2748
rect 7612 2692 7668 2748
rect 7668 2692 7672 2748
rect 7608 2688 7672 2692
rect 14337 2748 14401 2752
rect 14337 2692 14341 2748
rect 14341 2692 14397 2748
rect 14397 2692 14401 2748
rect 14337 2688 14401 2692
rect 14417 2748 14481 2752
rect 14417 2692 14421 2748
rect 14421 2692 14477 2748
rect 14477 2692 14481 2748
rect 14417 2688 14481 2692
rect 14497 2748 14561 2752
rect 14497 2692 14501 2748
rect 14501 2692 14557 2748
rect 14557 2692 14561 2748
rect 14497 2688 14561 2692
rect 14577 2748 14641 2752
rect 14577 2692 14581 2748
rect 14581 2692 14637 2748
rect 14637 2692 14641 2748
rect 14577 2688 14641 2692
rect 21306 2748 21370 2752
rect 21306 2692 21310 2748
rect 21310 2692 21366 2748
rect 21366 2692 21370 2748
rect 21306 2688 21370 2692
rect 21386 2748 21450 2752
rect 21386 2692 21390 2748
rect 21390 2692 21446 2748
rect 21446 2692 21450 2748
rect 21386 2688 21450 2692
rect 21466 2748 21530 2752
rect 21466 2692 21470 2748
rect 21470 2692 21526 2748
rect 21526 2692 21530 2748
rect 21466 2688 21530 2692
rect 21546 2748 21610 2752
rect 21546 2692 21550 2748
rect 21550 2692 21606 2748
rect 21606 2692 21610 2748
rect 21546 2688 21610 2692
rect 28275 2748 28339 2752
rect 28275 2692 28279 2748
rect 28279 2692 28335 2748
rect 28335 2692 28339 2748
rect 28275 2688 28339 2692
rect 28355 2748 28419 2752
rect 28355 2692 28359 2748
rect 28359 2692 28415 2748
rect 28415 2692 28419 2748
rect 28355 2688 28419 2692
rect 28435 2748 28499 2752
rect 28435 2692 28439 2748
rect 28439 2692 28495 2748
rect 28495 2692 28499 2748
rect 28435 2688 28499 2692
rect 28515 2748 28579 2752
rect 28515 2692 28519 2748
rect 28519 2692 28575 2748
rect 28575 2692 28579 2748
rect 28515 2688 28579 2692
rect 3884 2204 3948 2208
rect 3884 2148 3888 2204
rect 3888 2148 3944 2204
rect 3944 2148 3948 2204
rect 3884 2144 3948 2148
rect 3964 2204 4028 2208
rect 3964 2148 3968 2204
rect 3968 2148 4024 2204
rect 4024 2148 4028 2204
rect 3964 2144 4028 2148
rect 4044 2204 4108 2208
rect 4044 2148 4048 2204
rect 4048 2148 4104 2204
rect 4104 2148 4108 2204
rect 4044 2144 4108 2148
rect 4124 2204 4188 2208
rect 4124 2148 4128 2204
rect 4128 2148 4184 2204
rect 4184 2148 4188 2204
rect 4124 2144 4188 2148
rect 10853 2204 10917 2208
rect 10853 2148 10857 2204
rect 10857 2148 10913 2204
rect 10913 2148 10917 2204
rect 10853 2144 10917 2148
rect 10933 2204 10997 2208
rect 10933 2148 10937 2204
rect 10937 2148 10993 2204
rect 10993 2148 10997 2204
rect 10933 2144 10997 2148
rect 11013 2204 11077 2208
rect 11013 2148 11017 2204
rect 11017 2148 11073 2204
rect 11073 2148 11077 2204
rect 11013 2144 11077 2148
rect 11093 2204 11157 2208
rect 11093 2148 11097 2204
rect 11097 2148 11153 2204
rect 11153 2148 11157 2204
rect 11093 2144 11157 2148
rect 17822 2204 17886 2208
rect 17822 2148 17826 2204
rect 17826 2148 17882 2204
rect 17882 2148 17886 2204
rect 17822 2144 17886 2148
rect 17902 2204 17966 2208
rect 17902 2148 17906 2204
rect 17906 2148 17962 2204
rect 17962 2148 17966 2204
rect 17902 2144 17966 2148
rect 17982 2204 18046 2208
rect 17982 2148 17986 2204
rect 17986 2148 18042 2204
rect 18042 2148 18046 2204
rect 17982 2144 18046 2148
rect 18062 2204 18126 2208
rect 18062 2148 18066 2204
rect 18066 2148 18122 2204
rect 18122 2148 18126 2204
rect 18062 2144 18126 2148
rect 24791 2204 24855 2208
rect 24791 2148 24795 2204
rect 24795 2148 24851 2204
rect 24851 2148 24855 2204
rect 24791 2144 24855 2148
rect 24871 2204 24935 2208
rect 24871 2148 24875 2204
rect 24875 2148 24931 2204
rect 24931 2148 24935 2204
rect 24871 2144 24935 2148
rect 24951 2204 25015 2208
rect 24951 2148 24955 2204
rect 24955 2148 25011 2204
rect 25011 2148 25015 2204
rect 24951 2144 25015 2148
rect 25031 2204 25095 2208
rect 25031 2148 25035 2204
rect 25035 2148 25091 2204
rect 25091 2148 25095 2204
rect 25031 2144 25095 2148
rect 7368 1660 7432 1664
rect 7368 1604 7372 1660
rect 7372 1604 7428 1660
rect 7428 1604 7432 1660
rect 7368 1600 7432 1604
rect 7448 1660 7512 1664
rect 7448 1604 7452 1660
rect 7452 1604 7508 1660
rect 7508 1604 7512 1660
rect 7448 1600 7512 1604
rect 7528 1660 7592 1664
rect 7528 1604 7532 1660
rect 7532 1604 7588 1660
rect 7588 1604 7592 1660
rect 7528 1600 7592 1604
rect 7608 1660 7672 1664
rect 7608 1604 7612 1660
rect 7612 1604 7668 1660
rect 7668 1604 7672 1660
rect 7608 1600 7672 1604
rect 14337 1660 14401 1664
rect 14337 1604 14341 1660
rect 14341 1604 14397 1660
rect 14397 1604 14401 1660
rect 14337 1600 14401 1604
rect 14417 1660 14481 1664
rect 14417 1604 14421 1660
rect 14421 1604 14477 1660
rect 14477 1604 14481 1660
rect 14417 1600 14481 1604
rect 14497 1660 14561 1664
rect 14497 1604 14501 1660
rect 14501 1604 14557 1660
rect 14557 1604 14561 1660
rect 14497 1600 14561 1604
rect 14577 1660 14641 1664
rect 14577 1604 14581 1660
rect 14581 1604 14637 1660
rect 14637 1604 14641 1660
rect 14577 1600 14641 1604
rect 21306 1660 21370 1664
rect 21306 1604 21310 1660
rect 21310 1604 21366 1660
rect 21366 1604 21370 1660
rect 21306 1600 21370 1604
rect 21386 1660 21450 1664
rect 21386 1604 21390 1660
rect 21390 1604 21446 1660
rect 21446 1604 21450 1660
rect 21386 1600 21450 1604
rect 21466 1660 21530 1664
rect 21466 1604 21470 1660
rect 21470 1604 21526 1660
rect 21526 1604 21530 1660
rect 21466 1600 21530 1604
rect 21546 1660 21610 1664
rect 21546 1604 21550 1660
rect 21550 1604 21606 1660
rect 21606 1604 21610 1660
rect 21546 1600 21610 1604
rect 28275 1660 28339 1664
rect 28275 1604 28279 1660
rect 28279 1604 28335 1660
rect 28335 1604 28339 1660
rect 28275 1600 28339 1604
rect 28355 1660 28419 1664
rect 28355 1604 28359 1660
rect 28359 1604 28415 1660
rect 28415 1604 28419 1660
rect 28355 1600 28419 1604
rect 28435 1660 28499 1664
rect 28435 1604 28439 1660
rect 28439 1604 28495 1660
rect 28495 1604 28499 1660
rect 28435 1600 28499 1604
rect 28515 1660 28579 1664
rect 28515 1604 28519 1660
rect 28519 1604 28575 1660
rect 28575 1604 28579 1660
rect 28515 1600 28579 1604
rect 3884 1116 3948 1120
rect 3884 1060 3888 1116
rect 3888 1060 3944 1116
rect 3944 1060 3948 1116
rect 3884 1056 3948 1060
rect 3964 1116 4028 1120
rect 3964 1060 3968 1116
rect 3968 1060 4024 1116
rect 4024 1060 4028 1116
rect 3964 1056 4028 1060
rect 4044 1116 4108 1120
rect 4044 1060 4048 1116
rect 4048 1060 4104 1116
rect 4104 1060 4108 1116
rect 4044 1056 4108 1060
rect 4124 1116 4188 1120
rect 4124 1060 4128 1116
rect 4128 1060 4184 1116
rect 4184 1060 4188 1116
rect 4124 1056 4188 1060
rect 10853 1116 10917 1120
rect 10853 1060 10857 1116
rect 10857 1060 10913 1116
rect 10913 1060 10917 1116
rect 10853 1056 10917 1060
rect 10933 1116 10997 1120
rect 10933 1060 10937 1116
rect 10937 1060 10993 1116
rect 10993 1060 10997 1116
rect 10933 1056 10997 1060
rect 11013 1116 11077 1120
rect 11013 1060 11017 1116
rect 11017 1060 11073 1116
rect 11073 1060 11077 1116
rect 11013 1056 11077 1060
rect 11093 1116 11157 1120
rect 11093 1060 11097 1116
rect 11097 1060 11153 1116
rect 11153 1060 11157 1116
rect 11093 1056 11157 1060
rect 17822 1116 17886 1120
rect 17822 1060 17826 1116
rect 17826 1060 17882 1116
rect 17882 1060 17886 1116
rect 17822 1056 17886 1060
rect 17902 1116 17966 1120
rect 17902 1060 17906 1116
rect 17906 1060 17962 1116
rect 17962 1060 17966 1116
rect 17902 1056 17966 1060
rect 17982 1116 18046 1120
rect 17982 1060 17986 1116
rect 17986 1060 18042 1116
rect 18042 1060 18046 1116
rect 17982 1056 18046 1060
rect 18062 1116 18126 1120
rect 18062 1060 18066 1116
rect 18066 1060 18122 1116
rect 18122 1060 18126 1116
rect 18062 1056 18126 1060
rect 24791 1116 24855 1120
rect 24791 1060 24795 1116
rect 24795 1060 24851 1116
rect 24851 1060 24855 1116
rect 24791 1056 24855 1060
rect 24871 1116 24935 1120
rect 24871 1060 24875 1116
rect 24875 1060 24931 1116
rect 24931 1060 24935 1116
rect 24871 1056 24935 1060
rect 24951 1116 25015 1120
rect 24951 1060 24955 1116
rect 24955 1060 25011 1116
rect 25011 1060 25015 1116
rect 24951 1056 25015 1060
rect 25031 1116 25095 1120
rect 25031 1060 25035 1116
rect 25035 1060 25091 1116
rect 25091 1060 25095 1116
rect 25031 1056 25095 1060
rect 7368 572 7432 576
rect 7368 516 7372 572
rect 7372 516 7428 572
rect 7428 516 7432 572
rect 7368 512 7432 516
rect 7448 572 7512 576
rect 7448 516 7452 572
rect 7452 516 7508 572
rect 7508 516 7512 572
rect 7448 512 7512 516
rect 7528 572 7592 576
rect 7528 516 7532 572
rect 7532 516 7588 572
rect 7588 516 7592 572
rect 7528 512 7592 516
rect 7608 572 7672 576
rect 7608 516 7612 572
rect 7612 516 7668 572
rect 7668 516 7672 572
rect 7608 512 7672 516
rect 14337 572 14401 576
rect 14337 516 14341 572
rect 14341 516 14397 572
rect 14397 516 14401 572
rect 14337 512 14401 516
rect 14417 572 14481 576
rect 14417 516 14421 572
rect 14421 516 14477 572
rect 14477 516 14481 572
rect 14417 512 14481 516
rect 14497 572 14561 576
rect 14497 516 14501 572
rect 14501 516 14557 572
rect 14557 516 14561 572
rect 14497 512 14561 516
rect 14577 572 14641 576
rect 14577 516 14581 572
rect 14581 516 14637 572
rect 14637 516 14641 572
rect 14577 512 14641 516
rect 21306 572 21370 576
rect 21306 516 21310 572
rect 21310 516 21366 572
rect 21366 516 21370 572
rect 21306 512 21370 516
rect 21386 572 21450 576
rect 21386 516 21390 572
rect 21390 516 21446 572
rect 21446 516 21450 572
rect 21386 512 21450 516
rect 21466 572 21530 576
rect 21466 516 21470 572
rect 21470 516 21526 572
rect 21526 516 21530 572
rect 21466 512 21530 516
rect 21546 572 21610 576
rect 21546 516 21550 572
rect 21550 516 21606 572
rect 21606 516 21610 572
rect 21546 512 21610 516
rect 28275 572 28339 576
rect 28275 516 28279 572
rect 28279 516 28335 572
rect 28335 516 28339 572
rect 28275 512 28339 516
rect 28355 572 28419 576
rect 28355 516 28359 572
rect 28359 516 28415 572
rect 28415 516 28419 572
rect 28355 512 28419 516
rect 28435 572 28499 576
rect 28435 516 28439 572
rect 28439 516 28495 572
rect 28495 516 28499 572
rect 28435 512 28499 516
rect 28515 572 28579 576
rect 28515 516 28519 572
rect 28519 516 28575 572
rect 28575 516 28579 572
rect 28515 512 28579 516
<< metal4 >>
rect 3876 28320 4196 28336
rect 3876 28256 3884 28320
rect 3948 28256 3964 28320
rect 4028 28256 4044 28320
rect 4108 28256 4124 28320
rect 4188 28256 4196 28320
rect 3876 27232 4196 28256
rect 3876 27168 3884 27232
rect 3948 27168 3964 27232
rect 4028 27168 4044 27232
rect 4108 27168 4124 27232
rect 4188 27168 4196 27232
rect 3876 26144 4196 27168
rect 3876 26080 3884 26144
rect 3948 26080 3964 26144
rect 4028 26080 4044 26144
rect 4108 26080 4124 26144
rect 4188 26080 4196 26144
rect 3876 25056 4196 26080
rect 3876 24992 3884 25056
rect 3948 24992 3964 25056
rect 4028 24992 4044 25056
rect 4108 24992 4124 25056
rect 4188 24992 4196 25056
rect 3876 23968 4196 24992
rect 3876 23904 3884 23968
rect 3948 23904 3964 23968
rect 4028 23904 4044 23968
rect 4108 23904 4124 23968
rect 4188 23904 4196 23968
rect 3876 22880 4196 23904
rect 3876 22816 3884 22880
rect 3948 22816 3964 22880
rect 4028 22816 4044 22880
rect 4108 22816 4124 22880
rect 4188 22816 4196 22880
rect 3876 21792 4196 22816
rect 3876 21728 3884 21792
rect 3948 21728 3964 21792
rect 4028 21728 4044 21792
rect 4108 21728 4124 21792
rect 4188 21728 4196 21792
rect 3876 20704 4196 21728
rect 3876 20640 3884 20704
rect 3948 20640 3964 20704
rect 4028 20640 4044 20704
rect 4108 20640 4124 20704
rect 4188 20640 4196 20704
rect 3876 19616 4196 20640
rect 3876 19552 3884 19616
rect 3948 19552 3964 19616
rect 4028 19552 4044 19616
rect 4108 19552 4124 19616
rect 4188 19552 4196 19616
rect 3876 18528 4196 19552
rect 3876 18464 3884 18528
rect 3948 18464 3964 18528
rect 4028 18464 4044 18528
rect 4108 18464 4124 18528
rect 4188 18464 4196 18528
rect 3876 17440 4196 18464
rect 3876 17376 3884 17440
rect 3948 17376 3964 17440
rect 4028 17376 4044 17440
rect 4108 17376 4124 17440
rect 4188 17376 4196 17440
rect 3876 16352 4196 17376
rect 3876 16288 3884 16352
rect 3948 16288 3964 16352
rect 4028 16288 4044 16352
rect 4108 16288 4124 16352
rect 4188 16288 4196 16352
rect 3876 15264 4196 16288
rect 3876 15200 3884 15264
rect 3948 15200 3964 15264
rect 4028 15200 4044 15264
rect 4108 15200 4124 15264
rect 4188 15200 4196 15264
rect 3876 14176 4196 15200
rect 3876 14112 3884 14176
rect 3948 14112 3964 14176
rect 4028 14112 4044 14176
rect 4108 14112 4124 14176
rect 4188 14112 4196 14176
rect 3876 13088 4196 14112
rect 3876 13024 3884 13088
rect 3948 13024 3964 13088
rect 4028 13024 4044 13088
rect 4108 13024 4124 13088
rect 4188 13024 4196 13088
rect 3876 12000 4196 13024
rect 3876 11936 3884 12000
rect 3948 11936 3964 12000
rect 4028 11936 4044 12000
rect 4108 11936 4124 12000
rect 4188 11936 4196 12000
rect 3876 10912 4196 11936
rect 3876 10848 3884 10912
rect 3948 10848 3964 10912
rect 4028 10848 4044 10912
rect 4108 10848 4124 10912
rect 4188 10848 4196 10912
rect 3876 9824 4196 10848
rect 3876 9760 3884 9824
rect 3948 9760 3964 9824
rect 4028 9760 4044 9824
rect 4108 9760 4124 9824
rect 4188 9760 4196 9824
rect 3876 8736 4196 9760
rect 3876 8672 3884 8736
rect 3948 8672 3964 8736
rect 4028 8672 4044 8736
rect 4108 8672 4124 8736
rect 4188 8672 4196 8736
rect 3876 7648 4196 8672
rect 3876 7584 3884 7648
rect 3948 7584 3964 7648
rect 4028 7584 4044 7648
rect 4108 7584 4124 7648
rect 4188 7584 4196 7648
rect 3876 6560 4196 7584
rect 3876 6496 3884 6560
rect 3948 6496 3964 6560
rect 4028 6496 4044 6560
rect 4108 6496 4124 6560
rect 4188 6496 4196 6560
rect 3876 5472 4196 6496
rect 3876 5408 3884 5472
rect 3948 5408 3964 5472
rect 4028 5408 4044 5472
rect 4108 5408 4124 5472
rect 4188 5408 4196 5472
rect 3876 4384 4196 5408
rect 3876 4320 3884 4384
rect 3948 4320 3964 4384
rect 4028 4320 4044 4384
rect 4108 4320 4124 4384
rect 4188 4320 4196 4384
rect 3876 3296 4196 4320
rect 3876 3232 3884 3296
rect 3948 3232 3964 3296
rect 4028 3232 4044 3296
rect 4108 3232 4124 3296
rect 4188 3232 4196 3296
rect 3876 2208 4196 3232
rect 3876 2144 3884 2208
rect 3948 2144 3964 2208
rect 4028 2144 4044 2208
rect 4108 2144 4124 2208
rect 4188 2144 4196 2208
rect 3876 1120 4196 2144
rect 3876 1056 3884 1120
rect 3948 1056 3964 1120
rect 4028 1056 4044 1120
rect 4108 1056 4124 1120
rect 4188 1056 4196 1120
rect 3876 496 4196 1056
rect 7360 27776 7680 28336
rect 7360 27712 7368 27776
rect 7432 27712 7448 27776
rect 7512 27712 7528 27776
rect 7592 27712 7608 27776
rect 7672 27712 7680 27776
rect 7360 26688 7680 27712
rect 7360 26624 7368 26688
rect 7432 26624 7448 26688
rect 7512 26624 7528 26688
rect 7592 26624 7608 26688
rect 7672 26624 7680 26688
rect 7360 25600 7680 26624
rect 7360 25536 7368 25600
rect 7432 25536 7448 25600
rect 7512 25536 7528 25600
rect 7592 25536 7608 25600
rect 7672 25536 7680 25600
rect 7360 24512 7680 25536
rect 7360 24448 7368 24512
rect 7432 24448 7448 24512
rect 7512 24448 7528 24512
rect 7592 24448 7608 24512
rect 7672 24448 7680 24512
rect 7360 23424 7680 24448
rect 7360 23360 7368 23424
rect 7432 23360 7448 23424
rect 7512 23360 7528 23424
rect 7592 23360 7608 23424
rect 7672 23360 7680 23424
rect 7360 22336 7680 23360
rect 7360 22272 7368 22336
rect 7432 22272 7448 22336
rect 7512 22272 7528 22336
rect 7592 22272 7608 22336
rect 7672 22272 7680 22336
rect 7360 21248 7680 22272
rect 7360 21184 7368 21248
rect 7432 21184 7448 21248
rect 7512 21184 7528 21248
rect 7592 21184 7608 21248
rect 7672 21184 7680 21248
rect 7360 20160 7680 21184
rect 7360 20096 7368 20160
rect 7432 20096 7448 20160
rect 7512 20096 7528 20160
rect 7592 20096 7608 20160
rect 7672 20096 7680 20160
rect 7360 19072 7680 20096
rect 7360 19008 7368 19072
rect 7432 19008 7448 19072
rect 7512 19008 7528 19072
rect 7592 19008 7608 19072
rect 7672 19008 7680 19072
rect 7360 17984 7680 19008
rect 7360 17920 7368 17984
rect 7432 17920 7448 17984
rect 7512 17920 7528 17984
rect 7592 17920 7608 17984
rect 7672 17920 7680 17984
rect 7360 16896 7680 17920
rect 7360 16832 7368 16896
rect 7432 16832 7448 16896
rect 7512 16832 7528 16896
rect 7592 16832 7608 16896
rect 7672 16832 7680 16896
rect 7360 15808 7680 16832
rect 7360 15744 7368 15808
rect 7432 15744 7448 15808
rect 7512 15744 7528 15808
rect 7592 15744 7608 15808
rect 7672 15744 7680 15808
rect 7360 14720 7680 15744
rect 7360 14656 7368 14720
rect 7432 14656 7448 14720
rect 7512 14656 7528 14720
rect 7592 14656 7608 14720
rect 7672 14656 7680 14720
rect 7360 13632 7680 14656
rect 7360 13568 7368 13632
rect 7432 13568 7448 13632
rect 7512 13568 7528 13632
rect 7592 13568 7608 13632
rect 7672 13568 7680 13632
rect 7360 12544 7680 13568
rect 7360 12480 7368 12544
rect 7432 12480 7448 12544
rect 7512 12480 7528 12544
rect 7592 12480 7608 12544
rect 7672 12480 7680 12544
rect 7360 11456 7680 12480
rect 7360 11392 7368 11456
rect 7432 11392 7448 11456
rect 7512 11392 7528 11456
rect 7592 11392 7608 11456
rect 7672 11392 7680 11456
rect 7360 10368 7680 11392
rect 7360 10304 7368 10368
rect 7432 10304 7448 10368
rect 7512 10304 7528 10368
rect 7592 10304 7608 10368
rect 7672 10304 7680 10368
rect 7360 9280 7680 10304
rect 7360 9216 7368 9280
rect 7432 9216 7448 9280
rect 7512 9216 7528 9280
rect 7592 9216 7608 9280
rect 7672 9216 7680 9280
rect 7360 8192 7680 9216
rect 7360 8128 7368 8192
rect 7432 8128 7448 8192
rect 7512 8128 7528 8192
rect 7592 8128 7608 8192
rect 7672 8128 7680 8192
rect 7360 7104 7680 8128
rect 7360 7040 7368 7104
rect 7432 7040 7448 7104
rect 7512 7040 7528 7104
rect 7592 7040 7608 7104
rect 7672 7040 7680 7104
rect 7360 6016 7680 7040
rect 7360 5952 7368 6016
rect 7432 5952 7448 6016
rect 7512 5952 7528 6016
rect 7592 5952 7608 6016
rect 7672 5952 7680 6016
rect 7360 4928 7680 5952
rect 7360 4864 7368 4928
rect 7432 4864 7448 4928
rect 7512 4864 7528 4928
rect 7592 4864 7608 4928
rect 7672 4864 7680 4928
rect 7360 3840 7680 4864
rect 7360 3776 7368 3840
rect 7432 3776 7448 3840
rect 7512 3776 7528 3840
rect 7592 3776 7608 3840
rect 7672 3776 7680 3840
rect 7360 2752 7680 3776
rect 7360 2688 7368 2752
rect 7432 2688 7448 2752
rect 7512 2688 7528 2752
rect 7592 2688 7608 2752
rect 7672 2688 7680 2752
rect 7360 1664 7680 2688
rect 7360 1600 7368 1664
rect 7432 1600 7448 1664
rect 7512 1600 7528 1664
rect 7592 1600 7608 1664
rect 7672 1600 7680 1664
rect 7360 576 7680 1600
rect 7360 512 7368 576
rect 7432 512 7448 576
rect 7512 512 7528 576
rect 7592 512 7608 576
rect 7672 512 7680 576
rect 7360 496 7680 512
rect 10845 28320 11165 28336
rect 10845 28256 10853 28320
rect 10917 28256 10933 28320
rect 10997 28256 11013 28320
rect 11077 28256 11093 28320
rect 11157 28256 11165 28320
rect 10845 27232 11165 28256
rect 10845 27168 10853 27232
rect 10917 27168 10933 27232
rect 10997 27168 11013 27232
rect 11077 27168 11093 27232
rect 11157 27168 11165 27232
rect 10845 26144 11165 27168
rect 10845 26080 10853 26144
rect 10917 26080 10933 26144
rect 10997 26080 11013 26144
rect 11077 26080 11093 26144
rect 11157 26080 11165 26144
rect 10845 25056 11165 26080
rect 10845 24992 10853 25056
rect 10917 24992 10933 25056
rect 10997 24992 11013 25056
rect 11077 24992 11093 25056
rect 11157 24992 11165 25056
rect 10845 23968 11165 24992
rect 10845 23904 10853 23968
rect 10917 23904 10933 23968
rect 10997 23904 11013 23968
rect 11077 23904 11093 23968
rect 11157 23904 11165 23968
rect 10845 22880 11165 23904
rect 10845 22816 10853 22880
rect 10917 22816 10933 22880
rect 10997 22816 11013 22880
rect 11077 22816 11093 22880
rect 11157 22816 11165 22880
rect 10845 21792 11165 22816
rect 10845 21728 10853 21792
rect 10917 21728 10933 21792
rect 10997 21728 11013 21792
rect 11077 21728 11093 21792
rect 11157 21728 11165 21792
rect 10845 20704 11165 21728
rect 14329 27776 14649 28336
rect 14329 27712 14337 27776
rect 14401 27712 14417 27776
rect 14481 27712 14497 27776
rect 14561 27712 14577 27776
rect 14641 27712 14649 27776
rect 14329 26688 14649 27712
rect 14329 26624 14337 26688
rect 14401 26624 14417 26688
rect 14481 26624 14497 26688
rect 14561 26624 14577 26688
rect 14641 26624 14649 26688
rect 14329 25600 14649 26624
rect 14329 25536 14337 25600
rect 14401 25536 14417 25600
rect 14481 25536 14497 25600
rect 14561 25536 14577 25600
rect 14641 25536 14649 25600
rect 14329 24512 14649 25536
rect 14329 24448 14337 24512
rect 14401 24448 14417 24512
rect 14481 24448 14497 24512
rect 14561 24448 14577 24512
rect 14641 24448 14649 24512
rect 14329 23424 14649 24448
rect 14329 23360 14337 23424
rect 14401 23360 14417 23424
rect 14481 23360 14497 23424
rect 14561 23360 14577 23424
rect 14641 23360 14649 23424
rect 14329 22336 14649 23360
rect 14329 22272 14337 22336
rect 14401 22272 14417 22336
rect 14481 22272 14497 22336
rect 14561 22272 14577 22336
rect 14641 22272 14649 22336
rect 14329 21248 14649 22272
rect 14329 21184 14337 21248
rect 14401 21184 14417 21248
rect 14481 21184 14497 21248
rect 14561 21184 14577 21248
rect 14641 21184 14649 21248
rect 13491 20772 13557 20773
rect 13491 20708 13492 20772
rect 13556 20708 13557 20772
rect 13491 20707 13557 20708
rect 10845 20640 10853 20704
rect 10917 20640 10933 20704
rect 10997 20640 11013 20704
rect 11077 20640 11093 20704
rect 11157 20640 11165 20704
rect 10845 19616 11165 20640
rect 10845 19552 10853 19616
rect 10917 19552 10933 19616
rect 10997 19552 11013 19616
rect 11077 19552 11093 19616
rect 11157 19552 11165 19616
rect 10845 18528 11165 19552
rect 10845 18464 10853 18528
rect 10917 18464 10933 18528
rect 10997 18464 11013 18528
rect 11077 18464 11093 18528
rect 11157 18464 11165 18528
rect 10845 17440 11165 18464
rect 10845 17376 10853 17440
rect 10917 17376 10933 17440
rect 10997 17376 11013 17440
rect 11077 17376 11093 17440
rect 11157 17376 11165 17440
rect 10845 16352 11165 17376
rect 13494 16421 13554 20707
rect 14329 20160 14649 21184
rect 14329 20096 14337 20160
rect 14401 20096 14417 20160
rect 14481 20096 14497 20160
rect 14561 20096 14577 20160
rect 14641 20096 14649 20160
rect 14329 19072 14649 20096
rect 14329 19008 14337 19072
rect 14401 19008 14417 19072
rect 14481 19008 14497 19072
rect 14561 19008 14577 19072
rect 14641 19008 14649 19072
rect 14329 17984 14649 19008
rect 14329 17920 14337 17984
rect 14401 17920 14417 17984
rect 14481 17920 14497 17984
rect 14561 17920 14577 17984
rect 14641 17920 14649 17984
rect 14329 16896 14649 17920
rect 14329 16832 14337 16896
rect 14401 16832 14417 16896
rect 14481 16832 14497 16896
rect 14561 16832 14577 16896
rect 14641 16832 14649 16896
rect 13491 16420 13557 16421
rect 13491 16356 13492 16420
rect 13556 16356 13557 16420
rect 13491 16355 13557 16356
rect 10845 16288 10853 16352
rect 10917 16288 10933 16352
rect 10997 16288 11013 16352
rect 11077 16288 11093 16352
rect 11157 16288 11165 16352
rect 10845 15264 11165 16288
rect 10845 15200 10853 15264
rect 10917 15200 10933 15264
rect 10997 15200 11013 15264
rect 11077 15200 11093 15264
rect 11157 15200 11165 15264
rect 10845 14176 11165 15200
rect 10845 14112 10853 14176
rect 10917 14112 10933 14176
rect 10997 14112 11013 14176
rect 11077 14112 11093 14176
rect 11157 14112 11165 14176
rect 10845 13088 11165 14112
rect 10845 13024 10853 13088
rect 10917 13024 10933 13088
rect 10997 13024 11013 13088
rect 11077 13024 11093 13088
rect 11157 13024 11165 13088
rect 10845 12000 11165 13024
rect 10845 11936 10853 12000
rect 10917 11936 10933 12000
rect 10997 11936 11013 12000
rect 11077 11936 11093 12000
rect 11157 11936 11165 12000
rect 10845 10912 11165 11936
rect 10845 10848 10853 10912
rect 10917 10848 10933 10912
rect 10997 10848 11013 10912
rect 11077 10848 11093 10912
rect 11157 10848 11165 10912
rect 10845 9824 11165 10848
rect 10845 9760 10853 9824
rect 10917 9760 10933 9824
rect 10997 9760 11013 9824
rect 11077 9760 11093 9824
rect 11157 9760 11165 9824
rect 10845 8736 11165 9760
rect 10845 8672 10853 8736
rect 10917 8672 10933 8736
rect 10997 8672 11013 8736
rect 11077 8672 11093 8736
rect 11157 8672 11165 8736
rect 10845 7648 11165 8672
rect 10845 7584 10853 7648
rect 10917 7584 10933 7648
rect 10997 7584 11013 7648
rect 11077 7584 11093 7648
rect 11157 7584 11165 7648
rect 10845 6560 11165 7584
rect 10845 6496 10853 6560
rect 10917 6496 10933 6560
rect 10997 6496 11013 6560
rect 11077 6496 11093 6560
rect 11157 6496 11165 6560
rect 10845 5472 11165 6496
rect 10845 5408 10853 5472
rect 10917 5408 10933 5472
rect 10997 5408 11013 5472
rect 11077 5408 11093 5472
rect 11157 5408 11165 5472
rect 10845 4384 11165 5408
rect 10845 4320 10853 4384
rect 10917 4320 10933 4384
rect 10997 4320 11013 4384
rect 11077 4320 11093 4384
rect 11157 4320 11165 4384
rect 10845 3296 11165 4320
rect 10845 3232 10853 3296
rect 10917 3232 10933 3296
rect 10997 3232 11013 3296
rect 11077 3232 11093 3296
rect 11157 3232 11165 3296
rect 10845 2208 11165 3232
rect 10845 2144 10853 2208
rect 10917 2144 10933 2208
rect 10997 2144 11013 2208
rect 11077 2144 11093 2208
rect 11157 2144 11165 2208
rect 10845 1120 11165 2144
rect 10845 1056 10853 1120
rect 10917 1056 10933 1120
rect 10997 1056 11013 1120
rect 11077 1056 11093 1120
rect 11157 1056 11165 1120
rect 10845 496 11165 1056
rect 14329 15808 14649 16832
rect 14329 15744 14337 15808
rect 14401 15744 14417 15808
rect 14481 15744 14497 15808
rect 14561 15744 14577 15808
rect 14641 15744 14649 15808
rect 14329 14720 14649 15744
rect 14329 14656 14337 14720
rect 14401 14656 14417 14720
rect 14481 14656 14497 14720
rect 14561 14656 14577 14720
rect 14641 14656 14649 14720
rect 14329 13632 14649 14656
rect 14329 13568 14337 13632
rect 14401 13568 14417 13632
rect 14481 13568 14497 13632
rect 14561 13568 14577 13632
rect 14641 13568 14649 13632
rect 14329 12544 14649 13568
rect 14329 12480 14337 12544
rect 14401 12480 14417 12544
rect 14481 12480 14497 12544
rect 14561 12480 14577 12544
rect 14641 12480 14649 12544
rect 14329 11456 14649 12480
rect 14329 11392 14337 11456
rect 14401 11392 14417 11456
rect 14481 11392 14497 11456
rect 14561 11392 14577 11456
rect 14641 11392 14649 11456
rect 14329 10368 14649 11392
rect 14329 10304 14337 10368
rect 14401 10304 14417 10368
rect 14481 10304 14497 10368
rect 14561 10304 14577 10368
rect 14641 10304 14649 10368
rect 14329 9280 14649 10304
rect 14329 9216 14337 9280
rect 14401 9216 14417 9280
rect 14481 9216 14497 9280
rect 14561 9216 14577 9280
rect 14641 9216 14649 9280
rect 14329 8192 14649 9216
rect 14329 8128 14337 8192
rect 14401 8128 14417 8192
rect 14481 8128 14497 8192
rect 14561 8128 14577 8192
rect 14641 8128 14649 8192
rect 14329 7104 14649 8128
rect 14329 7040 14337 7104
rect 14401 7040 14417 7104
rect 14481 7040 14497 7104
rect 14561 7040 14577 7104
rect 14641 7040 14649 7104
rect 14329 6016 14649 7040
rect 14329 5952 14337 6016
rect 14401 5952 14417 6016
rect 14481 5952 14497 6016
rect 14561 5952 14577 6016
rect 14641 5952 14649 6016
rect 14329 4928 14649 5952
rect 14329 4864 14337 4928
rect 14401 4864 14417 4928
rect 14481 4864 14497 4928
rect 14561 4864 14577 4928
rect 14641 4864 14649 4928
rect 14329 3840 14649 4864
rect 14329 3776 14337 3840
rect 14401 3776 14417 3840
rect 14481 3776 14497 3840
rect 14561 3776 14577 3840
rect 14641 3776 14649 3840
rect 14329 2752 14649 3776
rect 14329 2688 14337 2752
rect 14401 2688 14417 2752
rect 14481 2688 14497 2752
rect 14561 2688 14577 2752
rect 14641 2688 14649 2752
rect 14329 1664 14649 2688
rect 14329 1600 14337 1664
rect 14401 1600 14417 1664
rect 14481 1600 14497 1664
rect 14561 1600 14577 1664
rect 14641 1600 14649 1664
rect 14329 576 14649 1600
rect 14329 512 14337 576
rect 14401 512 14417 576
rect 14481 512 14497 576
rect 14561 512 14577 576
rect 14641 512 14649 576
rect 14329 496 14649 512
rect 17814 28320 18134 28336
rect 17814 28256 17822 28320
rect 17886 28256 17902 28320
rect 17966 28256 17982 28320
rect 18046 28256 18062 28320
rect 18126 28256 18134 28320
rect 17814 27232 18134 28256
rect 17814 27168 17822 27232
rect 17886 27168 17902 27232
rect 17966 27168 17982 27232
rect 18046 27168 18062 27232
rect 18126 27168 18134 27232
rect 17814 26144 18134 27168
rect 17814 26080 17822 26144
rect 17886 26080 17902 26144
rect 17966 26080 17982 26144
rect 18046 26080 18062 26144
rect 18126 26080 18134 26144
rect 17814 25056 18134 26080
rect 17814 24992 17822 25056
rect 17886 24992 17902 25056
rect 17966 24992 17982 25056
rect 18046 24992 18062 25056
rect 18126 24992 18134 25056
rect 17814 23968 18134 24992
rect 17814 23904 17822 23968
rect 17886 23904 17902 23968
rect 17966 23904 17982 23968
rect 18046 23904 18062 23968
rect 18126 23904 18134 23968
rect 17814 22880 18134 23904
rect 17814 22816 17822 22880
rect 17886 22816 17902 22880
rect 17966 22816 17982 22880
rect 18046 22816 18062 22880
rect 18126 22816 18134 22880
rect 17814 21792 18134 22816
rect 17814 21728 17822 21792
rect 17886 21728 17902 21792
rect 17966 21728 17982 21792
rect 18046 21728 18062 21792
rect 18126 21728 18134 21792
rect 17814 20704 18134 21728
rect 17814 20640 17822 20704
rect 17886 20640 17902 20704
rect 17966 20640 17982 20704
rect 18046 20640 18062 20704
rect 18126 20640 18134 20704
rect 17814 19616 18134 20640
rect 17814 19552 17822 19616
rect 17886 19552 17902 19616
rect 17966 19552 17982 19616
rect 18046 19552 18062 19616
rect 18126 19552 18134 19616
rect 17814 18528 18134 19552
rect 17814 18464 17822 18528
rect 17886 18464 17902 18528
rect 17966 18464 17982 18528
rect 18046 18464 18062 18528
rect 18126 18464 18134 18528
rect 17814 17440 18134 18464
rect 17814 17376 17822 17440
rect 17886 17376 17902 17440
rect 17966 17376 17982 17440
rect 18046 17376 18062 17440
rect 18126 17376 18134 17440
rect 17814 16352 18134 17376
rect 17814 16288 17822 16352
rect 17886 16288 17902 16352
rect 17966 16288 17982 16352
rect 18046 16288 18062 16352
rect 18126 16288 18134 16352
rect 17814 15264 18134 16288
rect 17814 15200 17822 15264
rect 17886 15200 17902 15264
rect 17966 15200 17982 15264
rect 18046 15200 18062 15264
rect 18126 15200 18134 15264
rect 17814 14176 18134 15200
rect 17814 14112 17822 14176
rect 17886 14112 17902 14176
rect 17966 14112 17982 14176
rect 18046 14112 18062 14176
rect 18126 14112 18134 14176
rect 17814 13088 18134 14112
rect 17814 13024 17822 13088
rect 17886 13024 17902 13088
rect 17966 13024 17982 13088
rect 18046 13024 18062 13088
rect 18126 13024 18134 13088
rect 17814 12000 18134 13024
rect 17814 11936 17822 12000
rect 17886 11936 17902 12000
rect 17966 11936 17982 12000
rect 18046 11936 18062 12000
rect 18126 11936 18134 12000
rect 17814 10912 18134 11936
rect 17814 10848 17822 10912
rect 17886 10848 17902 10912
rect 17966 10848 17982 10912
rect 18046 10848 18062 10912
rect 18126 10848 18134 10912
rect 17814 9824 18134 10848
rect 17814 9760 17822 9824
rect 17886 9760 17902 9824
rect 17966 9760 17982 9824
rect 18046 9760 18062 9824
rect 18126 9760 18134 9824
rect 17814 8736 18134 9760
rect 17814 8672 17822 8736
rect 17886 8672 17902 8736
rect 17966 8672 17982 8736
rect 18046 8672 18062 8736
rect 18126 8672 18134 8736
rect 17814 7648 18134 8672
rect 17814 7584 17822 7648
rect 17886 7584 17902 7648
rect 17966 7584 17982 7648
rect 18046 7584 18062 7648
rect 18126 7584 18134 7648
rect 17814 6560 18134 7584
rect 17814 6496 17822 6560
rect 17886 6496 17902 6560
rect 17966 6496 17982 6560
rect 18046 6496 18062 6560
rect 18126 6496 18134 6560
rect 17814 5472 18134 6496
rect 17814 5408 17822 5472
rect 17886 5408 17902 5472
rect 17966 5408 17982 5472
rect 18046 5408 18062 5472
rect 18126 5408 18134 5472
rect 17814 4384 18134 5408
rect 17814 4320 17822 4384
rect 17886 4320 17902 4384
rect 17966 4320 17982 4384
rect 18046 4320 18062 4384
rect 18126 4320 18134 4384
rect 17814 3296 18134 4320
rect 17814 3232 17822 3296
rect 17886 3232 17902 3296
rect 17966 3232 17982 3296
rect 18046 3232 18062 3296
rect 18126 3232 18134 3296
rect 17814 2208 18134 3232
rect 17814 2144 17822 2208
rect 17886 2144 17902 2208
rect 17966 2144 17982 2208
rect 18046 2144 18062 2208
rect 18126 2144 18134 2208
rect 17814 1120 18134 2144
rect 17814 1056 17822 1120
rect 17886 1056 17902 1120
rect 17966 1056 17982 1120
rect 18046 1056 18062 1120
rect 18126 1056 18134 1120
rect 17814 496 18134 1056
rect 21298 27776 21618 28336
rect 21298 27712 21306 27776
rect 21370 27712 21386 27776
rect 21450 27712 21466 27776
rect 21530 27712 21546 27776
rect 21610 27712 21618 27776
rect 21298 26688 21618 27712
rect 21298 26624 21306 26688
rect 21370 26624 21386 26688
rect 21450 26624 21466 26688
rect 21530 26624 21546 26688
rect 21610 26624 21618 26688
rect 21298 25600 21618 26624
rect 21298 25536 21306 25600
rect 21370 25536 21386 25600
rect 21450 25536 21466 25600
rect 21530 25536 21546 25600
rect 21610 25536 21618 25600
rect 21298 24512 21618 25536
rect 21298 24448 21306 24512
rect 21370 24448 21386 24512
rect 21450 24448 21466 24512
rect 21530 24448 21546 24512
rect 21610 24448 21618 24512
rect 21298 23424 21618 24448
rect 21298 23360 21306 23424
rect 21370 23360 21386 23424
rect 21450 23360 21466 23424
rect 21530 23360 21546 23424
rect 21610 23360 21618 23424
rect 21298 22336 21618 23360
rect 21298 22272 21306 22336
rect 21370 22272 21386 22336
rect 21450 22272 21466 22336
rect 21530 22272 21546 22336
rect 21610 22272 21618 22336
rect 21298 21248 21618 22272
rect 21298 21184 21306 21248
rect 21370 21184 21386 21248
rect 21450 21184 21466 21248
rect 21530 21184 21546 21248
rect 21610 21184 21618 21248
rect 21298 20160 21618 21184
rect 21298 20096 21306 20160
rect 21370 20096 21386 20160
rect 21450 20096 21466 20160
rect 21530 20096 21546 20160
rect 21610 20096 21618 20160
rect 21298 19072 21618 20096
rect 21298 19008 21306 19072
rect 21370 19008 21386 19072
rect 21450 19008 21466 19072
rect 21530 19008 21546 19072
rect 21610 19008 21618 19072
rect 21298 17984 21618 19008
rect 21298 17920 21306 17984
rect 21370 17920 21386 17984
rect 21450 17920 21466 17984
rect 21530 17920 21546 17984
rect 21610 17920 21618 17984
rect 21298 16896 21618 17920
rect 21298 16832 21306 16896
rect 21370 16832 21386 16896
rect 21450 16832 21466 16896
rect 21530 16832 21546 16896
rect 21610 16832 21618 16896
rect 21298 15808 21618 16832
rect 21298 15744 21306 15808
rect 21370 15744 21386 15808
rect 21450 15744 21466 15808
rect 21530 15744 21546 15808
rect 21610 15744 21618 15808
rect 21298 14720 21618 15744
rect 21298 14656 21306 14720
rect 21370 14656 21386 14720
rect 21450 14656 21466 14720
rect 21530 14656 21546 14720
rect 21610 14656 21618 14720
rect 21298 13632 21618 14656
rect 21298 13568 21306 13632
rect 21370 13568 21386 13632
rect 21450 13568 21466 13632
rect 21530 13568 21546 13632
rect 21610 13568 21618 13632
rect 21298 12544 21618 13568
rect 21298 12480 21306 12544
rect 21370 12480 21386 12544
rect 21450 12480 21466 12544
rect 21530 12480 21546 12544
rect 21610 12480 21618 12544
rect 21298 11456 21618 12480
rect 21298 11392 21306 11456
rect 21370 11392 21386 11456
rect 21450 11392 21466 11456
rect 21530 11392 21546 11456
rect 21610 11392 21618 11456
rect 21298 10368 21618 11392
rect 21298 10304 21306 10368
rect 21370 10304 21386 10368
rect 21450 10304 21466 10368
rect 21530 10304 21546 10368
rect 21610 10304 21618 10368
rect 21298 9280 21618 10304
rect 21298 9216 21306 9280
rect 21370 9216 21386 9280
rect 21450 9216 21466 9280
rect 21530 9216 21546 9280
rect 21610 9216 21618 9280
rect 21298 8192 21618 9216
rect 21298 8128 21306 8192
rect 21370 8128 21386 8192
rect 21450 8128 21466 8192
rect 21530 8128 21546 8192
rect 21610 8128 21618 8192
rect 21298 7104 21618 8128
rect 21298 7040 21306 7104
rect 21370 7040 21386 7104
rect 21450 7040 21466 7104
rect 21530 7040 21546 7104
rect 21610 7040 21618 7104
rect 21298 6016 21618 7040
rect 21298 5952 21306 6016
rect 21370 5952 21386 6016
rect 21450 5952 21466 6016
rect 21530 5952 21546 6016
rect 21610 5952 21618 6016
rect 21298 4928 21618 5952
rect 21298 4864 21306 4928
rect 21370 4864 21386 4928
rect 21450 4864 21466 4928
rect 21530 4864 21546 4928
rect 21610 4864 21618 4928
rect 21298 3840 21618 4864
rect 21298 3776 21306 3840
rect 21370 3776 21386 3840
rect 21450 3776 21466 3840
rect 21530 3776 21546 3840
rect 21610 3776 21618 3840
rect 21298 2752 21618 3776
rect 21298 2688 21306 2752
rect 21370 2688 21386 2752
rect 21450 2688 21466 2752
rect 21530 2688 21546 2752
rect 21610 2688 21618 2752
rect 21298 1664 21618 2688
rect 21298 1600 21306 1664
rect 21370 1600 21386 1664
rect 21450 1600 21466 1664
rect 21530 1600 21546 1664
rect 21610 1600 21618 1664
rect 21298 576 21618 1600
rect 21298 512 21306 576
rect 21370 512 21386 576
rect 21450 512 21466 576
rect 21530 512 21546 576
rect 21610 512 21618 576
rect 21298 496 21618 512
rect 24783 28320 25103 28336
rect 24783 28256 24791 28320
rect 24855 28256 24871 28320
rect 24935 28256 24951 28320
rect 25015 28256 25031 28320
rect 25095 28256 25103 28320
rect 24783 27232 25103 28256
rect 24783 27168 24791 27232
rect 24855 27168 24871 27232
rect 24935 27168 24951 27232
rect 25015 27168 25031 27232
rect 25095 27168 25103 27232
rect 24783 26144 25103 27168
rect 24783 26080 24791 26144
rect 24855 26080 24871 26144
rect 24935 26080 24951 26144
rect 25015 26080 25031 26144
rect 25095 26080 25103 26144
rect 24783 25056 25103 26080
rect 24783 24992 24791 25056
rect 24855 24992 24871 25056
rect 24935 24992 24951 25056
rect 25015 24992 25031 25056
rect 25095 24992 25103 25056
rect 24783 23968 25103 24992
rect 24783 23904 24791 23968
rect 24855 23904 24871 23968
rect 24935 23904 24951 23968
rect 25015 23904 25031 23968
rect 25095 23904 25103 23968
rect 24783 22880 25103 23904
rect 24783 22816 24791 22880
rect 24855 22816 24871 22880
rect 24935 22816 24951 22880
rect 25015 22816 25031 22880
rect 25095 22816 25103 22880
rect 24783 21792 25103 22816
rect 24783 21728 24791 21792
rect 24855 21728 24871 21792
rect 24935 21728 24951 21792
rect 25015 21728 25031 21792
rect 25095 21728 25103 21792
rect 24783 20704 25103 21728
rect 24783 20640 24791 20704
rect 24855 20640 24871 20704
rect 24935 20640 24951 20704
rect 25015 20640 25031 20704
rect 25095 20640 25103 20704
rect 24783 19616 25103 20640
rect 24783 19552 24791 19616
rect 24855 19552 24871 19616
rect 24935 19552 24951 19616
rect 25015 19552 25031 19616
rect 25095 19552 25103 19616
rect 24783 18528 25103 19552
rect 24783 18464 24791 18528
rect 24855 18464 24871 18528
rect 24935 18464 24951 18528
rect 25015 18464 25031 18528
rect 25095 18464 25103 18528
rect 24783 17440 25103 18464
rect 24783 17376 24791 17440
rect 24855 17376 24871 17440
rect 24935 17376 24951 17440
rect 25015 17376 25031 17440
rect 25095 17376 25103 17440
rect 24783 16352 25103 17376
rect 24783 16288 24791 16352
rect 24855 16288 24871 16352
rect 24935 16288 24951 16352
rect 25015 16288 25031 16352
rect 25095 16288 25103 16352
rect 24783 15264 25103 16288
rect 24783 15200 24791 15264
rect 24855 15200 24871 15264
rect 24935 15200 24951 15264
rect 25015 15200 25031 15264
rect 25095 15200 25103 15264
rect 24783 14176 25103 15200
rect 24783 14112 24791 14176
rect 24855 14112 24871 14176
rect 24935 14112 24951 14176
rect 25015 14112 25031 14176
rect 25095 14112 25103 14176
rect 24783 13088 25103 14112
rect 24783 13024 24791 13088
rect 24855 13024 24871 13088
rect 24935 13024 24951 13088
rect 25015 13024 25031 13088
rect 25095 13024 25103 13088
rect 24783 12000 25103 13024
rect 24783 11936 24791 12000
rect 24855 11936 24871 12000
rect 24935 11936 24951 12000
rect 25015 11936 25031 12000
rect 25095 11936 25103 12000
rect 24783 10912 25103 11936
rect 24783 10848 24791 10912
rect 24855 10848 24871 10912
rect 24935 10848 24951 10912
rect 25015 10848 25031 10912
rect 25095 10848 25103 10912
rect 24783 9824 25103 10848
rect 24783 9760 24791 9824
rect 24855 9760 24871 9824
rect 24935 9760 24951 9824
rect 25015 9760 25031 9824
rect 25095 9760 25103 9824
rect 24783 8736 25103 9760
rect 24783 8672 24791 8736
rect 24855 8672 24871 8736
rect 24935 8672 24951 8736
rect 25015 8672 25031 8736
rect 25095 8672 25103 8736
rect 24783 7648 25103 8672
rect 24783 7584 24791 7648
rect 24855 7584 24871 7648
rect 24935 7584 24951 7648
rect 25015 7584 25031 7648
rect 25095 7584 25103 7648
rect 24783 6560 25103 7584
rect 24783 6496 24791 6560
rect 24855 6496 24871 6560
rect 24935 6496 24951 6560
rect 25015 6496 25031 6560
rect 25095 6496 25103 6560
rect 24783 5472 25103 6496
rect 24783 5408 24791 5472
rect 24855 5408 24871 5472
rect 24935 5408 24951 5472
rect 25015 5408 25031 5472
rect 25095 5408 25103 5472
rect 24783 4384 25103 5408
rect 24783 4320 24791 4384
rect 24855 4320 24871 4384
rect 24935 4320 24951 4384
rect 25015 4320 25031 4384
rect 25095 4320 25103 4384
rect 24783 3296 25103 4320
rect 24783 3232 24791 3296
rect 24855 3232 24871 3296
rect 24935 3232 24951 3296
rect 25015 3232 25031 3296
rect 25095 3232 25103 3296
rect 24783 2208 25103 3232
rect 24783 2144 24791 2208
rect 24855 2144 24871 2208
rect 24935 2144 24951 2208
rect 25015 2144 25031 2208
rect 25095 2144 25103 2208
rect 24783 1120 25103 2144
rect 24783 1056 24791 1120
rect 24855 1056 24871 1120
rect 24935 1056 24951 1120
rect 25015 1056 25031 1120
rect 25095 1056 25103 1120
rect 24783 496 25103 1056
rect 28267 27776 28587 28336
rect 28267 27712 28275 27776
rect 28339 27712 28355 27776
rect 28419 27712 28435 27776
rect 28499 27712 28515 27776
rect 28579 27712 28587 27776
rect 28267 26688 28587 27712
rect 28267 26624 28275 26688
rect 28339 26624 28355 26688
rect 28419 26624 28435 26688
rect 28499 26624 28515 26688
rect 28579 26624 28587 26688
rect 28267 25600 28587 26624
rect 28267 25536 28275 25600
rect 28339 25536 28355 25600
rect 28419 25536 28435 25600
rect 28499 25536 28515 25600
rect 28579 25536 28587 25600
rect 28267 24512 28587 25536
rect 28267 24448 28275 24512
rect 28339 24448 28355 24512
rect 28419 24448 28435 24512
rect 28499 24448 28515 24512
rect 28579 24448 28587 24512
rect 28267 23424 28587 24448
rect 28267 23360 28275 23424
rect 28339 23360 28355 23424
rect 28419 23360 28435 23424
rect 28499 23360 28515 23424
rect 28579 23360 28587 23424
rect 28267 22336 28587 23360
rect 28267 22272 28275 22336
rect 28339 22272 28355 22336
rect 28419 22272 28435 22336
rect 28499 22272 28515 22336
rect 28579 22272 28587 22336
rect 28267 21248 28587 22272
rect 28267 21184 28275 21248
rect 28339 21184 28355 21248
rect 28419 21184 28435 21248
rect 28499 21184 28515 21248
rect 28579 21184 28587 21248
rect 28267 20160 28587 21184
rect 28267 20096 28275 20160
rect 28339 20096 28355 20160
rect 28419 20096 28435 20160
rect 28499 20096 28515 20160
rect 28579 20096 28587 20160
rect 28267 19072 28587 20096
rect 28267 19008 28275 19072
rect 28339 19008 28355 19072
rect 28419 19008 28435 19072
rect 28499 19008 28515 19072
rect 28579 19008 28587 19072
rect 28267 17984 28587 19008
rect 28267 17920 28275 17984
rect 28339 17920 28355 17984
rect 28419 17920 28435 17984
rect 28499 17920 28515 17984
rect 28579 17920 28587 17984
rect 28267 16896 28587 17920
rect 28267 16832 28275 16896
rect 28339 16832 28355 16896
rect 28419 16832 28435 16896
rect 28499 16832 28515 16896
rect 28579 16832 28587 16896
rect 28267 15808 28587 16832
rect 28267 15744 28275 15808
rect 28339 15744 28355 15808
rect 28419 15744 28435 15808
rect 28499 15744 28515 15808
rect 28579 15744 28587 15808
rect 28267 14720 28587 15744
rect 28267 14656 28275 14720
rect 28339 14656 28355 14720
rect 28419 14656 28435 14720
rect 28499 14656 28515 14720
rect 28579 14656 28587 14720
rect 28267 13632 28587 14656
rect 28267 13568 28275 13632
rect 28339 13568 28355 13632
rect 28419 13568 28435 13632
rect 28499 13568 28515 13632
rect 28579 13568 28587 13632
rect 28267 12544 28587 13568
rect 28267 12480 28275 12544
rect 28339 12480 28355 12544
rect 28419 12480 28435 12544
rect 28499 12480 28515 12544
rect 28579 12480 28587 12544
rect 28267 11456 28587 12480
rect 28267 11392 28275 11456
rect 28339 11392 28355 11456
rect 28419 11392 28435 11456
rect 28499 11392 28515 11456
rect 28579 11392 28587 11456
rect 28267 10368 28587 11392
rect 28267 10304 28275 10368
rect 28339 10304 28355 10368
rect 28419 10304 28435 10368
rect 28499 10304 28515 10368
rect 28579 10304 28587 10368
rect 28267 9280 28587 10304
rect 28267 9216 28275 9280
rect 28339 9216 28355 9280
rect 28419 9216 28435 9280
rect 28499 9216 28515 9280
rect 28579 9216 28587 9280
rect 28267 8192 28587 9216
rect 28267 8128 28275 8192
rect 28339 8128 28355 8192
rect 28419 8128 28435 8192
rect 28499 8128 28515 8192
rect 28579 8128 28587 8192
rect 28267 7104 28587 8128
rect 28267 7040 28275 7104
rect 28339 7040 28355 7104
rect 28419 7040 28435 7104
rect 28499 7040 28515 7104
rect 28579 7040 28587 7104
rect 28267 6016 28587 7040
rect 28267 5952 28275 6016
rect 28339 5952 28355 6016
rect 28419 5952 28435 6016
rect 28499 5952 28515 6016
rect 28579 5952 28587 6016
rect 28267 4928 28587 5952
rect 28267 4864 28275 4928
rect 28339 4864 28355 4928
rect 28419 4864 28435 4928
rect 28499 4864 28515 4928
rect 28579 4864 28587 4928
rect 28267 3840 28587 4864
rect 28267 3776 28275 3840
rect 28339 3776 28355 3840
rect 28419 3776 28435 3840
rect 28499 3776 28515 3840
rect 28579 3776 28587 3840
rect 28267 2752 28587 3776
rect 28267 2688 28275 2752
rect 28339 2688 28355 2752
rect 28419 2688 28435 2752
rect 28499 2688 28515 2752
rect 28579 2688 28587 2752
rect 28267 1664 28587 2688
rect 28267 1600 28275 1664
rect 28339 1600 28355 1664
rect 28419 1600 28435 1664
rect 28499 1600 28515 1664
rect 28579 1600 28587 1664
rect 28267 576 28587 1600
rect 28267 512 28275 576
rect 28339 512 28355 576
rect 28419 512 28435 576
rect 28499 512 28515 576
rect 28579 512 28587 576
rect 28267 496 28587 512
use sky130_fd_sc_hd__or3_1  _0463_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13156 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0464_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13800 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0465_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14076 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0466_
timestamp 1704896540
transform -1 0 12972 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0467_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12604 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0468_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13156 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0469_
timestamp 1704896540
transform -1 0 2668 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0470_
timestamp 1704896540
transform -1 0 5060 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0471_
timestamp 1704896540
transform -1 0 4140 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0472_
timestamp 1704896540
transform 1 0 5152 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0473_
timestamp 1704896540
transform -1 0 7176 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0474_
timestamp 1704896540
transform 1 0 6348 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0475_
timestamp 1704896540
transform 1 0 8004 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0476_
timestamp 1704896540
transform -1 0 8740 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _0477_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8004 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0478_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9016 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0479_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16008 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0480_
timestamp 1704896540
transform 1 0 11776 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0481_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12328 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0482_
timestamp 1704896540
transform -1 0 12604 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0483_
timestamp 1704896540
transform -1 0 11868 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0484_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11868 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_1  _0485_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5796 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12972 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0487_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8372 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0488_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9292 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0489_
timestamp 1704896540
transform -1 0 14444 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10580 0 -1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9016 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13064 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0493_
timestamp 1704896540
transform -1 0 10120 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0494_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9660 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0495_
timestamp 1704896540
transform 1 0 11684 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0496_
timestamp 1704896540
transform -1 0 10856 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1704896540
transform -1 0 8464 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0498_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11684 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0499_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10948 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0500_
timestamp 1704896540
transform 1 0 6716 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0501_
timestamp 1704896540
transform -1 0 6992 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _0502_
timestamp 1704896540
transform 1 0 7176 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1704896540
transform -1 0 23368 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504_
timestamp 1704896540
transform -1 0 21160 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1704896540
transform -1 0 20240 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0506_
timestamp 1704896540
transform 1 0 18216 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0507_
timestamp 1704896540
transform -1 0 12972 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0508_
timestamp 1704896540
transform 1 0 12972 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0509_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12880 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0510_
timestamp 1704896540
transform -1 0 12788 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0511_
timestamp 1704896540
transform 1 0 5796 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0512_
timestamp 1704896540
transform 1 0 4140 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0513_
timestamp 1704896540
transform -1 0 9568 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0514_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6992 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0515_
timestamp 1704896540
transform -1 0 6532 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0516_
timestamp 1704896540
transform 1 0 5980 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0517_
timestamp 1704896540
transform 1 0 6532 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0518_
timestamp 1704896540
transform -1 0 7452 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0519_
timestamp 1704896540
transform -1 0 6900 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0520_
timestamp 1704896540
transform 1 0 6900 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0521_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6440 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0522_
timestamp 1704896540
transform 1 0 7912 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0523_
timestamp 1704896540
transform -1 0 12236 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0524_
timestamp 1704896540
transform 1 0 10580 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0525_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11132 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0526_
timestamp 1704896540
transform 1 0 8096 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0527_
timestamp 1704896540
transform 1 0 7820 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0528_
timestamp 1704896540
transform 1 0 8372 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0529_
timestamp 1704896540
transform 1 0 7268 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0530_
timestamp 1704896540
transform 1 0 7544 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0531_
timestamp 1704896540
transform 1 0 9108 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0532_
timestamp 1704896540
transform 1 0 9844 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _0533_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12144 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0534_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7084 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0535_
timestamp 1704896540
transform 1 0 7728 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0536_
timestamp 1704896540
transform 1 0 8556 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0537_
timestamp 1704896540
transform -1 0 6624 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0538_
timestamp 1704896540
transform 1 0 6164 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0539_
timestamp 1704896540
transform 1 0 7360 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0540_
timestamp 1704896540
transform 1 0 7360 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0541_
timestamp 1704896540
transform 1 0 8004 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0542_
timestamp 1704896540
transform 1 0 8740 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0543_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11776 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0544_
timestamp 1704896540
transform 1 0 11224 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0545_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11684 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0546_
timestamp 1704896540
transform -1 0 13156 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0547_
timestamp 1704896540
transform -1 0 7912 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0548_
timestamp 1704896540
transform -1 0 8740 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0549_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8556 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0550_
timestamp 1704896540
transform -1 0 16560 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0551_
timestamp 1704896540
transform 1 0 14260 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0552_
timestamp 1704896540
transform -1 0 15180 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0553_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14352 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0554_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12052 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0555_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12420 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0556_
timestamp 1704896540
transform 1 0 17848 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0557_
timestamp 1704896540
transform -1 0 5520 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _0558_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4416 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0559_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6072 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _0560_
timestamp 1704896540
transform 1 0 6716 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14904 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _0562_
timestamp 1704896540
transform -1 0 14076 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _0563_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14904 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0564_
timestamp 1704896540
transform -1 0 9384 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0565_
timestamp 1704896540
transform 1 0 4324 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0566_
timestamp 1704896540
transform 1 0 8648 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0567_
timestamp 1704896540
transform 1 0 8924 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0568_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9660 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0569_
timestamp 1704896540
transform -1 0 10028 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _0570_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6992 0 1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_1  _0571_
timestamp 1704896540
transform -1 0 13984 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0572_
timestamp 1704896540
transform 1 0 10948 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0573_
timestamp 1704896540
transform 1 0 9844 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0574_
timestamp 1704896540
transform -1 0 10764 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0575_
timestamp 1704896540
transform -1 0 4876 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0576_
timestamp 1704896540
transform -1 0 5152 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0577_
timestamp 1704896540
transform 1 0 4324 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0578_
timestamp 1704896540
transform 1 0 5796 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0579_
timestamp 1704896540
transform -1 0 4140 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0580_
timestamp 1704896540
transform 1 0 3864 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0581_
timestamp 1704896540
transform -1 0 3864 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0582_
timestamp 1704896540
transform 1 0 2760 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0583_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 23920 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0584_
timestamp 1704896540
transform 1 0 3312 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0585_
timestamp 1704896540
transform 1 0 2944 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0586_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12052 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0587_
timestamp 1704896540
transform -1 0 20700 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1704896540
transform 1 0 20608 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _0589_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 20700 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0590_
timestamp 1704896540
transform -1 0 21620 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0591_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21344 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0592_
timestamp 1704896540
transform -1 0 19596 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0593_
timestamp 1704896540
transform 1 0 18032 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0594_
timestamp 1704896540
transform -1 0 18584 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0595_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 21344 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 21620 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0597_
timestamp 1704896540
transform 1 0 21252 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0598_
timestamp 1704896540
transform 1 0 21712 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _0599_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 21344 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0600_
timestamp 1704896540
transform -1 0 22448 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0601_
timestamp 1704896540
transform -1 0 21160 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0602_
timestamp 1704896540
transform 1 0 19964 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _0603_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18768 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0604_
timestamp 1704896540
transform 1 0 18676 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0605_
timestamp 1704896540
transform 1 0 19596 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0606_
timestamp 1704896540
transform 1 0 22356 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _0607_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 22540 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0608_
timestamp 1704896540
transform -1 0 23368 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_2  _0609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21620 0 1 23392
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _0610_
timestamp 1704896540
transform -1 0 22540 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0611_
timestamp 1704896540
transform 1 0 22540 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0612_
timestamp 1704896540
transform -1 0 24472 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0613_
timestamp 1704896540
transform 1 0 23368 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0614_
timestamp 1704896540
transform 1 0 24472 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0615_
timestamp 1704896540
transform 1 0 22356 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0616_
timestamp 1704896540
transform 1 0 22080 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0617_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 22356 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0618_
timestamp 1704896540
transform 1 0 23092 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0619_
timestamp 1704896540
transform 1 0 23276 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0620_
timestamp 1704896540
transform 1 0 24288 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0621_
timestamp 1704896540
transform 1 0 21988 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0622_
timestamp 1704896540
transform 1 0 21252 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0623_
timestamp 1704896540
transform -1 0 21896 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0624_
timestamp 1704896540
transform 1 0 21712 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0625_
timestamp 1704896540
transform 1 0 21804 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0626_
timestamp 1704896540
transform -1 0 23460 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0627_
timestamp 1704896540
transform -1 0 24196 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _0628_
timestamp 1704896540
transform 1 0 22724 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0629_
timestamp 1704896540
transform 1 0 22080 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0630_
timestamp 1704896540
transform 1 0 22448 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0631_
timestamp 1704896540
transform 1 0 22540 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0632_
timestamp 1704896540
transform 1 0 23184 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1704896540
transform -1 0 18952 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0634_
timestamp 1704896540
transform -1 0 22356 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0635_
timestamp 1704896540
transform -1 0 22080 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0636_
timestamp 1704896540
transform 1 0 18584 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1704896540
transform 1 0 18676 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0638_
timestamp 1704896540
transform -1 0 18492 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0639_
timestamp 1704896540
transform -1 0 18584 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0640_
timestamp 1704896540
transform -1 0 21068 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0641_
timestamp 1704896540
transform -1 0 21160 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0642_
timestamp 1704896540
transform 1 0 20240 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0643_
timestamp 1704896540
transform 1 0 21252 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _0644_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 20240 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0645_
timestamp 1704896540
transform 1 0 19872 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0646_
timestamp 1704896540
transform -1 0 19780 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0647_
timestamp 1704896540
transform 1 0 20148 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0648_
timestamp 1704896540
transform -1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _0649_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18860 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0650_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19596 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0651_
timestamp 1704896540
transform 1 0 18308 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0652_
timestamp 1704896540
transform -1 0 19228 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1704896540
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11868 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0655_
timestamp 1704896540
transform 1 0 11316 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0656_
timestamp 1704896540
transform -1 0 20240 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0657_
timestamp 1704896540
transform -1 0 20240 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0658_
timestamp 1704896540
transform 1 0 13708 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0659_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18676 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0660_
timestamp 1704896540
transform 1 0 20240 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0661_
timestamp 1704896540
transform 1 0 20976 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0662_
timestamp 1704896540
transform -1 0 22080 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0663_
timestamp 1704896540
transform -1 0 21528 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0664_
timestamp 1704896540
transform -1 0 20148 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _0665_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 20884 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0666_
timestamp 1704896540
transform 1 0 18860 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0667_
timestamp 1704896540
transform 1 0 19044 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0668_
timestamp 1704896540
transform -1 0 19596 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0669_
timestamp 1704896540
transform 1 0 19688 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0670_
timestamp 1704896540
transform 1 0 20516 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0671_
timestamp 1704896540
transform 1 0 21252 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0672_
timestamp 1704896540
transform -1 0 21712 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0673_
timestamp 1704896540
transform 1 0 17848 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1704896540
transform 1 0 19228 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0675_
timestamp 1704896540
transform 1 0 19596 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0676_
timestamp 1704896540
transform 1 0 18584 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0677_
timestamp 1704896540
transform 1 0 19596 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0678_
timestamp 1704896540
transform 1 0 20240 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0679_
timestamp 1704896540
transform -1 0 20976 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1704896540
transform 1 0 18216 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0681_
timestamp 1704896540
transform 1 0 18676 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0682_
timestamp 1704896540
transform 1 0 18400 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0683_
timestamp 1704896540
transform -1 0 15916 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0684_
timestamp 1704896540
transform 1 0 15180 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0685_
timestamp 1704896540
transform 1 0 16100 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0686_
timestamp 1704896540
transform 1 0 15824 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0687_
timestamp 1704896540
transform 1 0 16744 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0688_
timestamp 1704896540
transform 1 0 17388 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0689_
timestamp 1704896540
transform 1 0 17848 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0690_
timestamp 1704896540
transform -1 0 15088 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0691_
timestamp 1704896540
transform -1 0 14076 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0692_
timestamp 1704896540
transform 1 0 13064 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0693_
timestamp 1704896540
transform 1 0 14260 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0694_
timestamp 1704896540
transform -1 0 11684 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0695_
timestamp 1704896540
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0696_
timestamp 1704896540
transform -1 0 12236 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1704896540
transform -1 0 11684 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0698_
timestamp 1704896540
transform -1 0 13248 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0699_
timestamp 1704896540
transform 1 0 12880 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0700_
timestamp 1704896540
transform 1 0 14076 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0701_
timestamp 1704896540
transform -1 0 13984 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0702_
timestamp 1704896540
transform -1 0 13892 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0703_
timestamp 1704896540
transform -1 0 13984 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0704_
timestamp 1704896540
transform 1 0 11868 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0705_
timestamp 1704896540
transform -1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0706_
timestamp 1704896540
transform -1 0 15364 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0707_
timestamp 1704896540
transform 1 0 14812 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0708_
timestamp 1704896540
transform 1 0 14536 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0709_
timestamp 1704896540
transform 1 0 14996 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0710_
timestamp 1704896540
transform 1 0 15640 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0711_
timestamp 1704896540
transform -1 0 16008 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0712_
timestamp 1704896540
transform -1 0 16468 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1704896540
transform -1 0 4876 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0714_
timestamp 1704896540
transform -1 0 5704 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0715_
timestamp 1704896540
transform 1 0 5796 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0716_
timestamp 1704896540
transform 1 0 2944 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0717_
timestamp 1704896540
transform 1 0 3588 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0718_
timestamp 1704896540
transform -1 0 4968 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0719_
timestamp 1704896540
transform -1 0 2484 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0720_
timestamp 1704896540
transform 1 0 1840 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0721_
timestamp 1704896540
transform 1 0 3956 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _0722_
timestamp 1704896540
transform 1 0 3680 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0723_
timestamp 1704896540
transform 1 0 2024 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0724_
timestamp 1704896540
transform 1 0 2576 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0725_
timestamp 1704896540
transform -1 0 3496 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0726_
timestamp 1704896540
transform 1 0 3588 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0727_
timestamp 1704896540
transform -1 0 4876 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0728_
timestamp 1704896540
transform -1 0 2576 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0729_
timestamp 1704896540
transform 1 0 1932 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0730_
timestamp 1704896540
transform -1 0 5336 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0731_
timestamp 1704896540
transform 1 0 3128 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0732_
timestamp 1704896540
transform 1 0 3220 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0733_
timestamp 1704896540
transform -1 0 4784 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0734_
timestamp 1704896540
transform 1 0 3220 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0735_
timestamp 1704896540
transform 1 0 3680 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0736_
timestamp 1704896540
transform 1 0 7912 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _0737_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4140 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0738_
timestamp 1704896540
transform -1 0 4140 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0739_
timestamp 1704896540
transform 1 0 8740 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0740_
timestamp 1704896540
transform 1 0 6808 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0741_
timestamp 1704896540
transform -1 0 7912 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0742_
timestamp 1704896540
transform 1 0 7912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0743_
timestamp 1704896540
transform -1 0 6440 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0744_
timestamp 1704896540
transform 1 0 5428 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0745_
timestamp 1704896540
transform 1 0 5796 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0746_
timestamp 1704896540
transform 1 0 6256 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0747_
timestamp 1704896540
transform -1 0 7544 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0748_
timestamp 1704896540
transform -1 0 7176 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0749_
timestamp 1704896540
transform -1 0 6900 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0750_
timestamp 1704896540
transform -1 0 8096 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0751_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6716 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0752_
timestamp 1704896540
transform 1 0 6716 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0753_
timestamp 1704896540
transform -1 0 7452 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0754_
timestamp 1704896540
transform 1 0 10488 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0755_
timestamp 1704896540
transform -1 0 10580 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0756_
timestamp 1704896540
transform 1 0 8740 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0757_
timestamp 1704896540
transform 1 0 9752 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0758_
timestamp 1704896540
transform 1 0 7176 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _0759_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9016 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0760_
timestamp 1704896540
transform -1 0 11040 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0761_
timestamp 1704896540
transform 1 0 9660 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0762_
timestamp 1704896540
transform 1 0 10028 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0763_
timestamp 1704896540
transform 1 0 10120 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0764_
timestamp 1704896540
transform 1 0 8464 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0765_
timestamp 1704896540
transform 1 0 8832 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0766_
timestamp 1704896540
transform 1 0 9200 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0767_
timestamp 1704896540
transform 1 0 8464 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0768_
timestamp 1704896540
transform -1 0 8372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0769_
timestamp 1704896540
transform 1 0 10212 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0770_
timestamp 1704896540
transform -1 0 9292 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0771_
timestamp 1704896540
transform 1 0 9476 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0772_
timestamp 1704896540
transform -1 0 10580 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0773_
timestamp 1704896540
transform 1 0 11316 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0774_
timestamp 1704896540
transform 1 0 10580 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0775_
timestamp 1704896540
transform 1 0 10396 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0776_
timestamp 1704896540
transform 1 0 11408 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1704896540
transform 1 0 17204 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0778_
timestamp 1704896540
transform 1 0 16560 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0779_
timestamp 1704896540
transform 1 0 17480 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1704896540
transform -1 0 19688 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0781_
timestamp 1704896540
transform 1 0 16560 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _0782_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17940 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0783_
timestamp 1704896540
transform -1 0 19320 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0784_
timestamp 1704896540
transform -1 0 19136 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0785_
timestamp 1704896540
transform -1 0 18124 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0786_
timestamp 1704896540
transform 1 0 16744 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0787_
timestamp 1704896540
transform 1 0 16192 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0788_
timestamp 1704896540
transform 1 0 15456 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0789_
timestamp 1704896540
transform 1 0 16192 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0790_
timestamp 1704896540
transform -1 0 17572 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0791_
timestamp 1704896540
transform -1 0 17296 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0792_
timestamp 1704896540
transform -1 0 10580 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0793_
timestamp 1704896540
transform 1 0 11592 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0794_
timestamp 1704896540
transform -1 0 11592 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0795_
timestamp 1704896540
transform -1 0 11408 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0796_
timestamp 1704896540
transform 1 0 8372 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0797_
timestamp 1704896540
transform -1 0 9016 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0798_
timestamp 1704896540
transform 1 0 7636 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0799_
timestamp 1704896540
transform -1 0 9660 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0800_
timestamp 1704896540
transform -1 0 9108 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0801_
timestamp 1704896540
transform 1 0 4324 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0802_
timestamp 1704896540
transform 1 0 5428 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0803_
timestamp 1704896540
transform 1 0 4416 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0804_
timestamp 1704896540
transform 1 0 4416 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0805_
timestamp 1704896540
transform 1 0 4784 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0806_
timestamp 1704896540
transform 1 0 4784 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0807_
timestamp 1704896540
transform 1 0 4140 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0808_
timestamp 1704896540
transform -1 0 6992 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _0809_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9200 0 -1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0810_
timestamp 1704896540
transform 1 0 6072 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0811_
timestamp 1704896540
transform 1 0 6532 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _0812_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6072 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _0813_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5796 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0814_
timestamp 1704896540
transform 1 0 6532 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0815_
timestamp 1704896540
transform 1 0 7176 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0816_
timestamp 1704896540
transform -1 0 7176 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0817_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7176 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0818_
timestamp 1704896540
transform 1 0 8280 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1704896540
transform -1 0 7360 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0820_
timestamp 1704896540
transform 1 0 5060 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0821_
timestamp 1704896540
transform -1 0 6532 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0822_
timestamp 1704896540
transform 1 0 6624 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0823_
timestamp 1704896540
transform -1 0 9292 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0824_
timestamp 1704896540
transform 1 0 9292 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0825_
timestamp 1704896540
transform -1 0 9476 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1704896540
transform 1 0 9568 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0827_
timestamp 1704896540
transform 1 0 9660 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0828_
timestamp 1704896540
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0829_
timestamp 1704896540
transform 1 0 12788 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1704896540
transform -1 0 13800 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0831_
timestamp 1704896540
transform -1 0 13616 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0832_
timestamp 1704896540
transform 1 0 12696 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1704896540
transform -1 0 10488 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0834_
timestamp 1704896540
transform 1 0 9660 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0835_
timestamp 1704896540
transform 1 0 9936 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0836_
timestamp 1704896540
transform -1 0 10396 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0837_
timestamp 1704896540
transform -1 0 16008 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0838_
timestamp 1704896540
transform -1 0 15456 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0839_
timestamp 1704896540
transform 1 0 13800 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0840_
timestamp 1704896540
transform 1 0 16192 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0841_
timestamp 1704896540
transform 1 0 15180 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0842_
timestamp 1704896540
transform 1 0 13800 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0843_
timestamp 1704896540
transform 1 0 14996 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0844_
timestamp 1704896540
transform 1 0 15456 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0845_
timestamp 1704896540
transform -1 0 15824 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0846_
timestamp 1704896540
transform 1 0 16744 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0847_
timestamp 1704896540
transform 1 0 15456 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0848_
timestamp 1704896540
transform -1 0 18032 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0849_
timestamp 1704896540
transform 1 0 16928 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0850_
timestamp 1704896540
transform -1 0 16008 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0851_
timestamp 1704896540
transform -1 0 17296 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0852_
timestamp 1704896540
transform 1 0 17296 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0853_
timestamp 1704896540
transform 1 0 16652 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0854_
timestamp 1704896540
transform 1 0 17296 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0855_
timestamp 1704896540
transform -1 0 19320 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0856_
timestamp 1704896540
transform -1 0 19320 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0857_
timestamp 1704896540
transform -1 0 18860 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0858_
timestamp 1704896540
transform 1 0 16744 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0859_
timestamp 1704896540
transform -1 0 18216 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _0860_
timestamp 1704896540
transform 1 0 16836 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0861_
timestamp 1704896540
transform -1 0 18216 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0862_
timestamp 1704896540
transform 1 0 17756 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0863_
timestamp 1704896540
transform 1 0 17020 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0864_
timestamp 1704896540
transform -1 0 9292 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0865_
timestamp 1704896540
transform -1 0 1656 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0866_
timestamp 1704896540
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0867_
timestamp 1704896540
transform -1 0 2484 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0868_
timestamp 1704896540
transform 1 0 1748 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0869_
timestamp 1704896540
transform 1 0 1748 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0870_
timestamp 1704896540
transform 1 0 2668 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0871_
timestamp 1704896540
transform -1 0 4140 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0872_
timestamp 1704896540
transform 1 0 3220 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0873_
timestamp 1704896540
transform 1 0 3036 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0874_
timestamp 1704896540
transform 1 0 3496 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0875_
timestamp 1704896540
transform 1 0 5796 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0876_
timestamp 1704896540
transform -1 0 5428 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0877_
timestamp 1704896540
transform 1 0 4692 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0878_
timestamp 1704896540
transform -1 0 5244 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0879_
timestamp 1704896540
transform 1 0 5244 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0880_
timestamp 1704896540
transform 1 0 5796 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0881_
timestamp 1704896540
transform -1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0882_
timestamp 1704896540
transform -1 0 3128 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0883_
timestamp 1704896540
transform -1 0 6348 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0884_
timestamp 1704896540
transform 1 0 4784 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0885_
timestamp 1704896540
transform 1 0 3956 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0886_
timestamp 1704896540
transform 1 0 4876 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0887_
timestamp 1704896540
transform -1 0 3680 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0888_
timestamp 1704896540
transform -1 0 4048 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0889_
timestamp 1704896540
transform 1 0 2392 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0890_
timestamp 1704896540
transform -1 0 3404 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0891_
timestamp 1704896540
transform -1 0 3128 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0892_
timestamp 1704896540
transform 1 0 1380 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0893_
timestamp 1704896540
transform 1 0 1564 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0894_
timestamp 1704896540
transform -1 0 2116 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0895_
timestamp 1704896540
transform -1 0 1840 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0896_
timestamp 1704896540
transform -1 0 18308 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0897_
timestamp 1704896540
transform -1 0 18032 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0898_
timestamp 1704896540
transform 1 0 16284 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0899_
timestamp 1704896540
transform -1 0 16652 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0900_
timestamp 1704896540
transform 1 0 15272 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _0901_
timestamp 1704896540
transform 1 0 15824 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0902_
timestamp 1704896540
transform 1 0 14812 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0903_
timestamp 1704896540
transform 1 0 14352 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0904_
timestamp 1704896540
transform -1 0 14260 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0905_
timestamp 1704896540
transform -1 0 15180 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0906_
timestamp 1704896540
transform -1 0 15364 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0907_
timestamp 1704896540
transform 1 0 13800 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0908_
timestamp 1704896540
transform 1 0 14628 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0909_
timestamp 1704896540
transform 1 0 14628 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0910_
timestamp 1704896540
transform -1 0 15916 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0911_
timestamp 1704896540
transform 1 0 13708 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1704896540
transform 1 0 13892 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0913_
timestamp 1704896540
transform 1 0 14260 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0914_
timestamp 1704896540
transform -1 0 15456 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0915_
timestamp 1704896540
transform 1 0 14168 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0916_
timestamp 1704896540
transform 1 0 14352 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0917_
timestamp 1704896540
transform 1 0 14812 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0918_
timestamp 1704896540
transform -1 0 16192 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0919_
timestamp 1704896540
transform 1 0 13616 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0920_
timestamp 1704896540
transform 1 0 14904 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0921_
timestamp 1704896540
transform 1 0 14904 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0922_
timestamp 1704896540
transform -1 0 16376 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0923_
timestamp 1704896540
transform -1 0 12972 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0924_
timestamp 1704896540
transform -1 0 12788 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0925_
timestamp 1704896540
transform 1 0 11684 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0926_
timestamp 1704896540
transform 1 0 11960 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0927_
timestamp 1704896540
transform 1 0 13064 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0928_
timestamp 1704896540
transform 1 0 11500 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0929_
timestamp 1704896540
transform 1 0 12972 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0930_
timestamp 1704896540
transform 1 0 14352 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0931_
timestamp 1704896540
transform 1 0 13708 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0932_
timestamp 1704896540
transform -1 0 15272 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0933_
timestamp 1704896540
transform -1 0 14076 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1704896540
transform -1 0 13156 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0935_
timestamp 1704896540
transform -1 0 14352 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0936_
timestamp 1704896540
transform 1 0 13524 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0937_
timestamp 1704896540
transform 1 0 12788 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0938_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9384 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0939_
timestamp 1704896540
transform 1 0 10488 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0940_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6348 0 1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0941_
timestamp 1704896540
transform 1 0 2300 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0942_
timestamp 1704896540
transform 1 0 1656 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0943_
timestamp 1704896540
transform -1 0 20148 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0944_
timestamp 1704896540
transform 1 0 21252 0 1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0945_
timestamp 1704896540
transform 1 0 19320 0 -1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0946_
timestamp 1704896540
transform 1 0 23828 0 -1 24480
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0947_
timestamp 1704896540
transform 1 0 23828 0 1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0948_
timestamp 1704896540
transform 1 0 22908 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0949_
timestamp 1704896540
transform 1 0 18676 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0950_
timestamp 1704896540
transform 1 0 19596 0 -1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0951_
timestamp 1704896540
transform 1 0 18768 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0952_
timestamp 1704896540
transform 1 0 9384 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0953_
timestamp 1704896540
transform 1 0 11132 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0954_
timestamp 1704896540
transform 1 0 13156 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0955_
timestamp 1704896540
transform -1 0 24380 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0956_
timestamp 1704896540
transform 1 0 23000 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0957_
timestamp 1704896540
transform -1 0 23000 0 -1 27744
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0958_
timestamp 1704896540
transform 1 0 20608 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0959_
timestamp 1704896540
transform -1 0 21160 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0960_
timestamp 1704896540
transform 1 0 19044 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0961_
timestamp 1704896540
transform 1 0 19136 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0962_
timestamp 1704896540
transform 1 0 17664 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0963_
timestamp 1704896540
transform -1 0 21988 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0964_
timestamp 1704896540
transform -1 0 23092 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0965_
timestamp 1704896540
transform -1 0 22632 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0966_
timestamp 1704896540
transform -1 0 21252 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0967_
timestamp 1704896540
transform -1 0 18124 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0968_
timestamp 1704896540
transform 1 0 11684 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0969_
timestamp 1704896540
transform 1 0 11224 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0970_
timestamp 1704896540
transform -1 0 18032 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0971_
timestamp 1704896540
transform -1 0 5244 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0972_
timestamp 1704896540
transform 1 0 1472 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0973_
timestamp 1704896540
transform 1 0 1472 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0974_
timestamp 1704896540
transform 1 0 2944 0 -1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0975_
timestamp 1704896540
transform 1 0 5888 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0976_
timestamp 1704896540
transform -1 0 7728 0 1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0977_
timestamp 1704896540
transform 1 0 9844 0 1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0978_
timestamp 1704896540
transform 1 0 7820 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1704896540
transform 1 0 11040 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1704896540
transform 1 0 10948 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0981_
timestamp 1704896540
transform -1 0 10856 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1704896540
transform 1 0 12512 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0983_
timestamp 1704896540
transform -1 0 11316 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1704896540
transform 1 0 17664 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1704896540
transform 1 0 828 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1704896540
transform 1 0 1472 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1704896540
transform 1 0 2944 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0988_
timestamp 1704896540
transform 1 0 4140 0 1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1704896540
transform 1 0 5520 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1704896540
transform 1 0 3220 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1704896540
transform 1 0 4140 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0992_
timestamp 1704896540
transform 1 0 1564 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1704896540
transform 1 0 1288 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0994_
timestamp 1704896540
transform 1 0 1012 0 1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1704896540
transform 1 0 14352 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0996_
timestamp 1704896540
transform 1 0 15364 0 1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0997_
timestamp 1704896540
transform 1 0 16100 0 -1 27744
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0998_
timestamp 1704896540
transform 1 0 16100 0 -1 24480
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0999_
timestamp 1704896540
transform 1 0 16192 0 1 24480
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1000_
timestamp 1704896540
transform 1 0 16468 0 -1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1704896540
transform 1 0 11684 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1002_
timestamp 1704896540
transform 1 0 11132 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1704896540
transform -1 0 16836 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1004_
timestamp 1704896540
transform 1 0 14076 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1704896540
transform 1 0 12512 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  _1006_
timestamp 1704896540
transform 1 0 15272 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1007_
timestamp 1704896540
transform 1 0 12604 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1008_
timestamp 1704896540
transform 1 0 11132 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1009_
timestamp 1704896540
transform 1 0 8740 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1010_
timestamp 1704896540
transform -1 0 7360 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1011_
timestamp 1704896540
transform -1 0 5704 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1012_
timestamp 1704896540
transform -1 0 4324 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1013_
timestamp 1704896540
transform -1 0 1932 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15364 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1704896540
transform -1 0 7636 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1704896540
transform 1 0 7820 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1704896540
transform -1 0 7636 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1704896540
transform 1 0 7820 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1704896540
transform 1 0 13524 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1704896540
transform 1 0 18676 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1704896540
transform -1 0 17480 0 1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1704896540
transform 1 0 18676 0 1 23392
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1704896540
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1704896540
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1704896540
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1704896540
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1704896540
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1704896540
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1704896540
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1704896540
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1704896540
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1704896540
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1704896540
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1704896540
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1704896540
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1704896540
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1704896540
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1704896540
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1704896540
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1704896540
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1704896540
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_293 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 27508 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_299
timestamp 1704896540
transform 1 0 28060 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1704896540
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1704896540
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1704896540
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1704896540
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1704896540
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1704896540
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1704896540
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1704896540
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1704896540
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1704896540
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1704896540
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1704896540
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1704896540
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1704896540
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1704896540
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1704896540
transform 1 0 22356 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1704896540
transform 1 0 23460 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1704896540
transform 1 0 24564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1704896540
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1704896540
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1704896540
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_293
timestamp 1704896540
transform 1 0 27508 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_299
timestamp 1704896540
transform 1 0 28060 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1704896540
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1704896540
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1704896540
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1704896540
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1704896540
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1704896540
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1704896540
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1704896540
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1704896540
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1704896540
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1704896540
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1704896540
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1704896540
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1704896540
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1704896540
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1704896540
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1704896540
transform 1 0 23092 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1704896540
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1704896540
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1704896540
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1704896540
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_289 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 27140 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_297
timestamp 1704896540
transform 1 0 27876 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1704896540
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1704896540
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1704896540
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1704896540
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1704896540
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1704896540
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1704896540
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1704896540
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1704896540
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1704896540
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1704896540
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1704896540
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1704896540
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1704896540
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1704896540
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1704896540
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1704896540
transform 1 0 23460 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1704896540
transform 1 0 24564 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1704896540
transform 1 0 25668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1704896540
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1704896540
transform 1 0 26404 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_293
timestamp 1704896540
transform 1 0 27508 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_299
timestamp 1704896540
transform 1 0 28060 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1704896540
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1704896540
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1704896540
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1704896540
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1704896540
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1704896540
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1704896540
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1704896540
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1704896540
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1704896540
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1704896540
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1704896540
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1704896540
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1704896540
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1704896540
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1704896540
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1704896540
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1704896540
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1704896540
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1704896540
transform 1 0 23092 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1704896540
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1704896540
transform 1 0 23828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1704896540
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1704896540
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_289
timestamp 1704896540
transform 1 0 27140 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_297
timestamp 1704896540
transform 1 0 27876 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1704896540
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1704896540
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1704896540
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1704896540
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1704896540
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1704896540
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1704896540
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1704896540
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1704896540
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1704896540
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1704896540
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1704896540
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1704896540
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1704896540
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1704896540
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1704896540
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1704896540
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1704896540
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1704896540
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1704896540
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1704896540
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1704896540
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1704896540
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1704896540
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1704896540
transform 1 0 26404 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_293
timestamp 1704896540
transform 1 0 27508 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_299
timestamp 1704896540
transform 1 0 28060 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1704896540
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1704896540
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1704896540
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1704896540
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1704896540
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1704896540
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1704896540
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1704896540
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1704896540
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1704896540
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1704896540
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1704896540
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1704896540
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1704896540
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1704896540
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1704896540
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1704896540
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1704896540
transform 1 0 21988 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1704896540
transform 1 0 23092 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1704896540
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1704896540
transform 1 0 23828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1704896540
transform 1 0 24932 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1704896540
transform 1 0 26036 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_289
timestamp 1704896540
transform 1 0 27140 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_297
timestamp 1704896540
transform 1 0 27876 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1704896540
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1704896540
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1704896540
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1704896540
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1704896540
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1704896540
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1704896540
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1704896540
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1704896540
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1704896540
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1704896540
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1704896540
transform 1 0 20516 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1704896540
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1704896540
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1704896540
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1704896540
transform 1 0 23460 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1704896540
transform 1 0 24564 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1704896540
transform 1 0 25668 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1704896540
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1704896540
transform 1 0 26404 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_293
timestamp 1704896540
transform 1 0 27508 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_299
timestamp 1704896540
transform 1 0 28060 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1704896540
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1704896540
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1704896540
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1704896540
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1704896540
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1704896540
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1704896540
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1704896540
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1704896540
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1704896540
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1704896540
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1704896540
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1704896540
transform 1 0 17940 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1704896540
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1704896540
transform 1 0 18676 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1704896540
transform 1 0 19780 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1704896540
transform 1 0 20884 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1704896540
transform 1 0 21988 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1704896540
transform 1 0 23092 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1704896540
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1704896540
transform 1 0 23828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1704896540
transform 1 0 24932 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1704896540
transform 1 0 26036 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_289
timestamp 1704896540
transform 1 0 27140 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_297
timestamp 1704896540
transform 1 0 27876 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1704896540
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1704896540
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1704896540
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1704896540
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1704896540
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1704896540
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1704896540
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1704896540
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1704896540
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1704896540
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1704896540
transform 1 0 12052 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1704896540
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1704896540
transform 1 0 14260 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1704896540
transform 1 0 15364 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1704896540
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1704896540
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1704896540
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1704896540
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1704896540
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1704896540
transform 1 0 20516 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1704896540
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1704896540
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1704896540
transform 1 0 22356 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1704896540
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1704896540
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1704896540
transform 1 0 25668 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1704896540
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1704896540
transform 1 0 26404 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_293
timestamp 1704896540
transform 1 0 27508 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_299
timestamp 1704896540
transform 1 0 28060 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1704896540
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1704896540
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1704896540
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1704896540
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1704896540
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1704896540
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1704896540
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1704896540
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1704896540
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1704896540
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1704896540
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1704896540
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1704896540
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1704896540
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1704896540
transform 1 0 17940 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1704896540
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1704896540
transform 1 0 18676 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1704896540
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1704896540
transform 1 0 20884 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1704896540
transform 1 0 21988 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1704896540
transform 1 0 23092 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1704896540
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1704896540
transform 1 0 23828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1704896540
transform 1 0 24932 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1704896540
transform 1 0 26036 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_289
timestamp 1704896540
transform 1 0 27140 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_297
timestamp 1704896540
transform 1 0 27876 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1704896540
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1704896540
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1704896540
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1704896540
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1704896540
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1704896540
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1704896540
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1704896540
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1704896540
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1704896540
transform 1 0 10212 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1704896540
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1704896540
transform 1 0 10948 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1704896540
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1704896540
transform 1 0 13156 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1704896540
transform 1 0 14260 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1704896540
transform 1 0 15364 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1704896540
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1704896540
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1704896540
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1704896540
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1704896540
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1704896540
transform 1 0 20516 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1704896540
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1704896540
transform 1 0 21252 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1704896540
transform 1 0 22356 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1704896540
transform 1 0 23460 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1704896540
transform 1 0 24564 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1704896540
transform 1 0 25668 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1704896540
transform 1 0 26220 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1704896540
transform 1 0 26404 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_293
timestamp 1704896540
transform 1 0 27508 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_299
timestamp 1704896540
transform 1 0 28060 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1704896540
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1704896540
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1704896540
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1704896540
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1704896540
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1704896540
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1704896540
transform 1 0 9476 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1704896540
transform 1 0 10580 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1704896540
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1704896540
transform 1 0 12788 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1704896540
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1704896540
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1704896540
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1704896540
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1704896540
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1704896540
transform 1 0 17940 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1704896540
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1704896540
transform 1 0 18676 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1704896540
transform 1 0 19780 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1704896540
transform 1 0 20884 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1704896540
transform 1 0 21988 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1704896540
transform 1 0 23092 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1704896540
transform 1 0 23644 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1704896540
transform 1 0 23828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1704896540
transform 1 0 24932 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1704896540
transform 1 0 26036 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_289
timestamp 1704896540
transform 1 0 27140 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_297
timestamp 1704896540
transform 1 0 27876 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1704896540
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1704896540
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1704896540
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1704896540
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1704896540
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1704896540
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1704896540
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1704896540
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1704896540
transform 1 0 10212 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1704896540
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1704896540
transform 1 0 10948 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1704896540
transform 1 0 12052 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1704896540
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1704896540
transform 1 0 14260 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1704896540
transform 1 0 15364 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1704896540
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1704896540
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1704896540
transform 1 0 17204 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1704896540
transform 1 0 18308 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1704896540
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1704896540
transform 1 0 20516 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1704896540
transform 1 0 21068 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1704896540
transform 1 0 21252 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1704896540
transform 1 0 22356 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1704896540
transform 1 0 23460 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1704896540
transform 1 0 24564 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1704896540
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1704896540
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1704896540
transform 1 0 26404 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_293
timestamp 1704896540
transform 1 0 27508 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_299
timestamp 1704896540
transform 1 0 28060 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1704896540
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1704896540
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1704896540
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1704896540
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1704896540
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1704896540
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1704896540
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8372 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1704896540
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1704896540
transform 1 0 10580 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1704896540
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1704896540
transform 1 0 12788 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1704896540
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1704896540
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1704896540
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1704896540
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1704896540
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1704896540
transform 1 0 17940 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1704896540
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1704896540
transform 1 0 18676 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1704896540
transform 1 0 19780 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1704896540
transform 1 0 20884 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1704896540
transform 1 0 21988 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1704896540
transform 1 0 23092 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1704896540
transform 1 0 23644 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1704896540
transform 1 0 23828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1704896540
transform 1 0 24932 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1704896540
transform 1 0 26036 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_289
timestamp 1704896540
transform 1 0 27140 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_297
timestamp 1704896540
transform 1 0 27876 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1704896540
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1704896540
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1704896540
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1704896540
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1704896540
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1704896540
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1704896540
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1704896540
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1704896540
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1704896540
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1704896540
transform 1 0 10212 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1704896540
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1704896540
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1704896540
transform 1 0 12052 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1704896540
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1704896540
transform 1 0 14260 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1704896540
transform 1 0 15364 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1704896540
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1704896540
transform 1 0 16100 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1704896540
transform 1 0 17204 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1704896540
transform 1 0 18308 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1704896540
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1704896540
transform 1 0 20516 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1704896540
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1704896540
transform 1 0 21252 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1704896540
transform 1 0 22356 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1704896540
transform 1 0 23460 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1704896540
transform 1 0 24564 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1704896540
transform 1 0 25668 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1704896540
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1704896540
transform 1 0 26404 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_293
timestamp 1704896540
transform 1 0 27508 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_299
timestamp 1704896540
transform 1 0 28060 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1704896540
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1704896540
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1704896540
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1704896540
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1704896540
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1704896540
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1704896540
transform 1 0 7636 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1704896540
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1704896540
transform 1 0 9476 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1704896540
transform 1 0 10580 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1704896540
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1704896540
transform 1 0 12788 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1704896540
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1704896540
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1704896540
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1704896540
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1704896540
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1704896540
transform 1 0 17940 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1704896540
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1704896540
transform 1 0 18676 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1704896540
transform 1 0 19780 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1704896540
transform 1 0 20884 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1704896540
transform 1 0 21988 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1704896540
transform 1 0 23092 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1704896540
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1704896540
transform 1 0 23828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1704896540
transform 1 0 24932 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1704896540
transform 1 0 26036 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_289
timestamp 1704896540
transform 1 0 27140 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_297
timestamp 1704896540
transform 1 0 27876 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1704896540
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1704896540
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1704896540
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1704896540
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1704896540
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1704896540
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1704896540
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_69
timestamp 1704896540
transform 1 0 6900 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_96
timestamp 1704896540
transform 1 0 9384 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_108
timestamp 1704896540
transform 1 0 10488 0 -1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1704896540
transform 1 0 10948 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1704896540
transform 1 0 12052 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1704896540
transform 1 0 13156 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1704896540
transform 1 0 14260 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1704896540
transform 1 0 15364 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1704896540
transform 1 0 15916 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1704896540
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1704896540
transform 1 0 17204 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1704896540
transform 1 0 18308 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1704896540
transform 1 0 19412 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1704896540
transform 1 0 20516 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1704896540
transform 1 0 21068 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1704896540
transform 1 0 21252 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1704896540
transform 1 0 22356 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1704896540
transform 1 0 23460 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1704896540
transform 1 0 24564 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1704896540
transform 1 0 25668 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1704896540
transform 1 0 26220 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1704896540
transform 1 0 26404 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_293
timestamp 1704896540
transform 1 0 27508 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_299
timestamp 1704896540
transform 1 0 28060 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1704896540
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1704896540
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1704896540
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_53
timestamp 1704896540
transform 1 0 5428 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_78
timestamp 1704896540
transform 1 0 7728 0 1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_97
timestamp 1704896540
transform 1 0 9476 0 1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1704896540
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1704896540
transform 1 0 12788 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1704896540
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1704896540
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1704896540
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_165
timestamp 1704896540
transform 1 0 15732 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_173
timestamp 1704896540
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_186
timestamp 1704896540
transform 1 0 17664 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1704896540
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1704896540
transform 1 0 18676 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1704896540
transform 1 0 19780 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1704896540
transform 1 0 20884 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 1704896540
transform 1 0 21988 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 1704896540
transform 1 0 23092 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1704896540
transform 1 0 23644 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1704896540
transform 1 0 23828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1704896540
transform 1 0 24932 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1704896540
transform 1 0 26036 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_289
timestamp 1704896540
transform 1 0 27140 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_297
timestamp 1704896540
transform 1 0 27876 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1704896540
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1704896540
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1704896540
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1704896540
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1704896540
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1704896540
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_57
timestamp 1704896540
transform 1 0 5796 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_65
timestamp 1704896540
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_75
timestamp 1704896540
transform 1 0 7452 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_81
timestamp 1704896540
transform 1 0 8004 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_85
timestamp 1704896540
transform 1 0 8372 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_94
timestamp 1704896540
transform 1 0 9200 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_102
timestamp 1704896540
transform 1 0 9936 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1704896540
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_137
timestamp 1704896540
transform 1 0 13156 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_147
timestamp 1704896540
transform 1 0 14076 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_151
timestamp 1704896540
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_160
timestamp 1704896540
transform 1 0 15272 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_190
timestamp 1704896540
transform 1 0 18032 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_202
timestamp 1704896540
transform 1 0 19136 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_214
timestamp 1704896540
transform 1 0 20240 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_222
timestamp 1704896540
transform 1 0 20976 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1704896540
transform 1 0 21252 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1704896540
transform 1 0 22356 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1704896540
transform 1 0 23460 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1704896540
transform 1 0 24564 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 1704896540
transform 1 0 25668 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1704896540
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1704896540
transform 1 0 26404 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_293
timestamp 1704896540
transform 1 0 27508 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_299
timestamp 1704896540
transform 1 0 28060 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1704896540
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1704896540
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3220 0 1 11424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_51
timestamp 1704896540
transform 1 0 5244 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_63
timestamp 1704896540
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_74
timestamp 1704896540
transform 1 0 7360 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1704896540
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8372 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_89
timestamp 1704896540
transform 1 0 8740 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_101
timestamp 1704896540
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_110
timestamp 1704896540
transform 1 0 10672 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_127
timestamp 1704896540
transform 1 0 12236 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_135
timestamp 1704896540
transform 1 0 12972 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_154
timestamp 1704896540
transform 1 0 14720 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_171
timestamp 1704896540
transform 1 0 16284 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_183
timestamp 1704896540
transform 1 0 17388 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_187
timestamp 1704896540
transform 1 0 17756 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1704896540
transform 1 0 18492 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_197
timestamp 1704896540
transform 1 0 18676 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_205
timestamp 1704896540
transform 1 0 19412 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_225
timestamp 1704896540
transform 1 0 21252 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_237
timestamp 1704896540
transform 1 0 22356 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_249
timestamp 1704896540
transform 1 0 23460 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1704896540
transform 1 0 23828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1704896540
transform 1 0 24932 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1704896540
transform 1 0 26036 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_289
timestamp 1704896540
transform 1 0 27140 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_297
timestamp 1704896540
transform 1 0 27876 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1704896540
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1704896540
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1704896540
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_39
timestamp 1704896540
transform 1 0 4140 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_43
timestamp 1704896540
transform 1 0 4508 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_47
timestamp 1704896540
transform 1 0 4876 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_65
timestamp 1704896540
transform 1 0 6532 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_82
timestamp 1704896540
transform 1 0 8096 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_88
timestamp 1704896540
transform 1 0 8648 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_95
timestamp 1704896540
transform 1 0 9292 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 1704896540
transform 1 0 10396 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1704896540
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_113
timestamp 1704896540
transform 1 0 10948 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_117
timestamp 1704896540
transform 1 0 11316 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_121
timestamp 1704896540
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_129
timestamp 1704896540
transform 1 0 12420 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_141
timestamp 1704896540
transform 1 0 13524 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_153
timestamp 1704896540
transform 1 0 14628 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_165
timestamp 1704896540
transform 1 0 15732 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1704896540
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1704896540
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_193
timestamp 1704896540
transform 1 0 18308 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_206
timestamp 1704896540
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 1704896540
transform 1 0 20976 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1704896540
transform 1 0 21252 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1704896540
transform 1 0 22356 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1704896540
transform 1 0 23460 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1704896540
transform 1 0 24564 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1704896540
transform 1 0 25668 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1704896540
transform 1 0 26220 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1704896540
transform 1 0 26404 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_293
timestamp 1704896540
transform 1 0 27508 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_299
timestamp 1704896540
transform 1 0 28060 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1704896540
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_15
timestamp 1704896540
transform 1 0 1932 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_21
timestamp 1704896540
transform 1 0 2484 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1704896540
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3220 0 1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_40
timestamp 1704896540
transform 1 0 4232 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_52
timestamp 1704896540
transform 1 0 5336 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_56
timestamp 1704896540
transform 1 0 5704 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_64
timestamp 1704896540
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1704896540
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8372 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_93
timestamp 1704896540
transform 1 0 9108 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_99
timestamp 1704896540
transform 1 0 9660 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_114
timestamp 1704896540
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_138
timestamp 1704896540
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_146
timestamp 1704896540
transform 1 0 13984 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_161
timestamp 1704896540
transform 1 0 15364 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_165
timestamp 1704896540
transform 1 0 15732 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_173
timestamp 1704896540
transform 1 0 16468 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_191
timestamp 1704896540
transform 1 0 18124 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1704896540
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1704896540
transform 1 0 18676 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1704896540
transform 1 0 19780 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1704896540
transform 1 0 20884 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1704896540
transform 1 0 21988 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 1704896540
transform 1 0 23092 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1704896540
transform 1 0 23644 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1704896540
transform 1 0 23828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1704896540
transform 1 0 24932 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1704896540
transform 1 0 26036 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_289
timestamp 1704896540
transform 1 0 27140 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_297
timestamp 1704896540
transform 1 0 27876 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_3
timestamp 1704896540
transform 1 0 828 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_9
timestamp 1704896540
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_33
timestamp 1704896540
transform 1 0 3588 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_48
timestamp 1704896540
transform 1 0 4968 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_77
timestamp 1704896540
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 1704896540
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_113
timestamp 1704896540
transform 1 0 10948 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_123
timestamp 1704896540
transform 1 0 11868 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_131
timestamp 1704896540
transform 1 0 12604 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_146
timestamp 1704896540
transform 1 0 13984 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_155
timestamp 1704896540
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1704896540
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_172
timestamp 1704896540
transform 1 0 16376 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_191
timestamp 1704896540
transform 1 0 18124 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_211
timestamp 1704896540
transform 1 0 19964 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1704896540
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_230
timestamp 1704896540
transform 1 0 21712 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_242
timestamp 1704896540
transform 1 0 22816 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_254
timestamp 1704896540
transform 1 0 23920 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_266
timestamp 1704896540
transform 1 0 25024 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_278
timestamp 1704896540
transform 1 0 26128 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1704896540
transform 1 0 26404 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_293
timestamp 1704896540
transform 1 0 27508 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_299
timestamp 1704896540
transform 1 0 28060 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_3
timestamp 1704896540
transform 1 0 828 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_11
timestamp 1704896540
transform 1 0 1564 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_17
timestamp 1704896540
transform 1 0 2116 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_25
timestamp 1704896540
transform 1 0 2852 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_29
timestamp 1704896540
transform 1 0 3220 0 1 13600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_40
timestamp 1704896540
transform 1 0 4232 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_52
timestamp 1704896540
transform 1 0 5336 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_60
timestamp 1704896540
transform 1 0 6072 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_80
timestamp 1704896540
transform 1 0 7912 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_85
timestamp 1704896540
transform 1 0 8372 0 1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_95
timestamp 1704896540
transform 1 0 9292 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_107
timestamp 1704896540
transform 1 0 10396 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_115
timestamp 1704896540
transform 1 0 11132 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1704896540
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1704896540
transform 1 0 12788 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1704896540
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1704896540
transform 1 0 13524 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_145
timestamp 1704896540
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_157
timestamp 1704896540
transform 1 0 14996 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_169
timestamp 1704896540
transform 1 0 16100 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_181
timestamp 1704896540
transform 1 0 17204 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_193
timestamp 1704896540
transform 1 0 18308 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_203
timestamp 1704896540
transform 1 0 19228 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_207
timestamp 1704896540
transform 1 0 19596 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_215
timestamp 1704896540
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_240
timestamp 1704896540
transform 1 0 22632 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1704896540
transform 1 0 23828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1704896540
transform 1 0 24932 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1704896540
transform 1 0 26036 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_289
timestamp 1704896540
transform 1 0 27140 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_297
timestamp 1704896540
transform 1 0 27876 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1704896540
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1704896540
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_27
timestamp 1704896540
transform 1 0 3036 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_32
timestamp 1704896540
transform 1 0 3496 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_40
timestamp 1704896540
transform 1 0 4232 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_52
timestamp 1704896540
transform 1 0 5336 0 -1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_65
timestamp 1704896540
transform 1 0 6532 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_77
timestamp 1704896540
transform 1 0 7636 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_85
timestamp 1704896540
transform 1 0 8372 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_92
timestamp 1704896540
transform 1 0 9016 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_104
timestamp 1704896540
transform 1 0 10120 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_113
timestamp 1704896540
transform 1 0 10948 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_150
timestamp 1704896540
transform 1 0 14352 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_159
timestamp 1704896540
transform 1 0 15180 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_174
timestamp 1704896540
transform 1 0 16560 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_183
timestamp 1704896540
transform 1 0 17388 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_195
timestamp 1704896540
transform 1 0 18492 0 -1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1704896540
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1704896540
transform 1 0 20516 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1704896540
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_225
timestamp 1704896540
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_230
timestamp 1704896540
transform 1 0 21712 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_242
timestamp 1704896540
transform 1 0 22816 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_254
timestamp 1704896540
transform 1 0 23920 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_266
timestamp 1704896540
transform 1 0 25024 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_278
timestamp 1704896540
transform 1 0 26128 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1704896540
transform 1 0 26404 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_293
timestamp 1704896540
transform 1 0 27508 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_299
timestamp 1704896540
transform 1 0 28060 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1704896540
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_15
timestamp 1704896540
transform 1 0 1932 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_47
timestamp 1704896540
transform 1 0 4876 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_55
timestamp 1704896540
transform 1 0 5612 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_74
timestamp 1704896540
transform 1 0 7360 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_85
timestamp 1704896540
transform 1 0 8372 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_95
timestamp 1704896540
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_104
timestamp 1704896540
transform 1 0 10120 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_124
timestamp 1704896540
transform 1 0 11960 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_132
timestamp 1704896540
transform 1 0 12696 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_141
timestamp 1704896540
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_157
timestamp 1704896540
transform 1 0 14996 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_161
timestamp 1704896540
transform 1 0 15364 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_169
timestamp 1704896540
transform 1 0 16100 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_181
timestamp 1704896540
transform 1 0 17204 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_189
timestamp 1704896540
transform 1 0 17940 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1704896540
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_213
timestamp 1704896540
transform 1 0 20148 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_221
timestamp 1704896540
transform 1 0 20884 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_234
timestamp 1704896540
transform 1 0 22080 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_246
timestamp 1704896540
transform 1 0 23184 0 1 14688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1704896540
transform 1 0 23828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1704896540
transform 1 0 24932 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1704896540
transform 1 0 26036 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_289
timestamp 1704896540
transform 1 0 27140 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_297
timestamp 1704896540
transform 1 0 27876 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1704896540
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_15
timestamp 1704896540
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_22
timestamp 1704896540
transform 1 0 2576 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_34
timestamp 1704896540
transform 1 0 3680 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_42
timestamp 1704896540
transform 1 0 4416 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_52
timestamp 1704896540
transform 1 0 5336 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_57
timestamp 1704896540
transform 1 0 5796 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_63
timestamp 1704896540
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_68
timestamp 1704896540
transform 1 0 6808 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_80
timestamp 1704896540
transform 1 0 7912 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_86
timestamp 1704896540
transform 1 0 8464 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_95
timestamp 1704896540
transform 1 0 9292 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_107
timestamp 1704896540
transform 1 0 10396 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1704896540
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1704896540
transform 1 0 10948 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1704896540
transform 1 0 12052 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_137
timestamp 1704896540
transform 1 0 13156 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_142
timestamp 1704896540
transform 1 0 13616 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_154
timestamp 1704896540
transform 1 0 14720 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1704896540
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_169
timestamp 1704896540
transform 1 0 16100 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_177
timestamp 1704896540
transform 1 0 16836 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_190
timestamp 1704896540
transform 1 0 18032 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_196
timestamp 1704896540
transform 1 0 18584 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_204
timestamp 1704896540
transform 1 0 19320 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_245
timestamp 1704896540
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_257
timestamp 1704896540
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_269
timestamp 1704896540
transform 1 0 25300 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_277
timestamp 1704896540
transform 1 0 26036 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1704896540
transform 1 0 26404 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_293
timestamp 1704896540
transform 1 0 27508 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_299
timestamp 1704896540
transform 1 0 28060 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_3
timestamp 1704896540
transform 1 0 828 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_9
timestamp 1704896540
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_26
timestamp 1704896540
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_36
timestamp 1704896540
transform 1 0 3864 0 1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_47
timestamp 1704896540
transform 1 0 4876 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_59
timestamp 1704896540
transform 1 0 5980 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_65
timestamp 1704896540
transform 1 0 6532 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_70
timestamp 1704896540
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_75
timestamp 1704896540
transform 1 0 7452 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1704896540
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_85
timestamp 1704896540
transform 1 0 8372 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_89
timestamp 1704896540
transform 1 0 8740 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_97
timestamp 1704896540
transform 1 0 9476 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_123
timestamp 1704896540
transform 1 0 11868 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_131
timestamp 1704896540
transform 1 0 12604 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_138
timestamp 1704896540
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_151
timestamp 1704896540
transform 1 0 14444 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_157
timestamp 1704896540
transform 1 0 14996 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_166
timestamp 1704896540
transform 1 0 15824 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_174
timestamp 1704896540
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_192
timestamp 1704896540
transform 1 0 18216 0 1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1704896540
transform 1 0 21988 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1704896540
transform 1 0 23092 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1704896540
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1704896540
transform 1 0 23828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1704896540
transform 1 0 24932 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1704896540
transform 1 0 26036 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_289
timestamp 1704896540
transform 1 0 27140 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_297
timestamp 1704896540
transform 1 0 27876 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1704896540
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_18
timestamp 1704896540
transform 1 0 2208 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_30
timestamp 1704896540
transform 1 0 3312 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_38
timestamp 1704896540
transform 1 0 4048 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_46
timestamp 1704896540
transform 1 0 4784 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_57
timestamp 1704896540
transform 1 0 5796 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_94
timestamp 1704896540
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_101
timestamp 1704896540
transform 1 0 9844 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_107
timestamp 1704896540
transform 1 0 10396 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1704896540
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_113
timestamp 1704896540
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_132
timestamp 1704896540
transform 1 0 12696 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1704896540
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_149
timestamp 1704896540
transform 1 0 14260 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_162
timestamp 1704896540
transform 1 0 15456 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_169
timestamp 1704896540
transform 1 0 16100 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_192
timestamp 1704896540
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_199
timestamp 1704896540
transform 1 0 18860 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_214
timestamp 1704896540
transform 1 0 20240 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_222
timestamp 1704896540
transform 1 0 20976 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1704896540
transform 1 0 21252 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1704896540
transform 1 0 22356 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1704896540
transform 1 0 23460 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1704896540
transform 1 0 24564 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1704896540
transform 1 0 25668 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1704896540
transform 1 0 26220 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1704896540
transform 1 0 26404 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_293
timestamp 1704896540
transform 1 0 27508 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_299
timestamp 1704896540
transform 1 0 28060 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1704896540
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1704896540
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1704896540
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_37
timestamp 1704896540
transform 1 0 3956 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_49
timestamp 1704896540
transform 1 0 5060 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_61
timestamp 1704896540
transform 1 0 6164 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_73
timestamp 1704896540
transform 1 0 7268 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1704896540
transform 1 0 8004 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_92
timestamp 1704896540
transform 1 0 9016 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_98
timestamp 1704896540
transform 1 0 9568 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_104
timestamp 1704896540
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_116
timestamp 1704896540
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_128
timestamp 1704896540
transform 1 0 12328 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_141
timestamp 1704896540
transform 1 0 13524 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_151
timestamp 1704896540
transform 1 0 14444 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_175
timestamp 1704896540
transform 1 0 16652 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1704896540
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_204
timestamp 1704896540
transform 1 0 19320 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_212
timestamp 1704896540
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_220
timestamp 1704896540
transform 1 0 20792 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_232
timestamp 1704896540
transform 1 0 21896 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_244
timestamp 1704896540
transform 1 0 23000 0 1 16864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1704896540
transform 1 0 23828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1704896540
transform 1 0 24932 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1704896540
transform 1 0 26036 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_289
timestamp 1704896540
transform 1 0 27140 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_297
timestamp 1704896540
transform 1 0 27876 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1704896540
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_15
timestamp 1704896540
transform 1 0 1932 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_23
timestamp 1704896540
transform 1 0 2668 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_43
timestamp 1704896540
transform 1 0 4508 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1704896540
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_66
timestamp 1704896540
transform 1 0 6624 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_70
timestamp 1704896540
transform 1 0 6992 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_74
timestamp 1704896540
transform 1 0 7360 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_82
timestamp 1704896540
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_92
timestamp 1704896540
transform 1 0 9016 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_116
timestamp 1704896540
transform 1 0 11224 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_127
timestamp 1704896540
transform 1 0 12236 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_160
timestamp 1704896540
transform 1 0 15272 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_177
timestamp 1704896540
transform 1 0 16836 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_185
timestamp 1704896540
transform 1 0 17572 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_202
timestamp 1704896540
transform 1 0 19136 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_206
timestamp 1704896540
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1704896540
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1704896540
transform 1 0 22356 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1704896540
transform 1 0 23460 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1704896540
transform 1 0 24564 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1704896540
transform 1 0 25668 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1704896540
transform 1 0 26220 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1704896540
transform 1 0 26404 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_293
timestamp 1704896540
transform 1 0 27508 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_299
timestamp 1704896540
transform 1 0 28060 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_3
timestamp 1704896540
transform 1 0 828 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_29
timestamp 1704896540
transform 1 0 3220 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_37
timestamp 1704896540
transform 1 0 3956 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_53
timestamp 1704896540
transform 1 0 5428 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_57
timestamp 1704896540
transform 1 0 5796 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_65
timestamp 1704896540
transform 1 0 6532 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_74
timestamp 1704896540
transform 1 0 7360 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_85
timestamp 1704896540
transform 1 0 8372 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_102
timestamp 1704896540
transform 1 0 9936 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_114
timestamp 1704896540
transform 1 0 11040 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_120
timestamp 1704896540
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_133
timestamp 1704896540
transform 1 0 12788 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_185
timestamp 1704896540
transform 1 0 17572 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_193
timestamp 1704896540
transform 1 0 18308 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_197
timestamp 1704896540
transform 1 0 18676 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_205
timestamp 1704896540
transform 1 0 19412 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1704896540
transform 1 0 19780 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1704896540
transform 1 0 20884 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1704896540
transform 1 0 21988 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1704896540
transform 1 0 23092 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1704896540
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1704896540
transform 1 0 23828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1704896540
transform 1 0 24932 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1704896540
transform 1 0 26036 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_289
timestamp 1704896540
transform 1 0 27140 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_297
timestamp 1704896540
transform 1 0 27876 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1704896540
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1704896540
transform 1 0 1932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_27
timestamp 1704896540
transform 1 0 3036 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_31
timestamp 1704896540
transform 1 0 3404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_40
timestamp 1704896540
transform 1 0 4232 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_50
timestamp 1704896540
transform 1 0 5152 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_57
timestamp 1704896540
transform 1 0 5796 0 -1 19040
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_72
timestamp 1704896540
transform 1 0 7176 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_84
timestamp 1704896540
transform 1 0 8280 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_88
timestamp 1704896540
transform 1 0 8648 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1704896540
transform 1 0 9108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1704896540
transform 1 0 10212 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1704896540
transform 1 0 10764 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_127
timestamp 1704896540
transform 1 0 12236 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_135
timestamp 1704896540
transform 1 0 12972 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_150
timestamp 1704896540
transform 1 0 14352 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_162
timestamp 1704896540
transform 1 0 15456 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_169
timestamp 1704896540
transform 1 0 16100 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_186
timestamp 1704896540
transform 1 0 17664 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_194
timestamp 1704896540
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_200
timestamp 1704896540
transform 1 0 18952 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_208
timestamp 1704896540
transform 1 0 19688 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1704896540
transform 1 0 21068 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_225
timestamp 1704896540
transform 1 0 21252 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_237
timestamp 1704896540
transform 1 0 22356 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_245
timestamp 1704896540
transform 1 0 23092 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_254
timestamp 1704896540
transform 1 0 23920 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_266
timestamp 1704896540
transform 1 0 25024 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_278
timestamp 1704896540
transform 1 0 26128 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1704896540
transform 1 0 26404 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_293
timestamp 1704896540
transform 1 0 27508 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_299
timestamp 1704896540
transform 1 0 28060 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_3
timestamp 1704896540
transform 1 0 828 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_16
timestamp 1704896540
transform 1 0 2024 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_38
timestamp 1704896540
transform 1 0 4048 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_55
timestamp 1704896540
transform 1 0 5612 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_63
timestamp 1704896540
transform 1 0 6348 0 1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_70
timestamp 1704896540
transform 1 0 6992 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_82
timestamp 1704896540
transform 1 0 8096 0 1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_108
timestamp 1704896540
transform 1 0 10488 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_120
timestamp 1704896540
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_137
timestamp 1704896540
transform 1 0 13156 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_161
timestamp 1704896540
transform 1 0 15364 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_169
timestamp 1704896540
transform 1 0 16100 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_181
timestamp 1704896540
transform 1 0 17204 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_223
timestamp 1704896540
transform 1 0 21068 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_237
timestamp 1704896540
transform 1 0 22356 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_244
timestamp 1704896540
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_249
timestamp 1704896540
transform 1 0 23460 0 1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1704896540
transform 1 0 23828 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 1704896540
transform 1 0 24932 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 1704896540
transform 1 0 26036 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_289
timestamp 1704896540
transform 1 0 27140 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_297
timestamp 1704896540
transform 1 0 27876 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_3
timestamp 1704896540
transform 1 0 828 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_7
timestamp 1704896540
transform 1 0 1196 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_24
timestamp 1704896540
transform 1 0 2760 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_31
timestamp 1704896540
transform 1 0 3404 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_44
timestamp 1704896540
transform 1 0 4600 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_53
timestamp 1704896540
transform 1 0 5428 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_57
timestamp 1704896540
transform 1 0 5796 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_77
timestamp 1704896540
transform 1 0 7636 0 -1 20128
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_86
timestamp 1704896540
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_98
timestamp 1704896540
transform 1 0 9568 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_107
timestamp 1704896540
transform 1 0 10396 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1704896540
transform 1 0 10764 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_129
timestamp 1704896540
transform 1 0 12420 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_133
timestamp 1704896540
transform 1 0 12788 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_164
timestamp 1704896540
transform 1 0 15640 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_169
timestamp 1704896540
transform 1 0 16100 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_182
timestamp 1704896540
transform 1 0 17296 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_194
timestamp 1704896540
transform 1 0 18400 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_200
timestamp 1704896540
transform 1 0 18952 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_214
timestamp 1704896540
transform 1 0 20240 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_218
timestamp 1704896540
transform 1 0 20608 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_229
timestamp 1704896540
transform 1 0 21620 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_235
timestamp 1704896540
transform 1 0 22172 0 -1 20128
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_260
timestamp 1704896540
transform 1 0 24472 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_272
timestamp 1704896540
transform 1 0 25576 0 -1 20128
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1704896540
transform 1 0 26404 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_293
timestamp 1704896540
transform 1 0 27508 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_299
timestamp 1704896540
transform 1 0 28060 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_3
timestamp 1704896540
transform 1 0 828 0 1 20128
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_14
timestamp 1704896540
transform 1 0 1840 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_26
timestamp 1704896540
transform 1 0 2944 0 1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1704896540
transform 1 0 3220 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1704896540
transform 1 0 4324 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_53
timestamp 1704896540
transform 1 0 5428 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_60
timestamp 1704896540
transform 1 0 6072 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_66
timestamp 1704896540
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_75
timestamp 1704896540
transform 1 0 7452 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1704896540
transform 1 0 8188 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_99
timestamp 1704896540
transform 1 0 9660 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_111
timestamp 1704896540
transform 1 0 10764 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_118
timestamp 1704896540
transform 1 0 11408 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_129
timestamp 1704896540
transform 1 0 12420 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_137
timestamp 1704896540
transform 1 0 13156 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_145
timestamp 1704896540
transform 1 0 13892 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_153
timestamp 1704896540
transform 1 0 14628 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_163
timestamp 1704896540
transform 1 0 15548 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_180
timestamp 1704896540
transform 1 0 17112 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_188
timestamp 1704896540
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1704896540
transform 1 0 18492 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_200
timestamp 1704896540
transform 1 0 18952 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_212
timestamp 1704896540
transform 1 0 20056 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_224
timestamp 1704896540
transform 1 0 21160 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_232
timestamp 1704896540
transform 1 0 21896 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 1704896540
transform 1 0 23092 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1704896540
transform 1 0 23644 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1704896540
transform 1 0 23828 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1704896540
transform 1 0 24932 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 1704896540
transform 1 0 26036 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_289
timestamp 1704896540
transform 1 0 27140 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_297
timestamp 1704896540
transform 1 0 27876 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_3
timestamp 1704896540
transform 1 0 828 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_11
timestamp 1704896540
transform 1 0 1564 0 -1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_17
timestamp 1704896540
transform 1 0 2116 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_33
timestamp 1704896540
transform 1 0 3588 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_45
timestamp 1704896540
transform 1 0 4692 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1704896540
transform 1 0 5612 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_77
timestamp 1704896540
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_109
timestamp 1704896540
transform 1 0 10580 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_126
timestamp 1704896540
transform 1 0 12144 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_151
timestamp 1704896540
transform 1 0 14444 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 1704896540
transform 1 0 15364 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1704896540
transform 1 0 15916 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_169
timestamp 1704896540
transform 1 0 16100 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_173
timestamp 1704896540
transform 1 0 16468 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_185
timestamp 1704896540
transform 1 0 17572 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_215
timestamp 1704896540
transform 1 0 20332 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1704896540
transform 1 0 21068 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_225
timestamp 1704896540
transform 1 0 21252 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_234
timestamp 1704896540
transform 1 0 22080 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_240
timestamp 1704896540
transform 1 0 22632 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 1704896540
transform 1 0 23460 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 1704896540
transform 1 0 24564 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 1704896540
transform 1 0 25668 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1704896540
transform 1 0 26220 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1704896540
transform 1 0 26404 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_293
timestamp 1704896540
transform 1 0 27508 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_299
timestamp 1704896540
transform 1 0 28060 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_3
timestamp 1704896540
transform 1 0 828 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_22
timestamp 1704896540
transform 1 0 2576 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_49
timestamp 1704896540
transform 1 0 5060 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_80
timestamp 1704896540
transform 1 0 7912 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_92
timestamp 1704896540
transform 1 0 9016 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_104
timestamp 1704896540
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_109
timestamp 1704896540
transform 1 0 10580 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_117
timestamp 1704896540
transform 1 0 11316 0 1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_125
timestamp 1704896540
transform 1 0 12052 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_137
timestamp 1704896540
transform 1 0 13156 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_141
timestamp 1704896540
transform 1 0 13524 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_145
timestamp 1704896540
transform 1 0 13892 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_149
timestamp 1704896540
transform 1 0 14260 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 1704896540
transform 1 0 18308 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_197
timestamp 1704896540
transform 1 0 18676 0 1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_203
timestamp 1704896540
transform 1 0 19228 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_215
timestamp 1704896540
transform 1 0 20332 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_219
timestamp 1704896540
transform 1 0 20700 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_231
timestamp 1704896540
transform 1 0 21804 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_238
timestamp 1704896540
transform 1 0 22448 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_249
timestamp 1704896540
transform 1 0 23460 0 1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_257
timestamp 1704896540
transform 1 0 24196 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_269
timestamp 1704896540
transform 1 0 25300 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_281
timestamp 1704896540
transform 1 0 26404 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_293
timestamp 1704896540
transform 1 0 27508 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_299
timestamp 1704896540
transform 1 0 28060 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_3
timestamp 1704896540
transform 1 0 828 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_9
timestamp 1704896540
transform 1 0 1380 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_14
timestamp 1704896540
transform 1 0 1840 0 -1 22304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_24
timestamp 1704896540
transform 1 0 2760 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_36
timestamp 1704896540
transform 1 0 3864 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_47
timestamp 1704896540
transform 1 0 4876 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1704896540
transform 1 0 5612 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_57
timestamp 1704896540
transform 1 0 5796 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_65
timestamp 1704896540
transform 1 0 6532 0 -1 22304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_72
timestamp 1704896540
transform 1 0 7176 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_89
timestamp 1704896540
transform 1 0 8740 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_99
timestamp 1704896540
transform 1 0 9660 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_107
timestamp 1704896540
transform 1 0 10396 0 -1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_121
timestamp 1704896540
transform 1 0 11684 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_133
timestamp 1704896540
transform 1 0 12788 0 -1 22304
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_144
timestamp 1704896540
transform 1 0 13800 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_156
timestamp 1704896540
transform 1 0 14904 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_169
timestamp 1704896540
transform 1 0 16100 0 -1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_177
timestamp 1704896540
transform 1 0 16836 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_189
timestamp 1704896540
transform 1 0 17940 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_197
timestamp 1704896540
transform 1 0 18676 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_219
timestamp 1704896540
transform 1 0 20700 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1704896540
transform 1 0 21068 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_225
timestamp 1704896540
transform 1 0 21252 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_244
timestamp 1704896540
transform 1 0 23000 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_252
timestamp 1704896540
transform 1 0 23736 0 -1 22304
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 1704896540
transform 1 0 24564 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 1704896540
transform 1 0 25668 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1704896540
transform 1 0 26220 0 -1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1704896540
transform 1 0 26404 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_293
timestamp 1704896540
transform 1 0 27508 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_299
timestamp 1704896540
transform 1 0 28060 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_3
timestamp 1704896540
transform 1 0 828 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_11
timestamp 1704896540
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_21
timestamp 1704896540
transform 1 0 2484 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1704896540
transform 1 0 3036 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_39
timestamp 1704896540
transform 1 0 4140 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_56
timestamp 1704896540
transform 1 0 5704 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_62
timestamp 1704896540
transform 1 0 6256 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_69
timestamp 1704896540
transform 1 0 6900 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_75
timestamp 1704896540
transform 1 0 7452 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_81
timestamp 1704896540
transform 1 0 8004 0 1 22304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_92
timestamp 1704896540
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_104
timestamp 1704896540
transform 1 0 10120 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_112
timestamp 1704896540
transform 1 0 10856 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_117
timestamp 1704896540
transform 1 0 11316 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_121
timestamp 1704896540
transform 1 0 11684 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_127
timestamp 1704896540
transform 1 0 12236 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_135
timestamp 1704896540
transform 1 0 12972 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1704896540
transform 1 0 13340 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_141
timestamp 1704896540
transform 1 0 13524 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_151
timestamp 1704896540
transform 1 0 14444 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_159
timestamp 1704896540
transform 1 0 15180 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_167
timestamp 1704896540
transform 1 0 15916 0 1 22304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_175
timestamp 1704896540
transform 1 0 16652 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_187
timestamp 1704896540
transform 1 0 17756 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1704896540
transform 1 0 18492 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_204
timestamp 1704896540
transform 1 0 19320 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_229
timestamp 1704896540
transform 1 0 21620 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_233
timestamp 1704896540
transform 1 0 21988 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_241
timestamp 1704896540
transform 1 0 22724 0 1 22304
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_270
timestamp 1704896540
transform 1 0 25392 0 1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_282
timestamp 1704896540
transform 1 0 26496 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_294
timestamp 1704896540
transform 1 0 27600 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_3
timestamp 1704896540
transform 1 0 828 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_12
timestamp 1704896540
transform 1 0 1656 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_18
timestamp 1704896540
transform 1 0 2208 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_26
timestamp 1704896540
transform 1 0 2944 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_35
timestamp 1704896540
transform 1 0 3772 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_41
timestamp 1704896540
transform 1 0 4324 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_45
timestamp 1704896540
transform 1 0 4692 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_53
timestamp 1704896540
transform 1 0 5428 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_57
timestamp 1704896540
transform 1 0 5796 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_63
timestamp 1704896540
transform 1 0 6348 0 -1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_71
timestamp 1704896540
transform 1 0 7084 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_86
timestamp 1704896540
transform 1 0 8464 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_121
timestamp 1704896540
transform 1 0 11684 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_140
timestamp 1704896540
transform 1 0 13432 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_146
timestamp 1704896540
transform 1 0 13984 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_162
timestamp 1704896540
transform 1 0 15456 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_169
timestamp 1704896540
transform 1 0 16100 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_173
timestamp 1704896540
transform 1 0 16468 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_184
timestamp 1704896540
transform 1 0 17480 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_191
timestamp 1704896540
transform 1 0 18124 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_202
timestamp 1704896540
transform 1 0 19136 0 -1 23392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_208
timestamp 1704896540
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_220
timestamp 1704896540
transform 1 0 20792 0 -1 23392
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_232
timestamp 1704896540
transform 1 0 21896 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_244
timestamp 1704896540
transform 1 0 23000 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_256
timestamp 1704896540
transform 1 0 24104 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_268
timestamp 1704896540
transform 1 0 25208 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1704896540
transform 1 0 26404 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_293
timestamp 1704896540
transform 1 0 27508 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_299
timestamp 1704896540
transform 1 0 28060 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_26
timestamp 1704896540
transform 1 0 2944 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_29
timestamp 1704896540
transform 1 0 3220 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_45
timestamp 1704896540
transform 1 0 4692 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_53
timestamp 1704896540
transform 1 0 5428 0 1 23392
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1704896540
transform 1 0 6532 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1704896540
transform 1 0 7636 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1704896540
transform 1 0 8188 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_85
timestamp 1704896540
transform 1 0 8372 0 1 23392
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_99
timestamp 1704896540
transform 1 0 9660 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_111
timestamp 1704896540
transform 1 0 10764 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_123
timestamp 1704896540
transform 1 0 11868 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_127
timestamp 1704896540
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_131
timestamp 1704896540
transform 1 0 12604 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1704896540
transform 1 0 13340 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_141
timestamp 1704896540
transform 1 0 13524 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_145
timestamp 1704896540
transform 1 0 13892 0 1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_149
timestamp 1704896540
transform 1 0 14260 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_161
timestamp 1704896540
transform 1 0 15364 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_192
timestamp 1704896540
transform 1 0 18216 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_224
timestamp 1704896540
transform 1 0 21160 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_228
timestamp 1704896540
transform 1 0 21528 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_246
timestamp 1704896540
transform 1 0 23184 0 1 23392
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_263
timestamp 1704896540
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_275
timestamp 1704896540
transform 1 0 25852 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_287
timestamp 1704896540
transform 1 0 26956 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_299
timestamp 1704896540
transform 1 0 28060 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_3
timestamp 1704896540
transform 1 0 828 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_9
timestamp 1704896540
transform 1 0 1380 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_54
timestamp 1704896540
transform 1 0 5520 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_70
timestamp 1704896540
transform 1 0 6992 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_85
timestamp 1704896540
transform 1 0 8372 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_91
timestamp 1704896540
transform 1 0 8924 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_103
timestamp 1704896540
transform 1 0 10028 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_107
timestamp 1704896540
transform 1 0 10396 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1704896540
transform 1 0 10764 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_123
timestamp 1704896540
transform 1 0 11868 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_127
timestamp 1704896540
transform 1 0 12236 0 -1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_131
timestamp 1704896540
transform 1 0 12604 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_148
timestamp 1704896540
transform 1 0 14168 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_156
timestamp 1704896540
transform 1 0 14904 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_162
timestamp 1704896540
transform 1 0 15456 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_186
timestamp 1704896540
transform 1 0 17664 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_196
timestamp 1704896540
transform 1 0 18584 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_206
timestamp 1704896540
transform 1 0 19504 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_210
timestamp 1704896540
transform 1 0 19872 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_220
timestamp 1704896540
transform 1 0 20792 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_225
timestamp 1704896540
transform 1 0 21252 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_270
timestamp 1704896540
transform 1 0 25392 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_278
timestamp 1704896540
transform 1 0 26128 0 -1 24480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1704896540
transform 1 0 26404 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_293
timestamp 1704896540
transform 1 0 27508 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_299
timestamp 1704896540
transform 1 0 28060 0 -1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1704896540
transform 1 0 828 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1704896540
transform 1 0 1932 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1704896540
transform 1 0 3036 0 1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1704896540
transform 1 0 3220 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1704896540
transform 1 0 4324 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_53
timestamp 1704896540
transform 1 0 5428 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_75
timestamp 1704896540
transform 1 0 7452 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1704896540
transform 1 0 8188 0 1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1704896540
transform 1 0 8372 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_97
timestamp 1704896540
transform 1 0 9476 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_124
timestamp 1704896540
transform 1 0 11960 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_134
timestamp 1704896540
transform 1 0 12880 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_141
timestamp 1704896540
transform 1 0 13524 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_162
timestamp 1704896540
transform 1 0 15456 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_166
timestamp 1704896540
transform 1 0 15824 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_187
timestamp 1704896540
transform 1 0 17756 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1704896540
transform 1 0 18492 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_210
timestamp 1704896540
transform 1 0 19872 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_218
timestamp 1704896540
transform 1 0 20608 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_229
timestamp 1704896540
transform 1 0 21620 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_241
timestamp 1704896540
transform 1 0 22724 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_249
timestamp 1704896540
transform 1 0 23460 0 1 24480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1704896540
transform 1 0 23828 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1704896540
transform 1 0 24932 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1704896540
transform 1 0 26036 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_289
timestamp 1704896540
transform 1 0 27140 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_297
timestamp 1704896540
transform 1 0 27876 0 1 24480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1704896540
transform 1 0 828 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_15
timestamp 1704896540
transform 1 0 1932 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_23
timestamp 1704896540
transform 1 0 2668 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_39
timestamp 1704896540
transform 1 0 4140 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_48
timestamp 1704896540
transform 1 0 4968 0 -1 25568
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1704896540
transform 1 0 5796 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_69
timestamp 1704896540
transform 1 0 6900 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_77
timestamp 1704896540
transform 1 0 7636 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_85
timestamp 1704896540
transform 1 0 8372 0 -1 25568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_94
timestamp 1704896540
transform 1 0 9200 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_106
timestamp 1704896540
transform 1 0 10304 0 -1 25568
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1704896540
transform 1 0 10948 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_125
timestamp 1704896540
transform 1 0 12052 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_133
timestamp 1704896540
transform 1 0 12788 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_141
timestamp 1704896540
transform 1 0 13524 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_147
timestamp 1704896540
transform 1 0 14076 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_153
timestamp 1704896540
transform 1 0 14628 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1704896540
transform 1 0 15364 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1704896540
transform 1 0 15916 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_169
timestamp 1704896540
transform 1 0 16100 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_173
timestamp 1704896540
transform 1 0 16468 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_181
timestamp 1704896540
transform 1 0 17204 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_189
timestamp 1704896540
transform 1 0 17940 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_203
timestamp 1704896540
transform 1 0 19228 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_221
timestamp 1704896540
transform 1 0 20884 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_233
timestamp 1704896540
transform 1 0 21988 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_241
timestamp 1704896540
transform 1 0 22724 0 -1 25568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_259
timestamp 1704896540
transform 1 0 24380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_271
timestamp 1704896540
transform 1 0 25484 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1704896540
transform 1 0 26220 0 -1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1704896540
transform 1 0 26404 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_293
timestamp 1704896540
transform 1 0 27508 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_299
timestamp 1704896540
transform 1 0 28060 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_3
timestamp 1704896540
transform 1 0 828 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_11
timestamp 1704896540
transform 1 0 1564 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_37
timestamp 1704896540
transform 1 0 3956 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_56
timestamp 1704896540
transform 1 0 5704 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_73
timestamp 1704896540
transform 1 0 7268 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_81
timestamp 1704896540
transform 1 0 8004 0 1 25568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_91
timestamp 1704896540
transform 1 0 8924 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_103
timestamp 1704896540
transform 1 0 10028 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_127
timestamp 1704896540
transform 1 0 12236 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_138
timestamp 1704896540
transform 1 0 13248 0 1 25568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1704896540
transform 1 0 13524 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_153
timestamp 1704896540
transform 1 0 14628 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_163
timestamp 1704896540
transform 1 0 15548 0 1 25568
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_172
timestamp 1704896540
transform 1 0 16376 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_184
timestamp 1704896540
transform 1 0 17480 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_192
timestamp 1704896540
transform 1 0 18216 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_213
timestamp 1704896540
transform 1 0 20148 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_222
timestamp 1704896540
transform 1 0 20976 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_242
timestamp 1704896540
transform 1 0 22816 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_250
timestamp 1704896540
transform 1 0 23552 0 1 25568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1704896540
transform 1 0 23828 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1704896540
transform 1 0 24932 0 1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1704896540
transform 1 0 26036 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_289
timestamp 1704896540
transform 1 0 27140 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_297
timestamp 1704896540
transform 1 0 27876 0 1 25568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1704896540
transform 1 0 828 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1704896540
transform 1 0 1932 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1704896540
transform 1 0 3036 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_39
timestamp 1704896540
transform 1 0 4140 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_46
timestamp 1704896540
transform 1 0 4784 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_54
timestamp 1704896540
transform 1 0 5520 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_57
timestamp 1704896540
transform 1 0 5796 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_66
timestamp 1704896540
transform 1 0 6624 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_72
timestamp 1704896540
transform 1 0 7176 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_83
timestamp 1704896540
transform 1 0 8188 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_91
timestamp 1704896540
transform 1 0 8924 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_100
timestamp 1704896540
transform 1 0 9752 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_108
timestamp 1704896540
transform 1 0 10488 0 -1 26656
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1704896540
transform 1 0 10948 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_125
timestamp 1704896540
transform 1 0 12052 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_133
timestamp 1704896540
transform 1 0 12788 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_141
timestamp 1704896540
transform 1 0 13524 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_149
timestamp 1704896540
transform 1 0 14260 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_159
timestamp 1704896540
transform 1 0 15180 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1704896540
transform 1 0 15916 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_169
timestamp 1704896540
transform 1 0 16100 0 -1 26656
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_190
timestamp 1704896540
transform 1 0 18032 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_202
timestamp 1704896540
transform 1 0 19136 0 -1 26656
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1704896540
transform 1 0 21252 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1704896540
transform 1 0 22356 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1704896540
transform 1 0 23460 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1704896540
transform 1 0 24564 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 1704896540
transform 1 0 25668 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1704896540
transform 1 0 26220 0 -1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1704896540
transform 1 0 26404 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_293
timestamp 1704896540
transform 1 0 27508 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_299
timestamp 1704896540
transform 1 0 28060 0 -1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1704896540
transform 1 0 828 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_15
timestamp 1704896540
transform 1 0 1932 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_23
timestamp 1704896540
transform 1 0 2668 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1704896540
transform 1 0 3036 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_42
timestamp 1704896540
transform 1 0 4416 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_63
timestamp 1704896540
transform 1 0 6348 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_71
timestamp 1704896540
transform 1 0 7084 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_80
timestamp 1704896540
transform 1 0 7912 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_85
timestamp 1704896540
transform 1 0 8372 0 1 26656
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_93
timestamp 1704896540
transform 1 0 9108 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_105
timestamp 1704896540
transform 1 0 10212 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_113
timestamp 1704896540
transform 1 0 10948 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_137
timestamp 1704896540
transform 1 0 13156 0 1 26656
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1704896540
transform 1 0 13524 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_186
timestamp 1704896540
transform 1 0 17664 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1704896540
transform 1 0 18492 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_197
timestamp 1704896540
transform 1 0 18676 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_217
timestamp 1704896540
transform 1 0 20516 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_234
timestamp 1704896540
transform 1 0 22080 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_248
timestamp 1704896540
transform 1 0 23368 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_253
timestamp 1704896540
transform 1 0 23828 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_257
timestamp 1704896540
transform 1 0 24196 0 1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_266
timestamp 1704896540
transform 1 0 25024 0 1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_278
timestamp 1704896540
transform 1 0 26128 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_290
timestamp 1704896540
transform 1 0 27232 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_298
timestamp 1704896540
transform 1 0 27968 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_3
timestamp 1704896540
transform 1 0 828 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_15
timestamp 1704896540
transform 1 0 1932 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_41
timestamp 1704896540
transform 1 0 4324 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_60
timestamp 1704896540
transform 1 0 6072 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_88
timestamp 1704896540
transform 1 0 8648 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_113
timestamp 1704896540
transform 1 0 10948 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_166
timestamp 1704896540
transform 1 0 15824 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_225
timestamp 1704896540
transform 1 0 21252 0 -1 27744
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_260
timestamp 1704896540
transform 1 0 24472 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_272
timestamp 1704896540
transform 1 0 25576 0 -1 27744
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1704896540
transform 1 0 26404 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_293
timestamp 1704896540
transform 1 0 27508 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_299
timestamp 1704896540
transform 1 0 28060 0 -1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1704896540
transform 1 0 828 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1704896540
transform 1 0 1932 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1704896540
transform 1 0 3036 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1704896540
transform 1 0 3220 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1704896540
transform 1 0 4324 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_53
timestamp 1704896540
transform 1 0 5428 0 1 27744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_57
timestamp 1704896540
transform 1 0 5796 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_69
timestamp 1704896540
transform 1 0 6900 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_81
timestamp 1704896540
transform 1 0 8004 0 1 27744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1704896540
transform 1 0 8372 0 1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1704896540
transform 1 0 9476 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_109
timestamp 1704896540
transform 1 0 10580 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_113
timestamp 1704896540
transform 1 0 10948 0 1 27744
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_119
timestamp 1704896540
transform 1 0 11500 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_131
timestamp 1704896540
transform 1 0 12604 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1704896540
transform 1 0 13340 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1704896540
transform 1 0 13524 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_153
timestamp 1704896540
transform 1 0 14628 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_161
timestamp 1704896540
transform 1 0 15364 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_167
timestamp 1704896540
transform 1 0 15916 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_169
timestamp 1704896540
transform 1 0 16100 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_181
timestamp 1704896540
transform 1 0 17204 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_188
timestamp 1704896540
transform 1 0 17848 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_197
timestamp 1704896540
transform 1 0 18676 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_217
timestamp 1704896540
transform 1 0 20516 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_223
timestamp 1704896540
transform 1 0 21068 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_225
timestamp 1704896540
transform 1 0 21252 0 1 27744
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_232
timestamp 1704896540
transform 1 0 21896 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_244
timestamp 1704896540
transform 1 0 23000 0 1 27744
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_256
timestamp 1704896540
transform 1 0 24104 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_268
timestamp 1704896540
transform 1 0 25208 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_272
timestamp 1704896540
transform 1 0 25576 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_279
timestamp 1704896540
transform 1 0 26220 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_281
timestamp 1704896540
transform 1 0 26404 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_293
timestamp 1704896540
transform 1 0 27508 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_299
timestamp 1704896540
transform 1 0 28060 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19228 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform 1 0 20240 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform 1 0 22356 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform -1 0 25024 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform -1 0 2760 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 3956 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform 1 0 16652 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform -1 0 11684 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1704896540
transform -1 0 16836 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1704896540
transform -1 0 17388 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1704896540
transform -1 0 20240 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1704896540
transform -1 0 15548 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1704896540
transform -1 0 19228 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1704896540
transform -1 0 13064 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1704896540
transform -1 0 17664 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1704896540
transform 1 0 3496 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1704896540
transform 1 0 10948 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1704896540
transform 1 0 25668 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1704896540
transform 1 0 23828 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1704896540
transform 1 0 21620 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform 1 0 20240 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1704896540
transform -1 0 17848 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13984 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1704896540
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1704896540
transform -1 0 28428 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1704896540
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1704896540
transform -1 0 28428 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1704896540
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1704896540
transform -1 0 28428 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1704896540
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1704896540
transform -1 0 28428 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1704896540
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1704896540
transform -1 0 28428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1704896540
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1704896540
transform -1 0 28428 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1704896540
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1704896540
transform -1 0 28428 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1704896540
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1704896540
transform -1 0 28428 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1704896540
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1704896540
transform -1 0 28428 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1704896540
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1704896540
transform -1 0 28428 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1704896540
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1704896540
transform -1 0 28428 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1704896540
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1704896540
transform -1 0 28428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1704896540
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1704896540
transform -1 0 28428 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1704896540
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1704896540
transform -1 0 28428 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1704896540
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1704896540
transform -1 0 28428 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1704896540
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1704896540
transform -1 0 28428 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1704896540
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1704896540
transform -1 0 28428 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1704896540
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1704896540
transform -1 0 28428 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1704896540
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1704896540
transform -1 0 28428 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1704896540
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1704896540
transform -1 0 28428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1704896540
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1704896540
transform -1 0 28428 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1704896540
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1704896540
transform -1 0 28428 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1704896540
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1704896540
transform -1 0 28428 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1704896540
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1704896540
transform -1 0 28428 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1704896540
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1704896540
transform -1 0 28428 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1704896540
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1704896540
transform -1 0 28428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1704896540
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1704896540
transform -1 0 28428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1704896540
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1704896540
transform -1 0 28428 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1704896540
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1704896540
transform -1 0 28428 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1704896540
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1704896540
transform -1 0 28428 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1704896540
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1704896540
transform -1 0 28428 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1704896540
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1704896540
transform -1 0 28428 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1704896540
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1704896540
transform -1 0 28428 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1704896540
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1704896540
transform -1 0 28428 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1704896540
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1704896540
transform -1 0 28428 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1704896540
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1704896540
transform -1 0 28428 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1704896540
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1704896540
transform -1 0 28428 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1704896540
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1704896540
transform -1 0 28428 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1704896540
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1704896540
transform -1 0 28428 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1704896540
transform 1 0 552 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1704896540
transform -1 0 28428 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1704896540
transform 1 0 552 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1704896540
transform -1 0 28428 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1704896540
transform 1 0 552 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1704896540
transform -1 0 28428 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1704896540
transform 1 0 552 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1704896540
transform -1 0 28428 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1704896540
transform 1 0 552 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1704896540
transform -1 0 28428 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1704896540
transform 1 0 552 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1704896540
transform -1 0 28428 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1704896540
transform 1 0 552 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1704896540
transform -1 0 28428 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1704896540
transform 1 0 552 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1704896540
transform -1 0 28428 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1704896540
transform 1 0 552 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1704896540
transform -1 0 28428 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1704896540
transform 1 0 552 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1704896540
transform -1 0 28428 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1704896540
transform 1 0 552 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1704896540
transform -1 0 28428 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1704896540
transform 1 0 552 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1704896540
transform -1 0 28428 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1704896540
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1704896540
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1704896540
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1704896540
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1704896540
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1704896540
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1704896540
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1704896540
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1704896540
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1704896540
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1704896540
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1704896540
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1704896540
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1704896540
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1704896540
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1704896540
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1704896540
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1704896540
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1704896540
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1704896540
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1704896540
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1704896540
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1704896540
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1704896540
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1704896540
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1704896540
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1704896540
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1704896540
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1704896540
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1704896540
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1704896540
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1704896540
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1704896540
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1704896540
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1704896540
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1704896540
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1704896540
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1704896540
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1704896540
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1704896540
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1704896540
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1704896540
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1704896540
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1704896540
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1704896540
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1704896540
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1704896540
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1704896540
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1704896540
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1704896540
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1704896540
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1704896540
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1704896540
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1704896540
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1704896540
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1704896540
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1704896540
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1704896540
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1704896540
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1704896540
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1704896540
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1704896540
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1704896540
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1704896540
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1704896540
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1704896540
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1704896540
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1704896540
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1704896540
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1704896540
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1704896540
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1704896540
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1704896540
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1704896540
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1704896540
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1704896540
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1704896540
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1704896540
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1704896540
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1704896540
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1704896540
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1704896540
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1704896540
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1704896540
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1704896540
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1704896540
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1704896540
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1704896540
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1704896540
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1704896540
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1704896540
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1704896540
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1704896540
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1704896540
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1704896540
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1704896540
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1704896540
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1704896540
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1704896540
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1704896540
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1704896540
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1704896540
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1704896540
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1704896540
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1704896540
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1704896540
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1704896540
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1704896540
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1704896540
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1704896540
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1704896540
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1704896540
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1704896540
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1704896540
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1704896540
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1704896540
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1704896540
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1704896540
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1704896540
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1704896540
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1704896540
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1704896540
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1704896540
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1704896540
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1704896540
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1704896540
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1704896540
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1704896540
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1704896540
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1704896540
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1704896540
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1704896540
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1704896540
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1704896540
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1704896540
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1704896540
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1704896540
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1704896540
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1704896540
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1704896540
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1704896540
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1704896540
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1704896540
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1704896540
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1704896540
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1704896540
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1704896540
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1704896540
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1704896540
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1704896540
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1704896540
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1704896540
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1704896540
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1704896540
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1704896540
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1704896540
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1704896540
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1704896540
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1704896540
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1704896540
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1704896540
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1704896540
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1704896540
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1704896540
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1704896540
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1704896540
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1704896540
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1704896540
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1704896540
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1704896540
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1704896540
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1704896540
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1704896540
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1704896540
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1704896540
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1704896540
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1704896540
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1704896540
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1704896540
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1704896540
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1704896540
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1704896540
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1704896540
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1704896540
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1704896540
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1704896540
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1704896540
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1704896540
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1704896540
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1704896540
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1704896540
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1704896540
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1704896540
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1704896540
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1704896540
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1704896540
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1704896540
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1704896540
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1704896540
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1704896540
transform 1 0 5704 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1704896540
transform 1 0 10856 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1704896540
transform 1 0 16008 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1704896540
transform 1 0 21160 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1704896540
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1704896540
transform 1 0 3128 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1704896540
transform 1 0 8280 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1704896540
transform 1 0 13432 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1704896540
transform 1 0 18584 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1704896540
transform 1 0 23736 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1704896540
transform 1 0 5704 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1704896540
transform 1 0 10856 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1704896540
transform 1 0 16008 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1704896540
transform 1 0 21160 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1704896540
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1704896540
transform 1 0 3128 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1704896540
transform 1 0 8280 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1704896540
transform 1 0 13432 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1704896540
transform 1 0 18584 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1704896540
transform 1 0 23736 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1704896540
transform 1 0 5704 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1704896540
transform 1 0 10856 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1704896540
transform 1 0 16008 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1704896540
transform 1 0 21160 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1704896540
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1704896540
transform 1 0 3128 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1704896540
transform 1 0 8280 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1704896540
transform 1 0 13432 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1704896540
transform 1 0 18584 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1704896540
transform 1 0 23736 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1704896540
transform 1 0 5704 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1704896540
transform 1 0 10856 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1704896540
transform 1 0 16008 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1704896540
transform 1 0 21160 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1704896540
transform 1 0 26312 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1704896540
transform 1 0 3128 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1704896540
transform 1 0 8280 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1704896540
transform 1 0 13432 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1704896540
transform 1 0 18584 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1704896540
transform 1 0 23736 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1704896540
transform 1 0 5704 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1704896540
transform 1 0 10856 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1704896540
transform 1 0 16008 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1704896540
transform 1 0 21160 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1704896540
transform 1 0 26312 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1704896540
transform 1 0 3128 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1704896540
transform 1 0 8280 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1704896540
transform 1 0 13432 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1704896540
transform 1 0 18584 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1704896540
transform 1 0 23736 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1704896540
transform 1 0 5704 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1704896540
transform 1 0 10856 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1704896540
transform 1 0 16008 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1704896540
transform 1 0 21160 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1704896540
transform 1 0 26312 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1704896540
transform 1 0 3128 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1704896540
transform 1 0 5704 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1704896540
transform 1 0 8280 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1704896540
transform 1 0 10856 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1704896540
transform 1 0 13432 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1704896540
transform 1 0 16008 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1704896540
transform 1 0 18584 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1704896540
transform 1 0 21160 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1704896540
transform 1 0 23736 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1704896540
transform 1 0 26312 0 1 27744
box -38 -48 130 592
<< labels >>
flabel metal4 s 7360 496 7680 28336 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 14329 496 14649 28336 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 21298 496 21618 28336 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 28267 496 28587 28336 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3876 496 4196 28336 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 10845 496 11165 28336 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 17814 496 18134 28336 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 24783 496 25103 28336 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 27618 28600 27674 29000 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal2 s 25594 28600 25650 29000 0 FreeSans 224 90 0 0 rst_n
port 3 nsew signal input
flabel metal2 s 23570 28600 23626 29000 0 FreeSans 224 90 0 0 ui_in[0]
port 4 nsew signal input
flabel metal2 s 21546 28600 21602 29000 0 FreeSans 224 90 0 0 ui_in[1]
port 5 nsew signal input
flabel metal2 s 19522 28600 19578 29000 0 FreeSans 224 90 0 0 ui_in[2]
port 6 nsew signal input
flabel metal2 s 17498 28600 17554 29000 0 FreeSans 224 90 0 0 ui_in[3]
port 7 nsew signal input
flabel metal2 s 15474 28600 15530 29000 0 FreeSans 224 90 0 0 uo_out[0]
port 8 nsew signal tristate
flabel metal2 s 13450 28600 13506 29000 0 FreeSans 224 90 0 0 uo_out[1]
port 9 nsew signal tristate
flabel metal2 s 11426 28600 11482 29000 0 FreeSans 224 90 0 0 uo_out[2]
port 10 nsew signal tristate
flabel metal2 s 9402 28600 9458 29000 0 FreeSans 224 90 0 0 uo_out[3]
port 11 nsew signal tristate
flabel metal2 s 7378 28600 7434 29000 0 FreeSans 224 90 0 0 uo_out[4]
port 12 nsew signal tristate
flabel metal2 s 5354 28600 5410 29000 0 FreeSans 224 90 0 0 uo_out[5]
port 13 nsew signal tristate
flabel metal2 s 3330 28600 3386 29000 0 FreeSans 224 90 0 0 uo_out[6]
port 14 nsew signal tristate
flabel metal2 s 1306 28600 1362 29000 0 FreeSans 224 90 0 0 uo_out[7]
port 15 nsew signal tristate
rlabel via1 14569 27744 14569 27744 0 VGND
rlabel metal1 14490 28288 14490 28288 0 VPWR
rlabel via1 9701 23222 9701 23222 0 _0000_
rlabel metal1 10764 24378 10764 24378 0 _0001_
rlabel via1 6030 26894 6030 26894 0 _0002_
rlabel metal2 2622 27302 2622 27302 0 _0003_
rlabel metal2 2438 25602 2438 25602 0 _0004_
rlabel metal1 19186 25738 19186 25738 0 _0005_
rlabel metal2 21758 25602 21758 25602 0 _0006_
rlabel metal2 19642 25126 19642 25126 0 _0007_
rlabel metal2 24518 24038 24518 24038 0 _0008_
rlabel metal2 24334 22338 24334 22338 0 _0009_
rlabel metal2 23230 19686 23230 19686 0 _0010_
rlabel viali 18993 19210 18993 19210 0 _0011_
rlabel metal1 19810 17782 19810 17782 0 _0012_
rlabel metal1 19044 21658 19044 21658 0 _0013_
rlabel metal2 20194 15810 20194 15810 0 _0014_
rlabel metal1 21482 15470 21482 15470 0 _0015_
rlabel metal2 22310 14008 22310 14008 0 _0016_
rlabel via1 20934 11662 20934 11662 0 _0017_
rlabel metal1 17802 12954 17802 12954 0 _0018_
rlabel metal1 11730 10778 11730 10778 0 _0019_
rlabel metal1 11725 12682 11725 12682 0 _0020_
rlabel metal1 17346 11186 17346 11186 0 _0021_
rlabel metal1 5024 11662 5024 11662 0 _0022_
rlabel via1 1789 13362 1789 13362 0 _0023_
rlabel via1 1789 16014 1789 16014 0 _0024_
rlabel metal2 3726 17510 3726 17510 0 _0025_
rlabel metal2 6302 14722 6302 14722 0 _0026_
rlabel via1 7410 10506 7410 10506 0 _0027_
rlabel via1 10161 10506 10161 10506 0 _0028_
rlabel metal1 8183 10166 8183 10166 0 _0029_
rlabel metal1 11408 14042 11408 14042 0 _0030_
rlabel metal1 11311 19958 11311 19958 0 _0031_
rlabel metal1 10779 17782 10779 17782 0 _0032_
rlabel via1 12829 14518 12829 14518 0 _0033_
rlabel metal1 10860 16014 10860 16014 0 _0034_
rlabel metal2 17066 17476 17066 17476 0 _0035_
rlabel via1 1145 23562 1145 23562 0 _0036_
rlabel metal1 2438 23834 2438 23834 0 _0037_
rlabel metal2 3542 23766 3542 23766 0 _0038_
rlabel metal2 4738 25602 4738 25602 0 _0039_
rlabel metal2 5842 20978 5842 20978 0 _0040_
rlabel metal1 3342 21386 3342 21386 0 _0041_
rlabel metal2 4922 19074 4922 19074 0 _0042_
rlabel metal1 2019 18190 2019 18190 0 _0043_
rlabel via1 1605 19958 1605 19958 0 _0044_
rlabel metal1 1559 21454 1559 21454 0 _0045_
rlabel metal2 14858 21250 14858 21250 0 _0046_
rlabel metal1 15440 26826 15440 26826 0 _0047_
rlabel metal1 16320 27506 16320 27506 0 _0048_
rlabel metal1 15900 24310 15900 24310 0 _0049_
rlabel metal1 16314 24650 16314 24650 0 _0050_
rlabel metal1 16468 26010 16468 26010 0 _0051_
rlabel metal2 12006 19074 12006 19074 0 _0052_
rlabel metal1 11495 16694 11495 16694 0 _0053_
rlabel metal1 15870 17578 15870 17578 0 _0054_
rlabel metal1 14260 18938 14260 18938 0 _0055_
rlabel via1 12829 20978 12829 20978 0 _0056_
rlabel metal1 14398 21046 14398 21046 0 _0057_
rlabel metal1 13570 22474 13570 22474 0 _0058_
rlabel metal1 12834 16660 12834 16660 0 _0059_
rlabel metal1 12604 22746 12604 22746 0 _0060_
rlabel viali 13205 23154 13205 23154 0 _0061_
rlabel metal2 2438 23018 2438 23018 0 _0062_
rlabel metal1 8326 21454 8326 21454 0 _0063_
rlabel metal1 6440 24242 6440 24242 0 _0064_
rlabel metal1 4646 22032 4646 22032 0 _0065_
rlabel metal1 5060 18190 5060 18190 0 _0066_
rlabel metal1 7314 22678 7314 22678 0 _0067_
rlabel metal2 9338 20196 9338 20196 0 _0068_
rlabel metal2 8326 21760 8326 21760 0 _0069_
rlabel metal1 9430 22032 9430 22032 0 _0070_
rlabel via2 15870 22933 15870 22933 0 _0071_
rlabel metal2 12190 22950 12190 22950 0 _0072_
rlabel metal2 13662 22814 13662 22814 0 _0073_
rlabel metal1 10166 26452 10166 26452 0 _0074_
rlabel metal1 11868 23154 11868 23154 0 _0075_
rlabel metal1 8694 22644 8694 22644 0 _0076_
rlabel metal2 8786 22508 8786 22508 0 _0077_
rlabel metal1 13846 19720 13846 19720 0 _0078_
rlabel metal1 9108 20570 9108 20570 0 _0079_
rlabel metal1 9752 20570 9752 20570 0 _0080_
rlabel metal1 14076 20774 14076 20774 0 _0081_
rlabel metal1 11132 22066 11132 22066 0 _0082_
rlabel metal1 9154 22066 9154 22066 0 _0083_
rlabel metal1 13938 19958 13938 19958 0 _0084_
rlabel metal2 9614 21862 9614 21862 0 _0085_
rlabel metal1 10534 21386 10534 21386 0 _0086_
rlabel metal1 8740 23086 8740 23086 0 _0087_
rlabel metal1 10856 22542 10856 22542 0 _0088_
rlabel metal1 7222 20026 7222 20026 0 _0089_
rlabel metal1 7084 19890 7084 19890 0 _0090_
rlabel metal2 12558 26214 12558 26214 0 _0091_
rlabel metal1 12650 26350 12650 26350 0 _0092_
rlabel metal2 12374 25602 12374 25602 0 _0093_
rlabel metal2 12282 25942 12282 25942 0 _0094_
rlabel metal1 6716 25670 6716 25670 0 _0095_
rlabel metal1 5474 23562 5474 23562 0 _0096_
rlabel metal1 6210 23664 6210 23664 0 _0097_
rlabel metal2 6486 23834 6486 23834 0 _0098_
rlabel metal1 7406 24650 7406 24650 0 _0099_
rlabel metal1 6670 24786 6670 24786 0 _0100_
rlabel metal1 7084 24786 7084 24786 0 _0101_
rlabel metal1 7130 25806 7130 25806 0 _0102_
rlabel metal1 6486 26010 6486 26010 0 _0103_
rlabel metal2 6762 24514 6762 24514 0 _0104_
rlabel metal1 8142 23018 8142 23018 0 _0105_
rlabel metal2 7774 26792 7774 26792 0 _0106_
rlabel metal1 11638 25670 11638 25670 0 _0107_
rlabel metal1 11224 25806 11224 25806 0 _0108_
rlabel metal1 9982 25670 9982 25670 0 _0109_
rlabel metal1 8510 25466 8510 25466 0 _0110_
rlabel metal2 7958 25636 7958 25636 0 _0111_
rlabel metal2 7912 26418 7912 26418 0 _0112_
rlabel metal1 7360 26554 7360 26554 0 _0113_
rlabel metal1 7590 26248 7590 26248 0 _0114_
rlabel metal1 9844 26282 9844 26282 0 _0115_
rlabel metal1 11270 27098 11270 27098 0 _0116_
rlabel metal1 12788 26350 12788 26350 0 _0117_
rlabel metal1 7774 24174 7774 24174 0 _0118_
rlabel metal1 8510 24378 8510 24378 0 _0119_
rlabel metal1 9062 25466 9062 25466 0 _0120_
rlabel metal2 6118 26996 6118 26996 0 _0121_
rlabel metal1 8234 27540 8234 27540 0 _0122_
rlabel metal2 7866 27268 7866 27268 0 _0123_
rlabel metal1 8142 27404 8142 27404 0 _0124_
rlabel metal1 8740 27438 8740 27438 0 _0125_
rlabel metal1 10994 26894 10994 26894 0 _0126_
rlabel metal1 12742 26928 12742 26928 0 _0127_
rlabel metal1 12650 26860 12650 26860 0 _0128_
rlabel metal2 12466 24446 12466 24446 0 _0129_
rlabel metal2 7498 15334 7498 15334 0 _0130_
rlabel metal1 8648 15130 8648 15130 0 _0131_
rlabel metal2 12006 15130 12006 15130 0 _0132_
rlabel metal2 16146 14722 16146 14722 0 _0133_
rlabel metal1 12558 14960 12558 14960 0 _0134_
rlabel metal1 14536 14450 14536 14450 0 _0135_
rlabel metal1 13340 14926 13340 14926 0 _0136_
rlabel metal2 12098 17051 12098 17051 0 _0137_
rlabel metal1 15318 25942 15318 25942 0 _0138_
rlabel metal1 7498 21556 7498 21556 0 _0139_
rlabel metal1 5382 21046 5382 21046 0 _0140_
rlabel metal2 7130 20910 7130 20910 0 _0141_
rlabel metal1 9062 20332 9062 20332 0 _0142_
rlabel metal1 14030 22610 14030 22610 0 _0143_
rlabel metal1 14076 22746 14076 22746 0 _0144_
rlabel metal1 15502 23154 15502 23154 0 _0145_
rlabel metal1 9062 22950 9062 22950 0 _0146_
rlabel metal1 6210 13362 6210 13362 0 _0147_
rlabel metal1 9024 23290 9024 23290 0 _0148_
rlabel metal1 9384 23290 9384 23290 0 _0149_
rlabel metal1 9752 24718 9752 24718 0 _0150_
rlabel metal2 7774 21709 7774 21709 0 _0151_
rlabel metal1 14030 23664 14030 23664 0 _0152_
rlabel metal1 10994 24344 10994 24344 0 _0153_
rlabel metal1 10488 24242 10488 24242 0 _0154_
rlabel metal1 4508 26214 4508 26214 0 _0155_
rlabel metal1 4797 26554 4797 26554 0 _0156_
rlabel metal1 5336 26282 5336 26282 0 _0157_
rlabel metal2 3726 26180 3726 26180 0 _0158_
rlabel metal1 3680 26758 3680 26758 0 _0159_
rlabel metal1 3128 26894 3128 26894 0 _0160_
rlabel metal1 13340 18802 13340 18802 0 _0161_
rlabel metal1 2990 25296 2990 25296 0 _0162_
rlabel metal1 20148 21454 20148 21454 0 _0163_
rlabel metal1 20516 21930 20516 21930 0 _0164_
rlabel viali 20390 22542 20390 22542 0 _0165_
rlabel metal1 21574 22576 21574 22576 0 _0166_
rlabel metal1 20838 21522 20838 21522 0 _0167_
rlabel metal1 20930 18768 20930 18768 0 _0168_
rlabel metal1 19090 18802 19090 18802 0 _0169_
rlabel metal2 18446 25636 18446 25636 0 _0170_
rlabel metal1 21206 21658 21206 21658 0 _0171_
rlabel metal1 21528 24922 21528 24922 0 _0172_
rlabel metal1 21804 25330 21804 25330 0 _0173_
rlabel metal1 21068 19142 21068 19142 0 _0174_
rlabel metal2 22770 21386 22770 21386 0 _0175_
rlabel metal2 20562 24004 20562 24004 0 _0176_
rlabel metal1 19504 24378 19504 24378 0 _0177_
rlabel metal2 18814 24480 18814 24480 0 _0178_
rlabel metal1 19458 24718 19458 24718 0 _0179_
rlabel metal1 22908 24242 22908 24242 0 _0180_
rlabel metal1 22540 22066 22540 22066 0 _0181_
rlabel metal1 23092 23630 23092 23630 0 _0182_
rlabel viali 22862 22073 22862 22073 0 _0183_
rlabel metal1 22586 23664 22586 23664 0 _0184_
rlabel metal1 24242 23528 24242 23528 0 _0185_
rlabel metal1 23736 23834 23736 23834 0 _0186_
rlabel metal1 24702 23664 24702 23664 0 _0187_
rlabel metal1 22218 22066 22218 22066 0 _0188_
rlabel metal1 21804 22066 21804 22066 0 _0189_
rlabel metal1 22816 21930 22816 21930 0 _0190_
rlabel metal1 23644 21930 23644 21930 0 _0191_
rlabel metal1 24104 22066 24104 22066 0 _0192_
rlabel metal1 2484 15470 2484 15470 0 _0193_
rlabel metal1 21666 20400 21666 20400 0 _0194_
rlabel metal1 20930 20298 20930 20298 0 _0195_
rlabel metal2 22126 20196 22126 20196 0 _0196_
rlabel metal2 22218 20672 22218 20672 0 _0197_
rlabel metal1 21114 19822 21114 19822 0 _0198_
rlabel metal1 23552 20978 23552 20978 0 _0199_
rlabel metal1 22908 20434 22908 20434 0 _0200_
rlabel metal1 22540 20298 22540 20298 0 _0201_
rlabel metal1 22816 19278 22816 19278 0 _0202_
rlabel metal1 23184 19278 23184 19278 0 _0203_
rlabel metal1 18860 18938 18860 18938 0 _0204_
rlabel metal1 22126 19346 22126 19346 0 _0205_
rlabel metal1 18814 18870 18814 18870 0 _0206_
rlabel metal1 18403 18938 18403 18938 0 _0207_
rlabel metal1 9246 20400 9246 20400 0 _0208_
rlabel metal1 12926 15980 12926 15980 0 _0209_
rlabel metal1 20562 18870 20562 18870 0 _0210_
rlabel metal1 20884 20026 20884 20026 0 _0211_
rlabel metal1 18630 13430 18630 13430 0 _0212_
rlabel metal1 20930 19482 20930 19482 0 _0213_
rlabel metal2 20470 18938 20470 18938 0 _0214_
rlabel metal1 19826 18190 19826 18190 0 _0215_
rlabel metal1 19504 21046 19504 21046 0 _0216_
rlabel metal1 19642 20910 19642 20910 0 _0217_
rlabel metal1 18630 20910 18630 20910 0 _0218_
rlabel metal1 19182 20842 19182 20842 0 _0219_
rlabel metal1 18906 21114 18906 21114 0 _0220_
rlabel metal2 19918 16082 19918 16082 0 _0221_
rlabel metal2 11454 14654 11454 14654 0 _0222_
rlabel metal1 20930 13770 20930 13770 0 _0223_
rlabel metal1 19734 15572 19734 15572 0 _0224_
rlabel metal2 13938 14008 13938 14008 0 _0225_
rlabel metal1 20608 14994 20608 14994 0 _0226_
rlabel metal1 21160 14926 21160 14926 0 _0227_
rlabel metal1 21712 14926 21712 14926 0 _0228_
rlabel metal1 21482 15130 21482 15130 0 _0229_
rlabel metal1 20148 15538 20148 15538 0 _0230_
rlabel metal1 20148 13838 20148 13838 0 _0231_
rlabel metal1 19366 13940 19366 13940 0 _0232_
rlabel metal2 19550 13668 19550 13668 0 _0233_
rlabel metal1 19320 13362 19320 13362 0 _0234_
rlabel metal1 20746 13872 20746 13872 0 _0235_
rlabel metal1 21298 13362 21298 13362 0 _0236_
rlabel metal2 21666 13974 21666 13974 0 _0237_
rlabel metal1 18860 11798 18860 11798 0 _0238_
rlabel metal1 18722 12274 18722 12274 0 _0239_
rlabel metal1 18906 12172 18906 12172 0 _0240_
rlabel metal1 19504 12410 19504 12410 0 _0241_
rlabel metal1 20470 12240 20470 12240 0 _0242_
rlabel metal1 20700 12274 20700 12274 0 _0243_
rlabel metal1 14812 13294 14812 13294 0 _0244_
rlabel metal2 18906 13498 18906 13498 0 _0245_
rlabel metal1 16054 12682 16054 12682 0 _0246_
rlabel metal2 16330 13430 16330 13430 0 _0247_
rlabel metal1 15318 13158 15318 13158 0 _0248_
rlabel metal1 14582 12750 14582 12750 0 _0249_
rlabel metal1 16974 12784 16974 12784 0 _0250_
rlabel metal1 17618 12784 17618 12784 0 _0251_
rlabel metal1 17940 12750 17940 12750 0 _0252_
rlabel metal1 14628 11662 14628 11662 0 _0253_
rlabel metal1 14260 11594 14260 11594 0 _0254_
rlabel metal1 13695 11730 13695 11730 0 _0255_
rlabel metal1 14214 11526 14214 11526 0 _0256_
rlabel metal1 13938 11798 13938 11798 0 _0257_
rlabel metal2 13478 11679 13478 11679 0 _0258_
rlabel metal1 11546 10574 11546 10574 0 _0259_
rlabel metal2 12834 12444 12834 12444 0 _0260_
rlabel metal1 13616 13430 13616 13430 0 _0261_
rlabel metal1 13892 13430 13892 13430 0 _0262_
rlabel metal1 13662 12954 13662 12954 0 _0263_
rlabel via1 13746 12682 13746 12682 0 _0264_
rlabel metal2 13570 12410 13570 12410 0 _0265_
rlabel metal1 17204 10778 17204 10778 0 _0266_
rlabel metal1 15134 11798 15134 11798 0 _0267_
rlabel metal1 15594 11594 15594 11594 0 _0268_
rlabel metal2 15410 11390 15410 11390 0 _0269_
rlabel metal1 15594 11254 15594 11254 0 _0270_
rlabel metal1 15962 11220 15962 11220 0 _0271_
rlabel metal1 16146 11152 16146 11152 0 _0272_
rlabel metal1 4692 12410 4692 12410 0 _0273_
rlabel metal1 6302 12206 6302 12206 0 _0274_
rlabel metal1 3726 13362 3726 13362 0 _0275_
rlabel metal1 4186 12920 4186 12920 0 _0276_
rlabel metal1 2254 12784 2254 12784 0 _0277_
rlabel metal2 2070 13396 2070 13396 0 _0278_
rlabel metal1 4232 13430 4232 13430 0 _0279_
rlabel metal2 3818 13838 3818 13838 0 _0280_
rlabel metal1 3266 14960 3266 14960 0 _0281_
rlabel metal1 3450 14994 3450 14994 0 _0282_
rlabel metal1 3818 14892 3818 14892 0 _0283_
rlabel metal1 4416 14382 4416 14382 0 _0284_
rlabel metal1 2553 15538 2553 15538 0 _0285_
rlabel metal2 2162 16150 2162 16150 0 _0286_
rlabel metal2 3910 14977 3910 14977 0 _0287_
rlabel metal1 3174 14348 3174 14348 0 _0288_
rlabel metal1 4140 16218 4140 16218 0 _0289_
rlabel metal1 3818 16762 3818 16762 0 _0290_
rlabel metal1 3772 17102 3772 17102 0 _0291_
rlabel metal1 6072 15946 6072 15946 0 _0292_
rlabel metal1 3910 14994 3910 14994 0 _0293_
rlabel metal1 6164 12750 6164 12750 0 _0294_
rlabel metal1 9844 14926 9844 14926 0 _0295_
rlabel metal1 7682 12716 7682 12716 0 _0296_
rlabel metal1 7360 12818 7360 12818 0 _0297_
rlabel metal1 6670 12818 6670 12818 0 _0298_
rlabel metal1 5750 12954 5750 12954 0 _0299_
rlabel metal2 6026 14246 6026 14246 0 _0300_
rlabel metal1 6348 14450 6348 14450 0 _0301_
rlabel metal1 7728 12954 7728 12954 0 _0302_
rlabel metal1 6854 12308 6854 12308 0 _0303_
rlabel metal1 6900 11662 6900 11662 0 _0304_
rlabel metal1 7038 11764 7038 11764 0 _0305_
rlabel metal2 6762 11356 6762 11356 0 _0306_
rlabel metal1 7176 11186 7176 11186 0 _0307_
rlabel metal1 10488 11322 10488 11322 0 _0308_
rlabel metal1 10028 12750 10028 12750 0 _0309_
rlabel metal1 9522 12410 9522 12410 0 _0310_
rlabel metal1 10442 12682 10442 12682 0 _0311_
rlabel metal1 10810 12920 10810 12920 0 _0312_
rlabel metal2 10166 13090 10166 13090 0 _0313_
rlabel metal1 10534 11866 10534 11866 0 _0314_
rlabel metal1 9614 11730 9614 11730 0 _0315_
rlabel metal2 10442 11356 10442 11356 0 _0316_
rlabel metal2 9062 13124 9062 13124 0 _0317_
rlabel metal1 9246 11118 9246 11118 0 _0318_
rlabel metal1 9016 11118 9016 11118 0 _0319_
rlabel metal1 8418 11186 8418 11186 0 _0320_
rlabel metal2 10350 14841 10350 14841 0 _0321_
rlabel metal1 10350 14926 10350 14926 0 _0322_
rlabel metal1 10626 14858 10626 14858 0 _0323_
rlabel metal1 10672 14994 10672 14994 0 _0324_
rlabel metal1 10902 14858 10902 14858 0 _0325_
rlabel viali 10627 14450 10627 14450 0 _0326_
rlabel metal1 11178 13838 11178 13838 0 _0327_
rlabel metal1 17618 23290 17618 23290 0 _0328_
rlabel metal1 17342 23630 17342 23630 0 _0329_
rlabel metal1 18124 22950 18124 22950 0 _0330_
rlabel metal1 18515 23154 18515 23154 0 _0331_
rlabel metal1 17342 23086 17342 23086 0 _0332_
rlabel metal1 18124 23154 18124 23154 0 _0333_
rlabel metal1 18906 22746 18906 22746 0 _0334_
rlabel metal1 18262 23222 18262 23222 0 _0335_
rlabel metal1 17434 20910 17434 20910 0 _0336_
rlabel metal1 16974 20230 16974 20230 0 _0337_
rlabel metal2 16790 20672 16790 20672 0 _0338_
rlabel metal2 16974 19958 16974 19958 0 _0339_
rlabel metal2 17710 21692 17710 21692 0 _0340_
rlabel metal1 17099 21046 17099 21046 0 _0341_
rlabel metal1 14812 20910 14812 20910 0 _0342_
rlabel metal1 10350 21386 10350 21386 0 _0343_
rlabel metal1 11408 20774 11408 20774 0 _0344_
rlabel metal1 11224 20366 11224 20366 0 _0345_
rlabel metal1 9062 18156 9062 18156 0 _0346_
rlabel metal1 8188 18258 8188 18258 0 _0347_
rlabel metal1 8648 17714 8648 17714 0 _0348_
rlabel metal2 9062 19006 9062 19006 0 _0349_
rlabel metal2 8786 18054 8786 18054 0 _0350_
rlabel metal1 5106 22576 5106 22576 0 _0351_
rlabel viali 5198 22543 5198 22543 0 _0352_
rlabel metal1 4876 22202 4876 22202 0 _0353_
rlabel metal1 4692 22542 4692 22542 0 _0354_
rlabel metal1 6624 18190 6624 18190 0 _0355_
rlabel metal1 5842 18190 5842 18190 0 _0356_
rlabel metal1 5474 18122 5474 18122 0 _0357_
rlabel metal2 6854 16490 6854 16490 0 _0358_
rlabel metal1 7820 16558 7820 16558 0 _0359_
rlabel metal1 6578 15572 6578 15572 0 _0360_
rlabel metal1 6578 15674 6578 15674 0 _0361_
rlabel metal1 6072 17714 6072 17714 0 _0362_
rlabel metal1 8602 17612 8602 17612 0 _0363_
rlabel metal1 6992 18190 6992 18190 0 _0364_
rlabel metal1 7360 16218 7360 16218 0 _0365_
rlabel metal1 7176 16626 7176 16626 0 _0366_
rlabel metal1 8142 16762 8142 16762 0 _0367_
rlabel metal1 9338 17850 9338 17850 0 _0368_
rlabel metal1 7130 17850 7130 17850 0 _0369_
rlabel metal1 5658 16524 5658 16524 0 _0370_
rlabel metal1 6544 18258 6544 18258 0 _0371_
rlabel metal1 8786 18292 8786 18292 0 _0372_
rlabel metal1 9384 18122 9384 18122 0 _0373_
rlabel metal2 9890 17680 9890 17680 0 _0374_
rlabel metal1 9522 16218 9522 16218 0 _0375_
rlabel metal2 9798 16864 9798 16864 0 _0376_
rlabel metal2 10074 17510 10074 17510 0 _0377_
rlabel metal1 13064 16014 13064 16014 0 _0378_
rlabel metal1 13616 15538 13616 15538 0 _0379_
rlabel metal1 13248 15674 13248 15674 0 _0380_
rlabel metal1 10258 19278 10258 19278 0 _0381_
rlabel metal1 9844 19414 9844 19414 0 _0382_
rlabel metal1 10258 16626 10258 16626 0 _0383_
rlabel metal1 15548 16014 15548 16014 0 _0384_
rlabel metal1 15962 16592 15962 16592 0 _0385_
rlabel metal1 15410 17068 15410 17068 0 _0386_
rlabel metal1 15778 17136 15778 17136 0 _0387_
rlabel viali 15594 17102 15594 17102 0 _0388_
rlabel metal1 16192 16014 16192 16014 0 _0389_
rlabel metal1 15456 16762 15456 16762 0 _0390_
rlabel metal1 17066 17102 17066 17102 0 _0391_
rlabel viali 17701 16014 17701 16014 0 _0392_
rlabel viali 17436 15538 17436 15538 0 _0393_
rlabel metal2 17250 15300 17250 15300 0 _0394_
rlabel metal1 16974 15470 16974 15470 0 _0395_
rlabel metal1 17802 15674 17802 15674 0 _0396_
rlabel via2 17894 15997 17894 15997 0 _0397_
rlabel metal1 17204 18326 17204 18326 0 _0398_
rlabel metal1 17526 18394 17526 18394 0 _0399_
rlabel metal1 17250 18768 17250 18768 0 _0400_
rlabel metal1 17710 16422 17710 16422 0 _0401_
rlabel metal2 18630 16694 18630 16694 0 _0402_
rlabel metal1 18668 16694 18668 16694 0 _0403_
rlabel metal1 17388 16014 17388 16014 0 _0404_
rlabel metal1 17986 15946 17986 15946 0 _0405_
rlabel metal1 17480 16218 17480 16218 0 _0406_
rlabel metal2 17526 16864 17526 16864 0 _0407_
rlabel metal1 17802 16762 17802 16762 0 _0408_
rlabel metal1 17710 17136 17710 17136 0 _0409_
rlabel metal1 1794 20944 1794 20944 0 _0410_
rlabel metal1 1242 23290 1242 23290 0 _0411_
rlabel metal1 2070 22678 2070 22678 0 _0412_
rlabel metal2 2162 22984 2162 22984 0 _0413_
rlabel metal2 2898 23324 2898 23324 0 _0414_
rlabel metal1 3542 22950 3542 22950 0 _0415_
rlabel metal2 3266 22984 3266 22984 0 _0416_
rlabel metal1 3588 23154 3588 23154 0 _0417_
rlabel metal1 5428 23834 5428 23834 0 _0418_
rlabel metal1 4876 23834 4876 23834 0 _0419_
rlabel metal1 5428 20842 5428 20842 0 _0420_
rlabel metal1 5750 20366 5750 20366 0 _0421_
rlabel metal1 3174 21114 3174 21114 0 _0422_
rlabel metal1 3910 19210 3910 19210 0 _0423_
rlabel metal1 4600 20026 4600 20026 0 _0424_
rlabel metal1 4830 18802 4830 18802 0 _0425_
rlabel metal1 3174 19210 3174 19210 0 _0426_
rlabel metal1 2530 19312 2530 19312 0 _0427_
rlabel metal1 1748 20774 1748 20774 0 _0428_
rlabel metal1 2254 19210 2254 19210 0 _0429_
rlabel metal2 1978 19924 1978 19924 0 _0430_
rlabel metal1 1840 21114 1840 21114 0 _0431_
rlabel metal1 17802 21420 17802 21420 0 _0432_
rlabel metal1 16928 21590 16928 21590 0 _0433_
rlabel metal2 16330 21012 16330 21012 0 _0434_
rlabel metal1 15916 22678 15916 22678 0 _0435_
rlabel metal1 16054 21658 16054 21658 0 _0436_
rlabel metal1 15548 20978 15548 20978 0 _0437_
rlabel metal1 14904 26894 14904 26894 0 _0438_
rlabel metal1 14122 21658 14122 21658 0 _0439_
rlabel metal1 15088 26554 15088 26554 0 _0440_
rlabel metal2 14214 26962 14214 26962 0 _0441_
rlabel metal2 15042 27336 15042 27336 0 _0442_
rlabel metal1 15456 27642 15456 27642 0 _0443_
rlabel metal1 14214 24718 14214 24718 0 _0444_
rlabel metal1 14444 24378 14444 24378 0 _0445_
rlabel metal1 15042 24242 15042 24242 0 _0446_
rlabel metal1 14950 25432 14950 25432 0 _0447_
rlabel metal1 14996 24582 14996 24582 0 _0448_
rlabel metal1 15686 24718 15686 24718 0 _0449_
rlabel metal2 14582 17697 14582 17697 0 _0450_
rlabel metal2 15318 25568 15318 25568 0 _0451_
rlabel metal1 15824 25806 15824 25806 0 _0452_
rlabel metal1 13110 18156 13110 18156 0 _0453_
rlabel metal1 12236 18054 12236 18054 0 _0454_
rlabel metal1 12236 18394 12236 18394 0 _0455_
rlabel metal1 11730 17646 11730 17646 0 _0456_
rlabel metal2 13386 18564 13386 18564 0 _0457_
rlabel metal1 14260 17850 14260 17850 0 _0458_
rlabel metal2 14996 17714 14996 17714 0 _0459_
rlabel metal2 13662 20196 13662 20196 0 _0460_
rlabel metal1 13800 18802 13800 18802 0 _0461_
rlabel metal1 13340 20298 13340 20298 0 _0462_
rlabel metal1 18906 19244 18906 19244 0 clk
rlabel metal1 16284 19414 16284 19414 0 clknet_0_clk
rlabel metal1 1564 13362 1564 13362 0 clknet_3_0__leaf_clk
rlabel metal1 12489 14382 12489 14382 0 clknet_3_1__leaf_clk
rlabel metal1 1104 21454 1104 21454 0 clknet_3_2__leaf_clk
rlabel metal1 5244 21522 5244 21522 0 clknet_3_3__leaf_clk
rlabel metal1 14030 19890 14030 19890 0 clknet_3_4__leaf_clk
rlabel metal1 19412 16218 19412 16218 0 clknet_3_5__leaf_clk
rlabel metal1 15042 21658 15042 21658 0 clknet_3_6__leaf_clk
rlabel metal1 20056 25806 20056 25806 0 clknet_3_7__leaf_clk
rlabel viali 19361 26826 19361 26826 0 down_key.d
rlabel metal2 20378 26282 20378 26282 0 down_key.dff1
rlabel metal1 20194 22134 20194 22134 0 down_key.dff2
rlabel metal1 2530 14926 2530 14926 0 game.ballDirX
rlabel metal1 13892 14586 13892 14586 0 game.ballDirY
rlabel metal2 3818 12585 3818 12585 0 game.ballX\[0\]
rlabel metal1 4876 13430 4876 13430 0 game.ballX\[1\]
rlabel metal1 2070 15062 2070 15062 0 game.ballX\[2\]
rlabel metal2 6762 16830 6762 16830 0 game.ballX\[3\]
rlabel metal1 7590 14926 7590 14926 0 game.ballX\[4\]
rlabel metal1 7038 15946 7038 15946 0 game.ballX\[5\]
rlabel metal1 10442 12954 10442 12954 0 game.ballX\[6\]
rlabel metal1 8694 14892 8694 14892 0 game.ballX\[7\]
rlabel metal1 9522 19312 9522 19312 0 game.ballX\[8\]
rlabel metal2 20562 17408 20562 17408 0 game.ballY\[0\]
rlabel metal1 17296 18190 17296 18190 0 game.ballY\[1\]
rlabel metal1 18952 14518 18952 14518 0 game.ballY\[2\]
rlabel via1 19090 13821 19090 13821 0 game.ballY\[3\]
rlabel metal1 16882 13158 16882 13158 0 game.ballY\[4\]
rlabel metal1 14352 14926 14352 14926 0 game.ballY\[5\]
rlabel metal1 12834 12954 12834 12954 0 game.ballY\[6\]
rlabel metal1 14582 14314 14582 14314 0 game.ballY\[7\]
rlabel metal1 13202 27098 13202 27098 0 game.blue
rlabel metal1 7452 22746 7452 22746 0 game.col0
rlabel metal1 10994 21930 10994 21930 0 game.green
rlabel metal1 2254 23732 2254 23732 0 game.h\[0\]
rlabel metal1 4462 24072 4462 24072 0 game.h\[1\]
rlabel metal1 4600 24378 4600 24378 0 game.h\[2\]
rlabel metal1 5152 18394 5152 18394 0 game.h\[3\]
rlabel metal1 6854 21318 6854 21318 0 game.h\[4\]
rlabel metal1 5014 21420 5014 21420 0 game.h\[5\]
rlabel metal1 8556 20366 8556 20366 0 game.h\[6\]
rlabel metal1 8234 16694 8234 16694 0 game.h\[7\]
rlabel metal1 7544 19278 7544 19278 0 game.h\[8\]
rlabel metal1 2438 21930 2438 21930 0 game.h\[9\]
rlabel metal2 12006 20196 12006 20196 0 game.hit
rlabel metal1 7590 19992 7590 19992 0 game.hsync
rlabel metal1 10718 19278 10718 19278 0 game.inBallX
rlabel metal1 13524 16014 13524 16014 0 game.inBallY
rlabel metal1 8970 21522 8970 21522 0 game.inPaddle
rlabel metal1 21022 18836 21022 18836 0 game.new_game_n
rlabel metal1 9154 23664 9154 23664 0 game.offset\[0\]
rlabel metal1 9982 24276 9982 24276 0 game.offset\[1\]
rlabel metal1 11040 25738 11040 25738 0 game.offset\[2\]
rlabel metal1 4094 26928 4094 26928 0 game.offset\[3\]
rlabel metal1 3818 25908 3818 25908 0 game.offset\[4\]
rlabel metal1 17986 25262 17986 25262 0 game.paddle\[0\]
rlabel metal2 18814 23664 18814 23664 0 game.paddle\[1\]
rlabel metal1 17802 23698 17802 23698 0 game.paddle\[2\]
rlabel metal1 20562 23154 20562 23154 0 game.paddle\[3\]
rlabel metal1 19182 22984 19182 22984 0 game.paddle\[4\]
rlabel metal1 18515 23630 18515 23630 0 game.paddle\[5\]
rlabel metal1 17894 20570 17894 20570 0 game.paddle\[6\]
rlabel metal1 20286 18768 20286 18768 0 game.paddle\[7\]
rlabel metal1 18952 20978 18952 20978 0 game.paddle\[8\]
rlabel metal2 22954 24157 22954 24157 0 game.pause_n
rlabel metal1 9798 21930 9798 21930 0 game.red
rlabel metal2 2254 25279 2254 25279 0 game.row0
rlabel metal1 11454 20570 11454 20570 0 game.speaker
rlabel metal1 20608 27506 20608 27506 0 game.up_key_n
rlabel metal1 17158 27030 17158 27030 0 game.v\[0\]
rlabel metal1 14858 26792 14858 26792 0 game.v\[1\]
rlabel metal1 17526 18224 17526 18224 0 game.v\[2\]
rlabel metal1 18860 17102 18860 17102 0 game.v\[3\]
rlabel metal2 19136 18802 19136 18802 0 game.v\[4\]
rlabel metal1 13156 19414 13156 19414 0 game.v\[5\]
rlabel metal2 13294 19856 13294 19856 0 game.v\[6\]
rlabel metal1 13110 19822 13110 19822 0 game.v\[7\]
rlabel metal1 13524 17034 13524 17034 0 game.v\[8\]
rlabel metal1 14076 20842 14076 20842 0 game.v\[9\]
rlabel metal1 7360 27506 7360 27506 0 game.vsync
rlabel metal1 14076 17510 14076 17510 0 net1
rlabel metal1 24160 25330 24160 25330 0 net10
rlabel metal2 2070 21420 2070 21420 0 net11
rlabel metal2 3174 25568 3174 25568 0 net12
rlabel metal1 17388 10574 17388 10574 0 net13
rlabel metal1 10856 11186 10856 11186 0 net14
rlabel metal1 13110 16592 13110 16592 0 net15
rlabel metal1 16146 21420 16146 21420 0 net16
rlabel metal1 19228 19890 19228 19890 0 net17
rlabel metal1 14444 18802 14444 18802 0 net18
rlabel metal1 18078 25364 18078 25364 0 net19
rlabel metal1 23598 26894 23598 26894 0 net2
rlabel metal1 12282 17714 12282 17714 0 net20
rlabel metal1 15134 26452 15134 26452 0 net21
rlabel metal1 4094 18938 4094 18938 0 net22
rlabel metal1 11684 18802 11684 18802 0 net23
rlabel metal1 21390 27506 21390 27506 0 net3
rlabel metal1 20240 27982 20240 27982 0 net4
rlabel metal1 18216 26894 18216 26894 0 net5
rlabel metal1 14214 21420 14214 21420 0 net6
rlabel metal1 19683 27574 19683 27574 0 net7
rlabel metal1 20884 26010 20884 26010 0 net8
rlabel metal1 22954 27098 22954 27098 0 net9
rlabel via1 20925 26894 20925 26894 0 new_game.d
rlabel metal1 22402 26996 22402 26996 0 new_game.dff1
rlabel metal1 23276 27098 23276 27098 0 pause.d
rlabel metal1 24656 26962 24656 26962 0 pause.dff1
rlabel metal1 15272 27574 15272 27574 0 qb
rlabel metal1 12650 27506 12650 27506 0 qg
rlabel metal1 10994 27302 10994 27302 0 qr
rlabel metal1 25714 27982 25714 27982 0 rst_n
rlabel metal1 23828 27982 23828 27982 0 ui_in[0]
rlabel metal1 21712 27982 21712 27982 0 ui_in[1]
rlabel metal1 20470 28016 20470 28016 0 ui_in[2]
rlabel metal1 17572 27982 17572 27982 0 ui_in[3]
rlabel metal1 15640 27574 15640 27574 0 uo_out[0]
rlabel metal1 13248 27302 13248 27302 0 uo_out[1]
rlabel metal1 11408 28186 11408 28186 0 uo_out[2]
rlabel metal1 9200 27098 9200 27098 0 uo_out[3]
rlabel metal1 7176 27370 7176 27370 0 uo_out[4]
rlabel metal1 5290 27574 5290 27574 0 uo_out[5]
rlabel metal1 3588 27574 3588 27574 0 uo_out[6]
rlabel metal1 1380 27574 1380 27574 0 uo_out[7]
rlabel metal2 18354 27302 18354 27302 0 up_key.d
rlabel metal1 19182 27642 19182 27642 0 up_key.dff1
<< properties >>
string FIXED_BBOX 0 0 29000 29000
<< end >>
